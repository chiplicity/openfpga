magic
tech EFS8A
magscale 1 2
timestamp 1602873675
<< locali >>
rect 857 6647 891 16949
rect 949 14535 983 20213
rect 4019 17697 4146 17731
rect 15611 17697 15646 17731
rect 2547 16609 2582 16643
rect 23523 16609 23650 16643
rect 13737 16031 13771 16201
rect 13185 15929 13311 15963
rect 13277 15895 13311 15929
rect 10241 14807 10275 15113
rect 10333 14875 10367 14977
rect 4111 14433 4238 14467
rect 24627 14433 24662 14467
rect 22511 13345 22638 13379
rect 7481 12767 7515 12937
rect 21465 12767 21499 12937
rect 13363 12393 13369 12427
rect 13363 12325 13397 12393
rect 25087 12257 25122 12291
rect 949 9503 983 11509
rect 13455 11305 13461 11339
rect 12817 11135 12851 11305
rect 13455 11237 13489 11305
rect 25363 11169 25398 11203
rect 13455 10455 13489 10523
rect 13455 10421 13461 10455
rect 15577 9435 15611 9605
rect 24219 8041 24225 8075
rect 24219 7973 24253 8041
rect 18153 7735 18187 7973
rect 23213 7395 23247 7497
rect 22563 5865 22569 5899
rect 22563 5797 22597 5865
rect 12633 5559 12667 5661
rect 4445 5151 4479 5321
rect 8763 5015 8797 5083
rect 8763 4981 8769 5015
rect 21275 4777 21281 4811
rect 21275 4709 21309 4777
rect 1593 3417 1685 3451
rect 10609 3383 10643 3553
rect 18699 2601 18705 2635
rect 18699 2533 18733 2601
rect 23673 2295 23707 2533
<< viali >>
rect 1593 23817 1627 23851
rect 24777 23817 24811 23851
rect 1409 23613 1443 23647
rect 24593 23613 24627 23647
rect 25145 23613 25179 23647
rect 2053 23477 2087 23511
rect 1593 21641 1627 21675
rect 24777 21641 24811 21675
rect 1409 21437 1443 21471
rect 1961 21437 1995 21471
rect 24593 21437 24627 21471
rect 25145 21437 25179 21471
rect 1444 20349 1478 20383
rect 1869 20349 1903 20383
rect 949 20213 983 20247
rect 1547 20213 1581 20247
rect 857 16949 891 16983
rect 1444 19873 1478 19907
rect 1547 19669 1581 19703
rect 2237 19465 2271 19499
rect 2559 19397 2593 19431
rect 1476 19261 1510 19295
rect 1869 19261 1903 19295
rect 2488 19261 2522 19295
rect 1547 19125 1581 19159
rect 2973 19125 3007 19159
rect 1444 18785 1478 18819
rect 2456 18785 2490 18819
rect 1547 18581 1581 18615
rect 2559 18581 2593 18615
rect 2329 18241 2363 18275
rect 1444 18173 1478 18207
rect 2605 18173 2639 18207
rect 3868 18173 3902 18207
rect 6904 18173 6938 18207
rect 1869 18105 1903 18139
rect 4353 18105 4387 18139
rect 7297 18105 7331 18139
rect 1547 18037 1581 18071
rect 2789 18037 2823 18071
rect 3939 18037 3973 18071
rect 6975 18037 7009 18071
rect 1593 17833 1627 17867
rect 24777 17833 24811 17867
rect 1409 17697 1443 17731
rect 2580 17697 2614 17731
rect 3985 17697 4019 17731
rect 5156 17697 5190 17731
rect 6745 17697 6779 17731
rect 13461 17697 13495 17731
rect 13921 17697 13955 17731
rect 15577 17697 15611 17731
rect 24593 17697 24627 17731
rect 12357 17629 12391 17663
rect 14105 17629 14139 17663
rect 2651 17493 2685 17527
rect 4215 17493 4249 17527
rect 5227 17493 5261 17527
rect 6929 17493 6963 17527
rect 15715 17493 15749 17527
rect 2329 17289 2363 17323
rect 2559 17289 2593 17323
rect 13461 17289 13495 17323
rect 6975 17221 7009 17255
rect 9229 17221 9263 17255
rect 11805 17221 11839 17255
rect 3985 17153 4019 17187
rect 13001 17153 13035 17187
rect 15577 17153 15611 17187
rect 1444 17085 1478 17119
rect 1869 17085 1903 17119
rect 2488 17085 2522 17119
rect 2881 17085 2915 17119
rect 3500 17085 3534 17119
rect 4512 17085 4546 17119
rect 5524 17085 5558 17119
rect 6904 17085 6938 17119
rect 8815 17085 8849 17119
rect 8907 17085 8941 17119
rect 10860 17085 10894 17119
rect 11345 17085 11379 17119
rect 12265 17085 12299 17119
rect 12449 17085 12483 17119
rect 12909 17085 12943 17119
rect 14381 17085 14415 17119
rect 15025 17085 15059 17119
rect 15945 17085 15979 17119
rect 16405 17085 16439 17119
rect 4261 17017 4295 17051
rect 14289 17017 14323 17051
rect 1547 16949 1581 16983
rect 3249 16949 3283 16983
rect 3571 16949 3605 16983
rect 4583 16949 4617 16983
rect 4905 16949 4939 16983
rect 5273 16949 5307 16983
rect 5595 16949 5629 16983
rect 6009 16949 6043 16983
rect 6653 16949 6687 16983
rect 7389 16949 7423 16983
rect 7665 16949 7699 16983
rect 9781 16949 9815 16983
rect 10931 16949 10965 16983
rect 13921 16949 13955 16983
rect 16129 16949 16163 16983
rect 23765 16949 23799 16983
rect 24593 16949 24627 16983
rect 1593 16745 1627 16779
rect 7757 16745 7791 16779
rect 9965 16745 9999 16779
rect 13645 16745 13679 16779
rect 23719 16745 23753 16779
rect 1409 16609 1443 16643
rect 2513 16609 2547 16643
rect 4144 16609 4178 16643
rect 5641 16609 5675 16643
rect 6720 16609 6754 16643
rect 7849 16609 7883 16643
rect 8125 16609 8159 16643
rect 9689 16609 9723 16643
rect 10149 16609 10183 16643
rect 12633 16609 12667 16643
rect 13645 16609 13679 16643
rect 14105 16609 14139 16643
rect 15301 16609 15335 16643
rect 15577 16609 15611 16643
rect 16865 16609 16899 16643
rect 23489 16609 23523 16643
rect 24660 16609 24694 16643
rect 15761 16541 15795 16575
rect 20913 16541 20947 16575
rect 6791 16473 6825 16507
rect 15393 16473 15427 16507
rect 24731 16473 24765 16507
rect 2651 16405 2685 16439
rect 4215 16405 4249 16439
rect 5825 16405 5859 16439
rect 7481 16405 7515 16439
rect 10885 16405 10919 16439
rect 12265 16405 12299 16439
rect 13001 16405 13035 16439
rect 17049 16405 17083 16439
rect 1593 16201 1627 16235
rect 4675 16201 4709 16235
rect 8769 16201 8803 16235
rect 13737 16201 13771 16235
rect 13829 16201 13863 16235
rect 16313 16201 16347 16235
rect 16681 16201 16715 16235
rect 24593 16201 24627 16235
rect 25237 16201 25271 16235
rect 2053 16133 2087 16167
rect 11897 16133 11931 16167
rect 6285 16065 6319 16099
rect 12541 16065 12575 16099
rect 13553 16065 13587 16099
rect 17141 16133 17175 16167
rect 24133 16133 24167 16167
rect 15301 16065 15335 16099
rect 23029 16065 23063 16099
rect 1409 15997 1443 16031
rect 2559 15997 2593 16031
rect 2973 15997 3007 16031
rect 3592 15997 3626 16031
rect 4604 15997 4638 16031
rect 4997 15997 5031 16031
rect 5733 15997 5767 16031
rect 7941 15997 7975 16031
rect 8125 15997 8159 16031
rect 9137 15997 9171 16031
rect 9229 15997 9263 16031
rect 9781 15997 9815 16031
rect 10701 15997 10735 16031
rect 10793 15997 10827 16031
rect 11253 15997 11287 16031
rect 12449 15997 12483 16031
rect 12725 15997 12759 16031
rect 13737 15997 13771 16031
rect 14048 15997 14082 16031
rect 14841 15997 14875 16031
rect 15853 15997 15887 16031
rect 16957 15997 16991 16031
rect 17785 15997 17819 16031
rect 18061 15997 18095 16031
rect 18521 15997 18555 16031
rect 22620 15997 22654 16031
rect 24752 15997 24786 16031
rect 3341 15929 3375 15963
rect 3985 15929 4019 15963
rect 7573 15929 7607 15963
rect 11529 15929 11563 15963
rect 14151 15929 14185 15963
rect 22707 15929 22741 15963
rect 2651 15861 2685 15895
rect 3663 15861 3697 15895
rect 4445 15861 4479 15895
rect 5917 15861 5951 15895
rect 6561 15861 6595 15895
rect 7113 15861 7147 15895
rect 7941 15861 7975 15895
rect 9321 15861 9355 15895
rect 10241 15861 10275 15895
rect 12265 15861 12299 15895
rect 13277 15861 13311 15895
rect 15209 15861 15243 15895
rect 17417 15861 17451 15895
rect 18245 15861 18279 15895
rect 21097 15861 21131 15895
rect 23673 15861 23707 15895
rect 24823 15861 24857 15895
rect 1593 15657 1627 15691
rect 7573 15657 7607 15691
rect 13645 15657 13679 15691
rect 15761 15657 15795 15691
rect 9321 15589 9355 15623
rect 9965 15589 9999 15623
rect 14289 15589 14323 15623
rect 2053 15521 2087 15555
rect 2237 15521 2271 15555
rect 2789 15521 2823 15555
rect 4144 15521 4178 15555
rect 5124 15521 5158 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 8125 15521 8159 15555
rect 8401 15521 8435 15555
rect 10885 15521 10919 15555
rect 11069 15521 11103 15555
rect 12173 15521 12207 15555
rect 12449 15521 12483 15555
rect 13772 15521 13806 15555
rect 15301 15521 15335 15555
rect 15577 15521 15611 15555
rect 17233 15521 17267 15555
rect 18429 15521 18463 15555
rect 20980 15521 21014 15555
rect 23708 15521 23742 15555
rect 2329 15453 2363 15487
rect 7021 15453 7055 15487
rect 8585 15453 8619 15487
rect 11161 15453 11195 15487
rect 12633 15453 12667 15487
rect 15117 15453 15151 15487
rect 16865 15453 16899 15487
rect 19441 15453 19475 15487
rect 21925 15453 21959 15487
rect 24685 15453 24719 15487
rect 5227 15385 5261 15419
rect 12265 15385 12299 15419
rect 13875 15385 13909 15419
rect 15393 15385 15427 15419
rect 4215 15317 4249 15351
rect 5549 15317 5583 15351
rect 16313 15317 16347 15351
rect 18613 15317 18647 15351
rect 21051 15317 21085 15351
rect 23811 15317 23845 15351
rect 2973 15113 3007 15147
rect 6377 15113 6411 15147
rect 10241 15113 10275 15147
rect 22293 15113 22327 15147
rect 24777 15113 24811 15147
rect 8861 15045 8895 15079
rect 1869 14909 1903 14943
rect 2237 14909 2271 14943
rect 2513 14909 2547 14943
rect 3433 14909 3467 14943
rect 3525 14909 3559 14943
rect 3985 14909 4019 14943
rect 5365 14909 5399 14943
rect 5641 14909 5675 14943
rect 7757 14909 7791 14943
rect 7941 14909 7975 14943
rect 9045 14909 9079 14943
rect 9505 14909 9539 14943
rect 7389 14841 7423 14875
rect 8585 14841 8619 14875
rect 17785 15045 17819 15079
rect 19809 15045 19843 15079
rect 10333 14977 10367 15011
rect 16037 14977 16071 15011
rect 10609 14909 10643 14943
rect 11069 14909 11103 14943
rect 11897 14909 11931 14943
rect 12265 14909 12299 14943
rect 12817 14909 12851 14943
rect 14105 14909 14139 14943
rect 15577 14909 15611 14943
rect 15669 14909 15703 14943
rect 15853 14909 15887 14943
rect 18061 14909 18095 14943
rect 18521 14909 18555 14943
rect 19625 14909 19659 14943
rect 20856 14909 20890 14943
rect 20959 14909 20993 14943
rect 21884 14909 21918 14943
rect 24593 14909 24627 14943
rect 25145 14909 25179 14943
rect 10333 14841 10367 14875
rect 10425 14841 10459 14875
rect 13185 14841 13219 14875
rect 14749 14841 14783 14875
rect 15117 14841 15151 14875
rect 20085 14841 20119 14875
rect 21281 14841 21315 14875
rect 21971 14841 22005 14875
rect 2053 14773 2087 14807
rect 3617 14773 3651 14807
rect 4537 14773 4571 14807
rect 4905 14773 4939 14807
rect 5181 14773 5215 14807
rect 7573 14773 7607 14807
rect 9321 14773 9355 14807
rect 10149 14773 10183 14807
rect 10241 14773 10275 14807
rect 10701 14773 10735 14807
rect 13461 14773 13495 14807
rect 13921 14773 13955 14807
rect 15485 14773 15519 14807
rect 16957 14773 16991 14807
rect 18153 14773 18187 14807
rect 19073 14773 19107 14807
rect 21741 14773 21775 14807
rect 23857 14773 23891 14807
rect 1869 14569 1903 14603
rect 3525 14569 3559 14603
rect 5181 14569 5215 14603
rect 5457 14569 5491 14603
rect 6469 14569 6503 14603
rect 7757 14569 7791 14603
rect 10793 14569 10827 14603
rect 12633 14569 12667 14603
rect 16405 14569 16439 14603
rect 23719 14569 23753 14603
rect 949 14501 983 14535
rect 2329 14501 2363 14535
rect 2421 14501 2455 14535
rect 9873 14501 9907 14535
rect 11437 14501 11471 14535
rect 12357 14501 12391 14535
rect 4077 14433 4111 14467
rect 5549 14433 5583 14467
rect 5917 14433 5951 14467
rect 8125 14433 8159 14467
rect 8309 14433 8343 14467
rect 12817 14433 12851 14467
rect 13093 14433 13127 14467
rect 15301 14433 15335 14467
rect 15577 14433 15611 14467
rect 17392 14433 17426 14467
rect 18889 14433 18923 14467
rect 20948 14433 20982 14467
rect 21992 14433 22026 14467
rect 23648 14433 23682 14467
rect 24593 14433 24627 14467
rect 2697 14365 2731 14399
rect 8585 14365 8619 14399
rect 9781 14365 9815 14399
rect 10425 14365 10459 14399
rect 11345 14365 11379 14399
rect 11989 14365 12023 14399
rect 13277 14365 13311 14399
rect 16037 14365 16071 14399
rect 12909 14297 12943 14331
rect 15393 14297 15427 14331
rect 22063 14297 22097 14331
rect 4307 14229 4341 14263
rect 4721 14229 4755 14263
rect 6929 14229 6963 14263
rect 9045 14229 9079 14263
rect 11161 14229 11195 14263
rect 13829 14229 13863 14263
rect 14657 14229 14691 14263
rect 15117 14229 15151 14263
rect 16773 14229 16807 14263
rect 17463 14229 17497 14263
rect 18153 14229 18187 14263
rect 18613 14229 18647 14263
rect 19441 14229 19475 14263
rect 21051 14229 21085 14263
rect 24731 14229 24765 14263
rect 1593 14025 1627 14059
rect 2053 14025 2087 14059
rect 4905 14025 4939 14059
rect 7941 14025 7975 14059
rect 11345 14025 11379 14059
rect 12265 14025 12299 14059
rect 18889 14025 18923 14059
rect 24501 14025 24535 14059
rect 16221 13957 16255 13991
rect 18245 13957 18279 13991
rect 24777 13957 24811 13991
rect 3525 13889 3559 13923
rect 5365 13889 5399 13923
rect 6101 13889 6135 13923
rect 9689 13889 9723 13923
rect 10885 13889 10919 13923
rect 11621 13889 11655 13923
rect 12541 13889 12575 13923
rect 12817 13889 12851 13923
rect 25145 13889 25179 13923
rect 1409 13821 1443 13855
rect 2421 13821 2455 13855
rect 6561 13821 6595 13855
rect 6837 13821 6871 13855
rect 7297 13821 7331 13855
rect 8728 13821 8762 13855
rect 9505 13821 9539 13855
rect 13829 13821 13863 13855
rect 14381 13821 14415 13855
rect 15301 13821 15335 13855
rect 16129 13821 16163 13855
rect 16405 13821 16439 13855
rect 18061 13821 18095 13855
rect 18521 13821 18555 13855
rect 19441 13821 19475 13855
rect 20764 13821 20798 13855
rect 21189 13821 21223 13855
rect 22636 13821 22670 13855
rect 24593 13821 24627 13855
rect 2881 13753 2915 13787
rect 2973 13753 3007 13787
rect 3801 13753 3835 13787
rect 5089 13753 5123 13787
rect 5181 13753 5215 13787
rect 10051 13753 10085 13787
rect 12610 13753 12644 13787
rect 14702 13753 14736 13787
rect 15577 13753 15611 13787
rect 21557 13753 21591 13787
rect 4169 13685 4203 13719
rect 6929 13685 6963 13719
rect 8217 13685 8251 13719
rect 8815 13685 8849 13719
rect 9229 13685 9263 13719
rect 10609 13685 10643 13719
rect 13461 13685 13495 13719
rect 14197 13685 14231 13719
rect 15945 13685 15979 13719
rect 16589 13685 16623 13719
rect 17417 13685 17451 13719
rect 19441 13685 19475 13719
rect 20867 13685 20901 13719
rect 22017 13685 22051 13719
rect 22707 13685 22741 13719
rect 23029 13685 23063 13719
rect 23857 13685 23891 13719
rect 1685 13481 1719 13515
rect 2053 13481 2087 13515
rect 3157 13481 3191 13515
rect 3525 13481 3559 13515
rect 4905 13481 4939 13515
rect 5917 13481 5951 13515
rect 8769 13481 8803 13515
rect 9873 13481 9907 13515
rect 12081 13481 12115 13515
rect 12449 13481 12483 13515
rect 14013 13481 14047 13515
rect 24777 13481 24811 13515
rect 2599 13413 2633 13447
rect 5318 13413 5352 13447
rect 8211 13413 8245 13447
rect 9505 13413 9539 13447
rect 11523 13413 11557 13447
rect 15622 13413 15656 13447
rect 18797 13413 18831 13447
rect 2237 13345 2271 13379
rect 4997 13345 5031 13379
rect 6904 13345 6938 13379
rect 7849 13345 7883 13379
rect 12909 13345 12943 13379
rect 13185 13345 13219 13379
rect 15301 13345 15335 13379
rect 17049 13345 17083 13379
rect 17325 13345 17359 13379
rect 21005 13345 21039 13379
rect 22477 13345 22511 13379
rect 23648 13345 23682 13379
rect 24593 13345 24627 13379
rect 10149 13277 10183 13311
rect 11161 13277 11195 13311
rect 13369 13277 13403 13311
rect 14473 13277 14507 13311
rect 17785 13277 17819 13311
rect 18705 13277 18739 13311
rect 13001 13209 13035 13243
rect 15025 13209 15059 13243
rect 17141 13209 17175 13243
rect 19257 13209 19291 13243
rect 20177 13209 20211 13243
rect 3801 13141 3835 13175
rect 6975 13141 7009 13175
rect 10701 13141 10735 13175
rect 16221 13141 16255 13175
rect 16497 13141 16531 13175
rect 21373 13141 21407 13175
rect 22707 13141 22741 13175
rect 23719 13141 23753 13175
rect 3157 12937 3191 12971
rect 4721 12937 4755 12971
rect 5089 12937 5123 12971
rect 7113 12937 7147 12971
rect 7481 12937 7515 12971
rect 10517 12937 10551 12971
rect 14933 12937 14967 12971
rect 17785 12937 17819 12971
rect 18521 12937 18555 12971
rect 19717 12937 19751 12971
rect 21465 12937 21499 12971
rect 21557 12937 21591 12971
rect 24409 12937 24443 12971
rect 3433 12869 3467 12903
rect 2145 12801 2179 12835
rect 3709 12801 3743 12835
rect 3985 12801 4019 12835
rect 5549 12801 5583 12835
rect 8125 12869 8159 12903
rect 9505 12869 9539 12903
rect 11713 12869 11747 12903
rect 16221 12869 16255 12903
rect 19257 12869 19291 12903
rect 21189 12869 21223 12903
rect 8217 12801 8251 12835
rect 10977 12801 11011 12835
rect 12679 12801 12713 12835
rect 20269 12801 20303 12835
rect 20637 12801 20671 12835
rect 24777 12869 24811 12903
rect 7272 12733 7306 12767
rect 7481 12733 7515 12767
rect 12576 12733 12610 12767
rect 13553 12733 13587 12767
rect 21465 12733 21499 12767
rect 21741 12733 21775 12767
rect 22201 12733 22235 12767
rect 24593 12733 24627 12767
rect 25145 12733 25179 12767
rect 1961 12665 1995 12699
rect 2237 12665 2271 12699
rect 2789 12665 2823 12699
rect 3801 12665 3835 12699
rect 5273 12665 5307 12699
rect 5365 12665 5399 12699
rect 8579 12665 8613 12699
rect 10149 12665 10183 12699
rect 10701 12665 10735 12699
rect 10793 12665 10827 12699
rect 13915 12665 13949 12699
rect 15301 12665 15335 12699
rect 15669 12665 15703 12699
rect 15761 12665 15795 12699
rect 17417 12665 17451 12699
rect 18705 12665 18739 12699
rect 18797 12665 18831 12699
rect 20361 12665 20395 12699
rect 6193 12597 6227 12631
rect 7343 12597 7377 12631
rect 7757 12597 7791 12631
rect 9137 12597 9171 12631
rect 12173 12597 12207 12631
rect 13001 12597 13035 12631
rect 13369 12597 13403 12631
rect 14473 12597 14507 12631
rect 16589 12597 16623 12631
rect 17049 12597 17083 12631
rect 19993 12597 20027 12631
rect 21833 12597 21867 12631
rect 22753 12597 22787 12631
rect 23949 12597 23983 12631
rect 1685 12393 1719 12427
rect 2053 12393 2087 12427
rect 3709 12393 3743 12427
rect 7941 12393 7975 12427
rect 9045 12393 9079 12427
rect 11805 12393 11839 12427
rect 13369 12393 13403 12427
rect 14289 12393 14323 12427
rect 18705 12393 18739 12427
rect 18981 12393 19015 12427
rect 20729 12393 20763 12427
rect 2421 12325 2455 12359
rect 5911 12325 5945 12359
rect 8125 12325 8159 12359
rect 8217 12325 8251 12359
rect 10517 12325 10551 12359
rect 10609 12325 10643 12359
rect 15485 12325 15519 12359
rect 16037 12325 16071 12359
rect 18106 12325 18140 12359
rect 4077 12257 4111 12291
rect 5273 12257 5307 12291
rect 6469 12257 6503 12291
rect 8769 12257 8803 12291
rect 12024 12257 12058 12291
rect 19349 12257 19383 12291
rect 19876 12257 19910 12291
rect 21281 12257 21315 12291
rect 23581 12257 23615 12291
rect 25053 12257 25087 12291
rect 2329 12189 2363 12223
rect 2605 12189 2639 12223
rect 5549 12189 5583 12223
rect 10793 12189 10827 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 15393 12189 15427 12223
rect 17785 12189 17819 12223
rect 23489 12189 23523 12223
rect 4261 12121 4295 12155
rect 12127 12053 12161 12087
rect 12541 12053 12575 12087
rect 13921 12053 13955 12087
rect 15117 12053 15151 12087
rect 16313 12053 16347 12087
rect 19947 12053 19981 12087
rect 21465 12053 21499 12087
rect 25191 12053 25225 12087
rect 2881 11849 2915 11883
rect 3157 11849 3191 11883
rect 3525 11849 3559 11883
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 6285 11849 6319 11883
rect 8125 11849 8159 11883
rect 10241 11849 10275 11883
rect 11437 11849 11471 11883
rect 11897 11849 11931 11883
rect 13461 11849 13495 11883
rect 15393 11849 15427 11883
rect 17509 11849 17543 11883
rect 17785 11849 17819 11883
rect 19165 11849 19199 11883
rect 19441 11849 19475 11883
rect 21097 11849 21131 11883
rect 21373 11849 21407 11883
rect 23489 11849 23523 11883
rect 25421 11849 25455 11883
rect 6561 11781 6595 11815
rect 19901 11781 19935 11815
rect 20637 11781 20671 11815
rect 1961 11713 1995 11747
rect 3801 11713 3835 11747
rect 4077 11713 4111 11747
rect 6929 11713 6963 11747
rect 7205 11713 7239 11747
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 12541 11713 12575 11747
rect 15025 11713 15059 11747
rect 16405 11713 16439 11747
rect 20085 11713 20119 11747
rect 21649 11713 21683 11747
rect 21925 11713 21959 11747
rect 5800 11645 5834 11679
rect 8769 11645 8803 11679
rect 8953 11645 8987 11679
rect 12449 11645 12483 11679
rect 12725 11645 12759 11679
rect 18245 11645 18279 11679
rect 23121 11645 23155 11679
rect 23765 11645 23799 11679
rect 25237 11645 25271 11679
rect 25789 11645 25823 11679
rect 1869 11577 1903 11611
rect 2282 11577 2316 11611
rect 3893 11577 3927 11611
rect 7021 11577 7055 11611
rect 10609 11577 10643 11611
rect 14381 11577 14415 11611
rect 14473 11577 14507 11611
rect 15945 11577 15979 11611
rect 16037 11577 16071 11611
rect 18566 11577 18600 11611
rect 20177 11577 20211 11611
rect 21741 11577 21775 11611
rect 25145 11577 25179 11611
rect 949 11509 983 11543
rect 4813 11509 4847 11543
rect 5871 11509 5905 11543
rect 9137 11509 9171 11543
rect 9873 11509 9907 11543
rect 12173 11509 12207 11543
rect 12909 11509 12943 11543
rect 14197 11509 14231 11543
rect 15761 11509 15795 11543
rect 17141 11509 17175 11543
rect 24133 11509 24167 11543
rect 1409 11305 1443 11339
rect 2329 11305 2363 11339
rect 3801 11305 3835 11339
rect 4997 11305 5031 11339
rect 6377 11305 6411 11339
rect 6837 11305 6871 11339
rect 7665 11305 7699 11339
rect 10241 11305 10275 11339
rect 12817 11305 12851 11339
rect 12909 11305 12943 11339
rect 13461 11305 13495 11339
rect 14381 11305 14415 11339
rect 15117 11305 15151 11339
rect 17233 11305 17267 11339
rect 20269 11305 20303 11339
rect 22017 11305 22051 11339
rect 2605 11237 2639 11271
rect 3157 11237 3191 11271
rect 5819 11237 5853 11271
rect 8211 11237 8245 11271
rect 10609 11237 10643 11271
rect 4077 11169 4111 11203
rect 5457 11169 5491 11203
rect 7849 11169 7883 11203
rect 12116 11169 12150 11203
rect 12219 11169 12253 11203
rect 15669 11237 15703 11271
rect 21189 11237 21223 11271
rect 21741 11237 21775 11271
rect 17417 11169 17451 11203
rect 17877 11169 17911 11203
rect 17969 11169 18003 11203
rect 18521 11169 18555 11203
rect 19876 11169 19910 11203
rect 22604 11169 22638 11203
rect 23857 11169 23891 11203
rect 25329 11169 25363 11203
rect 2513 11101 2547 11135
rect 10517 11101 10551 11135
rect 10793 11101 10827 11135
rect 12817 11101 12851 11135
rect 13093 11101 13127 11135
rect 15577 11101 15611 11135
rect 16037 11101 16071 11135
rect 21097 11101 21131 11135
rect 23765 11101 23799 11135
rect 4261 11033 4295 11067
rect 25467 11033 25501 11067
rect 1869 10965 1903 10999
rect 8769 10965 8803 10999
rect 9965 10965 9999 10999
rect 12633 10965 12667 10999
rect 14013 10965 14047 10999
rect 18889 10965 18923 10999
rect 19349 10965 19383 10999
rect 19947 10965 19981 10999
rect 22707 10965 22741 10999
rect 2973 10761 3007 10795
rect 6285 10761 6319 10795
rect 7941 10761 7975 10795
rect 9321 10761 9355 10795
rect 11253 10761 11287 10795
rect 14013 10761 14047 10795
rect 17509 10761 17543 10795
rect 17877 10761 17911 10795
rect 19625 10761 19659 10795
rect 20729 10761 20763 10795
rect 21005 10761 21039 10795
rect 21373 10761 21407 10795
rect 22569 10761 22603 10795
rect 23121 10761 23155 10795
rect 23489 10761 23523 10795
rect 24961 10761 24995 10795
rect 6975 10693 7009 10727
rect 16037 10693 16071 10727
rect 18705 10693 18739 10727
rect 1685 10625 1719 10659
rect 2329 10625 2363 10659
rect 3157 10625 3191 10659
rect 4997 10625 5031 10659
rect 5273 10625 5307 10659
rect 8125 10625 8159 10659
rect 9689 10625 9723 10659
rect 10241 10625 10275 10659
rect 12081 10625 12115 10659
rect 13093 10625 13127 10659
rect 14289 10625 14323 10659
rect 15301 10625 15335 10659
rect 16957 10625 16991 10659
rect 18153 10625 18187 10659
rect 21649 10625 21683 10659
rect 24041 10625 24075 10659
rect 24317 10625 24351 10659
rect 25421 10625 25455 10659
rect 4077 10557 4111 10591
rect 4721 10557 4755 10591
rect 6872 10557 6906 10591
rect 7297 10557 7331 10591
rect 19809 10557 19843 10591
rect 25580 10557 25614 10591
rect 1777 10489 1811 10523
rect 3478 10489 3512 10523
rect 5089 10489 5123 10523
rect 6009 10489 6043 10523
rect 8446 10489 8480 10523
rect 9965 10489 9999 10523
rect 10057 10489 10091 10523
rect 10977 10489 11011 10523
rect 15485 10489 15519 10523
rect 15577 10489 15611 10523
rect 16497 10489 16531 10523
rect 18245 10489 18279 10523
rect 20130 10489 20164 10523
rect 21741 10489 21775 10523
rect 22293 10489 22327 10523
rect 24133 10489 24167 10523
rect 2605 10421 2639 10455
rect 4445 10421 4479 10455
rect 9045 10421 9079 10455
rect 13001 10421 13035 10455
rect 13461 10421 13495 10455
rect 14933 10421 14967 10455
rect 16865 10421 16899 10455
rect 19257 10421 19291 10455
rect 25651 10421 25685 10455
rect 26065 10421 26099 10455
rect 1547 10217 1581 10251
rect 2329 10217 2363 10251
rect 3525 10217 3559 10251
rect 5733 10217 5767 10251
rect 7849 10217 7883 10251
rect 15117 10217 15151 10251
rect 19165 10217 19199 10251
rect 21833 10217 21867 10251
rect 22109 10217 22143 10251
rect 24593 10217 24627 10251
rect 2513 10149 2547 10183
rect 2605 10149 2639 10183
rect 4169 10149 4203 10183
rect 4261 10149 4295 10183
rect 8125 10149 8159 10183
rect 8217 10149 8251 10183
rect 8769 10149 8803 10183
rect 11345 10149 11379 10183
rect 11897 10149 11931 10183
rect 13185 10149 13219 10183
rect 13737 10149 13771 10183
rect 15485 10149 15519 10183
rect 18889 10149 18923 10183
rect 21234 10149 21268 10183
rect 23581 10149 23615 10183
rect 23673 10149 23707 10183
rect 24225 10149 24259 10183
rect 1476 10081 1510 10115
rect 5917 10081 5951 10115
rect 6193 10081 6227 10115
rect 9724 10081 9758 10115
rect 17693 10081 17727 10115
rect 17877 10081 17911 10115
rect 18245 10081 18279 10115
rect 18797 10081 18831 10115
rect 19768 10081 19802 10115
rect 25120 10081 25154 10115
rect 3157 10013 3191 10047
rect 4445 10013 4479 10047
rect 10149 10013 10183 10047
rect 11253 10013 11287 10047
rect 13645 10013 13679 10047
rect 15393 10013 15427 10047
rect 15669 10013 15703 10047
rect 19855 10013 19889 10047
rect 20913 10013 20947 10047
rect 12725 9945 12759 9979
rect 14197 9945 14231 9979
rect 16773 9945 16807 9979
rect 17141 9945 17175 9979
rect 19533 9945 19567 9979
rect 1961 9877 1995 9911
rect 5273 9877 5307 9911
rect 9827 9877 9861 9911
rect 10885 9877 10919 9911
rect 16313 9877 16347 9911
rect 20269 9877 20303 9911
rect 22569 9877 22603 9911
rect 25191 9877 25225 9911
rect 4445 9673 4479 9707
rect 5089 9673 5123 9707
rect 6193 9673 6227 9707
rect 8401 9673 8435 9707
rect 9045 9673 9079 9707
rect 10149 9673 10183 9707
rect 11805 9673 11839 9707
rect 13093 9673 13127 9707
rect 13461 9673 13495 9707
rect 14657 9673 14691 9707
rect 15393 9673 15427 9707
rect 18521 9673 18555 9707
rect 21005 9673 21039 9707
rect 21465 9673 21499 9707
rect 22661 9673 22695 9707
rect 23121 9673 23155 9707
rect 23489 9673 23523 9707
rect 24041 9673 24075 9707
rect 10609 9605 10643 9639
rect 12725 9605 12759 9639
rect 15577 9605 15611 9639
rect 15669 9605 15703 9639
rect 17141 9605 17175 9639
rect 22293 9605 22327 9639
rect 3065 9537 3099 9571
rect 3433 9537 3467 9571
rect 5273 9537 5307 9571
rect 8125 9537 8159 9571
rect 9229 9537 9263 9571
rect 10885 9537 10919 9571
rect 11529 9537 11563 9571
rect 13645 9537 13679 9571
rect 14289 9537 14323 9571
rect 15025 9537 15059 9571
rect 949 9469 983 9503
rect 1685 9469 1719 9503
rect 1961 9469 1995 9503
rect 6653 9469 6687 9503
rect 7113 9469 7147 9503
rect 7297 9469 7331 9503
rect 12541 9469 12575 9503
rect 15945 9537 15979 9571
rect 16405 9537 16439 9571
rect 17509 9537 17543 9571
rect 21741 9537 21775 9571
rect 24317 9537 24351 9571
rect 24593 9537 24627 9571
rect 17785 9469 17819 9503
rect 18705 9469 18739 9503
rect 19165 9469 19199 9503
rect 19533 9469 19567 9503
rect 19901 9469 19935 9503
rect 2881 9401 2915 9435
rect 3157 9401 3191 9435
rect 5365 9401 5399 9435
rect 5917 9401 5951 9435
rect 9321 9401 9355 9435
rect 9873 9401 9907 9435
rect 10977 9401 11011 9435
rect 13737 9401 13771 9435
rect 15577 9401 15611 9435
rect 16037 9401 16071 9435
rect 21833 9401 21867 9435
rect 24409 9401 24443 9435
rect 1685 9333 1719 9367
rect 2421 9333 2455 9367
rect 4169 9333 4203 9367
rect 6929 9333 6963 9367
rect 12265 9333 12299 9367
rect 18981 9333 19015 9367
rect 20453 9333 20487 9367
rect 25329 9333 25363 9367
rect 2973 9129 3007 9163
rect 3341 9129 3375 9163
rect 5089 9129 5123 9163
rect 6193 9129 6227 9163
rect 7159 9129 7193 9163
rect 7849 9129 7883 9163
rect 9229 9129 9263 9163
rect 10195 9129 10229 9163
rect 14197 9129 14231 9163
rect 16313 9129 16347 9163
rect 18061 9129 18095 9163
rect 18429 9129 18463 9163
rect 21649 9129 21683 9163
rect 22937 9129 22971 9163
rect 25559 9129 25593 9163
rect 2098 9061 2132 9095
rect 3709 9061 3743 9095
rect 5635 9061 5669 9095
rect 6929 9061 6963 9095
rect 8125 9061 8159 9095
rect 8217 9061 8251 9095
rect 11431 9061 11465 9095
rect 19993 9061 20027 9095
rect 22338 9061 22372 9095
rect 24041 9061 24075 9095
rect 4077 8993 4111 9027
rect 5273 8993 5307 9027
rect 7088 8993 7122 9027
rect 10092 8993 10126 9027
rect 11069 8993 11103 9027
rect 11989 8993 12023 9027
rect 13461 8993 13495 9027
rect 13921 8993 13955 9027
rect 16497 8993 16531 9027
rect 16681 8993 16715 9027
rect 17141 8993 17175 9027
rect 17601 8993 17635 9027
rect 18521 8993 18555 9027
rect 18981 8993 19015 9027
rect 19349 8993 19383 9027
rect 19717 8993 19751 9027
rect 20729 8993 20763 9027
rect 21072 8993 21106 9027
rect 23673 8993 23707 9027
rect 25488 8993 25522 9027
rect 1777 8925 1811 8959
rect 8769 8925 8803 8959
rect 10609 8925 10643 8959
rect 12817 8925 12851 8959
rect 20269 8925 20303 8959
rect 22017 8925 22051 8959
rect 23949 8925 23983 8959
rect 24225 8925 24259 8959
rect 4261 8857 4295 8891
rect 12449 8857 12483 8891
rect 1685 8789 1719 8823
rect 2697 8789 2731 8823
rect 15761 8789 15795 8823
rect 16129 8789 16163 8823
rect 21143 8789 21177 8823
rect 4353 8585 4387 8619
rect 4721 8585 4755 8619
rect 7849 8585 7883 8619
rect 8309 8585 8343 8619
rect 9781 8585 9815 8619
rect 11621 8585 11655 8619
rect 13461 8585 13495 8619
rect 15301 8585 15335 8619
rect 16865 8585 16899 8619
rect 17233 8585 17267 8619
rect 18245 8585 18279 8619
rect 22385 8585 22419 8619
rect 22753 8585 22787 8619
rect 23489 8585 23523 8619
rect 24869 8585 24903 8619
rect 25605 8585 25639 8619
rect 10057 8517 10091 8551
rect 16405 8517 16439 8551
rect 17877 8517 17911 8551
rect 20821 8517 20855 8551
rect 2605 8449 2639 8483
rect 5549 8449 5583 8483
rect 6193 8449 6227 8483
rect 6929 8449 6963 8483
rect 7205 8449 7239 8483
rect 8861 8449 8895 8483
rect 10701 8449 10735 8483
rect 12541 8449 12575 8483
rect 14565 8449 14599 8483
rect 20545 8449 20579 8483
rect 21465 8449 21499 8483
rect 21833 8449 21867 8483
rect 23949 8449 23983 8483
rect 24225 8449 24259 8483
rect 18061 8381 18095 8415
rect 18521 8381 18555 8415
rect 19073 8381 19107 8415
rect 19533 8381 19567 8415
rect 19901 8381 19935 8415
rect 20269 8381 20303 8415
rect 25421 8381 25455 8415
rect 25973 8381 26007 8415
rect 2329 8313 2363 8347
rect 2421 8313 2455 8347
rect 3709 8313 3743 8347
rect 5273 8313 5307 8347
rect 5365 8313 5399 8347
rect 7021 8313 7055 8347
rect 9182 8313 9216 8347
rect 10793 8313 10827 8347
rect 11345 8313 11379 8347
rect 12633 8313 12667 8347
rect 13185 8313 13219 8347
rect 14289 8313 14323 8347
rect 14381 8313 14415 8347
rect 15853 8313 15887 8347
rect 15945 8313 15979 8347
rect 21557 8313 21591 8347
rect 24041 8313 24075 8347
rect 1869 8245 1903 8279
rect 3249 8245 3283 8279
rect 3801 8245 3835 8279
rect 5089 8245 5123 8279
rect 6653 8245 6687 8279
rect 8769 8245 8803 8279
rect 10517 8245 10551 8279
rect 12265 8245 12299 8279
rect 14105 8245 14139 8279
rect 15669 8245 15703 8279
rect 18889 8245 18923 8279
rect 21189 8245 21223 8279
rect 25329 8245 25363 8279
rect 1777 8041 1811 8075
rect 2973 8041 3007 8075
rect 6929 8041 6963 8075
rect 7849 8041 7883 8075
rect 11069 8041 11103 8075
rect 14289 8041 14323 8075
rect 16129 8041 16163 8075
rect 16313 8041 16347 8075
rect 17969 8041 18003 8075
rect 20269 8041 20303 8075
rect 21925 8041 21959 8075
rect 23029 8041 23063 8075
rect 23673 8041 23707 8075
rect 24225 8041 24259 8075
rect 24777 8041 24811 8075
rect 2145 7973 2179 8007
rect 4169 7973 4203 8007
rect 4261 7973 4295 8007
rect 5641 7973 5675 8007
rect 6371 7973 6405 8007
rect 7297 7973 7331 8007
rect 9873 7973 9907 8007
rect 11437 7973 11471 8007
rect 12909 7973 12943 8007
rect 13001 7973 13035 8007
rect 18153 7973 18187 8007
rect 18429 7973 18463 8007
rect 22471 7973 22505 8007
rect 7757 7905 7791 7939
rect 8217 7905 8251 7939
rect 8953 7905 8987 7939
rect 15761 7905 15795 7939
rect 16497 7905 16531 7939
rect 16681 7905 16715 7939
rect 17049 7905 17083 7939
rect 17601 7905 17635 7939
rect 2053 7837 2087 7871
rect 4445 7837 4479 7871
rect 6009 7837 6043 7871
rect 9781 7837 9815 7871
rect 10057 7837 10091 7871
rect 11345 7837 11379 7871
rect 13185 7837 13219 7871
rect 2605 7769 2639 7803
rect 9413 7769 9447 7803
rect 11897 7769 11931 7803
rect 18521 7905 18555 7939
rect 18981 7905 19015 7939
rect 19349 7905 19383 7939
rect 19717 7905 19751 7939
rect 21132 7905 21166 7939
rect 19993 7837 20027 7871
rect 22109 7837 22143 7871
rect 23857 7837 23891 7871
rect 21235 7769 21269 7803
rect 5181 7701 5215 7735
rect 12725 7701 12759 7735
rect 15117 7701 15151 7735
rect 18153 7701 18187 7735
rect 20729 7701 20763 7735
rect 21557 7701 21591 7735
rect 2789 7497 2823 7531
rect 3157 7497 3191 7531
rect 5181 7497 5215 7531
rect 5871 7497 5905 7531
rect 9045 7497 9079 7531
rect 10149 7497 10183 7531
rect 11897 7497 11931 7531
rect 14565 7497 14599 7531
rect 14841 7497 14875 7531
rect 17417 7497 17451 7531
rect 21189 7497 21223 7531
rect 23029 7497 23063 7531
rect 23213 7497 23247 7531
rect 24961 7497 24995 7531
rect 9781 7429 9815 7463
rect 12173 7429 12207 7463
rect 14289 7429 14323 7463
rect 15577 7429 15611 7463
rect 18245 7429 18279 7463
rect 18889 7429 18923 7463
rect 22569 7429 22603 7463
rect 1869 7361 1903 7395
rect 3617 7361 3651 7395
rect 7389 7361 7423 7395
rect 9229 7361 9263 7395
rect 13829 7361 13863 7395
rect 20545 7361 20579 7395
rect 23213 7361 23247 7395
rect 24041 7361 24075 7395
rect 24317 7361 24351 7395
rect 5768 7293 5802 7327
rect 6193 7293 6227 7327
rect 6929 7293 6963 7327
rect 7297 7293 7331 7327
rect 8217 7293 8251 7327
rect 10701 7293 10735 7327
rect 11437 7293 11471 7327
rect 12633 7293 12667 7327
rect 14381 7293 14415 7327
rect 15945 7293 15979 7327
rect 16129 7293 16163 7327
rect 16497 7293 16531 7327
rect 17049 7293 17083 7327
rect 18061 7293 18095 7327
rect 18521 7293 18555 7327
rect 19073 7293 19107 7327
rect 19533 7293 19567 7327
rect 19901 7293 19935 7327
rect 20269 7293 20303 7327
rect 21373 7293 21407 7327
rect 23397 7293 23431 7327
rect 25513 7293 25547 7327
rect 26065 7293 26099 7327
rect 1777 7225 1811 7259
rect 2231 7225 2265 7259
rect 3525 7225 3559 7259
rect 3979 7225 4013 7259
rect 4905 7225 4939 7259
rect 9321 7225 9355 7259
rect 11529 7225 11563 7259
rect 12954 7225 12988 7259
rect 17785 7225 17819 7259
rect 21694 7225 21728 7259
rect 24133 7225 24167 7259
rect 4537 7157 4571 7191
rect 5641 7157 5675 7191
rect 6653 7157 6687 7191
rect 7849 7157 7883 7191
rect 13553 7157 13587 7191
rect 15761 7157 15795 7191
rect 20913 7157 20947 7191
rect 22293 7157 22327 7191
rect 25697 7157 25731 7191
rect 1869 6953 1903 6987
rect 3617 6953 3651 6987
rect 7665 6953 7699 6987
rect 9137 6953 9171 6987
rect 11713 6953 11747 6987
rect 13369 6953 13403 6987
rect 14381 6953 14415 6987
rect 16405 6953 16439 6987
rect 19073 6953 19107 6987
rect 22109 6953 22143 6987
rect 24041 6953 24075 6987
rect 2145 6885 2179 6919
rect 4261 6885 4295 6919
rect 6187 6885 6221 6919
rect 9873 6885 9907 6919
rect 12541 6885 12575 6919
rect 13093 6885 13127 6919
rect 18705 6885 18739 6919
rect 19993 6885 20027 6919
rect 21281 6885 21315 6919
rect 21833 6885 21867 6919
rect 24317 6885 24351 6919
rect 24409 6885 24443 6919
rect 5825 6817 5859 6851
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 14197 6817 14231 6851
rect 15301 6817 15335 6851
rect 16589 6817 16623 6851
rect 16773 6817 16807 6851
rect 17141 6817 17175 6851
rect 17509 6817 17543 6851
rect 18337 6817 18371 6851
rect 19901 6817 19935 6851
rect 22753 6817 22787 6851
rect 2053 6749 2087 6783
rect 2329 6749 2363 6783
rect 4158 6749 4192 6783
rect 9781 6749 9815 6783
rect 10057 6749 10091 6783
rect 11253 6749 11287 6783
rect 12449 6749 12483 6783
rect 15761 6749 15795 6783
rect 16221 6749 16255 6783
rect 21189 6749 21223 6783
rect 22477 6749 22511 6783
rect 23397 6749 23431 6783
rect 24777 6749 24811 6783
rect 2973 6681 3007 6715
rect 4721 6681 4755 6715
rect 6745 6681 6779 6715
rect 15117 6681 15151 6715
rect 857 6613 891 6647
rect 7021 6613 7055 6647
rect 10793 6613 10827 6647
rect 15485 6613 15519 6647
rect 20269 6613 20303 6647
rect 20637 6613 20671 6647
rect 1685 6409 1719 6443
rect 2053 6409 2087 6443
rect 3341 6409 3375 6443
rect 4905 6409 4939 6443
rect 5549 6409 5583 6443
rect 5917 6409 5951 6443
rect 6285 6409 6319 6443
rect 8217 6409 8251 6443
rect 9781 6409 9815 6443
rect 10057 6409 10091 6443
rect 12633 6409 12667 6443
rect 14105 6409 14139 6443
rect 15485 6409 15519 6443
rect 17325 6409 17359 6443
rect 17785 6409 17819 6443
rect 18889 6409 18923 6443
rect 20821 6409 20855 6443
rect 22753 6409 22787 6443
rect 25145 6409 25179 6443
rect 11805 6341 11839 6375
rect 16221 6341 16255 6375
rect 25513 6341 25547 6375
rect 2421 6273 2455 6307
rect 3065 6273 3099 6307
rect 3985 6273 4019 6307
rect 4261 6273 4295 6307
rect 8861 6273 8895 6307
rect 10701 6273 10735 6307
rect 12909 6273 12943 6307
rect 13277 6273 13311 6307
rect 14565 6273 14599 6307
rect 16405 6273 16439 6307
rect 16773 6273 16807 6307
rect 23857 6273 23891 6307
rect 24501 6273 24535 6307
rect 5733 6205 5767 6239
rect 6837 6205 6871 6239
rect 7297 6205 7331 6239
rect 12173 6205 12207 6239
rect 16313 6205 16347 6239
rect 16589 6205 16623 6239
rect 18061 6205 18095 6239
rect 18521 6205 18555 6239
rect 19073 6205 19107 6239
rect 19533 6205 19567 6239
rect 19993 6205 20027 6239
rect 20269 6205 20303 6239
rect 21465 6205 21499 6239
rect 25329 6205 25363 6239
rect 25881 6205 25915 6239
rect 2513 6137 2547 6171
rect 4077 6137 4111 6171
rect 8769 6137 8803 6171
rect 9223 6137 9257 6171
rect 10793 6137 10827 6171
rect 11345 6137 11379 6171
rect 13001 6137 13035 6171
rect 14473 6137 14507 6171
rect 14927 6137 14961 6171
rect 20545 6137 20579 6171
rect 22109 6137 22143 6171
rect 23489 6137 23523 6171
rect 23949 6137 23983 6171
rect 3709 6069 3743 6103
rect 6653 6069 6687 6103
rect 6929 6069 6963 6103
rect 7941 6069 7975 6103
rect 10425 6069 10459 6103
rect 15853 6069 15887 6103
rect 18245 6069 18279 6103
rect 21281 6069 21315 6103
rect 24777 6069 24811 6103
rect 3433 5865 3467 5899
rect 4445 5865 4479 5899
rect 4721 5865 4755 5899
rect 7205 5865 7239 5899
rect 9137 5865 9171 5899
rect 9505 5865 9539 5899
rect 10241 5865 10275 5899
rect 11897 5865 11931 5899
rect 14565 5865 14599 5899
rect 15761 5865 15795 5899
rect 16405 5865 16439 5899
rect 17049 5865 17083 5899
rect 17693 5865 17727 5899
rect 19993 5865 20027 5899
rect 20361 5865 20395 5899
rect 22569 5865 22603 5899
rect 23121 5865 23155 5899
rect 23857 5865 23891 5899
rect 2605 5797 2639 5831
rect 5635 5797 5669 5831
rect 8211 5797 8245 5831
rect 11339 5797 11373 5831
rect 12449 5797 12483 5831
rect 12909 5797 12943 5831
rect 17325 5797 17359 5831
rect 18061 5797 18095 5831
rect 19717 5797 19751 5831
rect 24317 5797 24351 5831
rect 1444 5729 1478 5763
rect 4261 5729 4295 5763
rect 7849 5729 7883 5763
rect 9724 5729 9758 5763
rect 10977 5729 11011 5763
rect 15301 5729 15335 5763
rect 15577 5729 15611 5763
rect 16865 5729 16899 5763
rect 18245 5729 18279 5763
rect 18705 5729 18739 5763
rect 19073 5729 19107 5763
rect 19441 5729 19475 5763
rect 21097 5729 21131 5763
rect 22201 5729 22235 5763
rect 2513 5661 2547 5695
rect 5273 5661 5307 5695
rect 12633 5661 12667 5695
rect 12817 5661 12851 5695
rect 13093 5661 13127 5695
rect 15393 5661 15427 5695
rect 16681 5661 16715 5695
rect 24225 5661 24259 5695
rect 24501 5661 24535 5695
rect 1547 5593 1581 5627
rect 3065 5593 3099 5627
rect 9827 5593 9861 5627
rect 21281 5593 21315 5627
rect 2145 5525 2179 5559
rect 6193 5525 6227 5559
rect 6837 5525 6871 5559
rect 8769 5525 8803 5559
rect 10517 5525 10551 5559
rect 12633 5525 12667 5559
rect 13737 5525 13771 5559
rect 21833 5525 21867 5559
rect 1593 5321 1627 5355
rect 1961 5321 1995 5355
rect 4077 5321 4111 5355
rect 4445 5321 4479 5355
rect 4721 5321 4755 5355
rect 9689 5321 9723 5355
rect 11529 5321 11563 5355
rect 13461 5321 13495 5355
rect 15393 5321 15427 5355
rect 17417 5321 17451 5355
rect 18245 5321 18279 5355
rect 18797 5321 18831 5355
rect 21097 5321 21131 5355
rect 21741 5321 21775 5355
rect 22753 5321 22787 5355
rect 24041 5321 24075 5355
rect 25237 5321 25271 5355
rect 2145 5185 2179 5219
rect 5825 5253 5859 5287
rect 10793 5253 10827 5287
rect 12173 5253 12207 5287
rect 14657 5253 14691 5287
rect 17785 5253 17819 5287
rect 23029 5253 23063 5287
rect 25605 5253 25639 5287
rect 5273 5185 5307 5219
rect 6193 5185 6227 5219
rect 7205 5185 7239 5219
rect 8401 5185 8435 5219
rect 10241 5185 10275 5219
rect 11253 5185 11287 5219
rect 20453 5185 20487 5219
rect 21833 5185 21867 5219
rect 24777 5185 24811 5219
rect 4169 5117 4203 5151
rect 4445 5117 4479 5151
rect 12449 5117 12483 5151
rect 12909 5117 12943 5151
rect 15669 5117 15703 5151
rect 19073 5117 19107 5151
rect 19717 5117 19751 5151
rect 19993 5117 20027 5151
rect 20177 5117 20211 5151
rect 2466 5049 2500 5083
rect 3341 5049 3375 5083
rect 5365 5049 5399 5083
rect 6929 5049 6963 5083
rect 7021 5049 7055 5083
rect 10333 5049 10367 5083
rect 14105 5049 14139 5083
rect 14197 5049 14231 5083
rect 15577 5049 15611 5083
rect 16957 5049 16991 5083
rect 20729 5049 20763 5083
rect 22154 5049 22188 5083
rect 23489 5049 23523 5083
rect 24317 5049 24351 5083
rect 24409 5049 24443 5083
rect 3065 4981 3099 5015
rect 4353 4981 4387 5015
rect 5089 4981 5123 5015
rect 6653 4981 6687 5015
rect 7941 4981 7975 5015
rect 8309 4981 8343 5015
rect 8769 4981 8803 5015
rect 9321 4981 9355 5015
rect 12541 4981 12575 5015
rect 13921 4981 13955 5015
rect 1547 4777 1581 4811
rect 1961 4777 1995 4811
rect 5273 4777 5307 4811
rect 5549 4777 5583 4811
rect 6929 4777 6963 4811
rect 7849 4777 7883 4811
rect 9045 4777 9079 4811
rect 11345 4777 11379 4811
rect 12909 4777 12943 4811
rect 14105 4777 14139 4811
rect 16405 4777 16439 4811
rect 17693 4777 17727 4811
rect 17969 4777 18003 4811
rect 19901 4777 19935 4811
rect 20637 4777 20671 4811
rect 21281 4777 21315 4811
rect 22201 4777 22235 4811
rect 24133 4777 24167 4811
rect 24685 4777 24719 4811
rect 2329 4709 2363 4743
rect 2605 4709 2639 4743
rect 3157 4709 3191 4743
rect 4158 4709 4192 4743
rect 4270 4709 4304 4743
rect 6095 4709 6129 4743
rect 7573 4709 7607 4743
rect 8125 4709 8159 4743
rect 8217 4709 8251 4743
rect 9873 4709 9907 4743
rect 12449 4709 12483 4743
rect 20361 4709 20395 4743
rect 22753 4709 22787 4743
rect 22845 4709 22879 4743
rect 1476 4641 1510 4675
rect 11253 4641 11287 4675
rect 11713 4641 11747 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 15577 4641 15611 4675
rect 16681 4641 16715 4675
rect 18245 4641 18279 4675
rect 18613 4641 18647 4675
rect 18981 4641 19015 4675
rect 19349 4641 19383 4675
rect 24869 4641 24903 4675
rect 2513 4573 2547 4607
rect 3433 4573 3467 4607
rect 4445 4573 4479 4607
rect 5733 4573 5767 4607
rect 8769 4573 8803 4607
rect 9413 4573 9447 4607
rect 9781 4573 9815 4607
rect 10057 4573 10091 4607
rect 15117 4573 15151 4607
rect 16129 4573 16163 4607
rect 17325 4573 17359 4607
rect 19625 4573 19659 4607
rect 20913 4573 20947 4607
rect 23029 4573 23063 4607
rect 14749 4505 14783 4539
rect 21833 4505 21867 4539
rect 6653 4437 6687 4471
rect 15761 4437 15795 4471
rect 4445 4233 4479 4267
rect 7205 4233 7239 4267
rect 9781 4233 9815 4267
rect 11345 4233 11379 4267
rect 11713 4233 11747 4267
rect 13461 4233 13495 4267
rect 17417 4233 17451 4267
rect 17785 4233 17819 4267
rect 18245 4233 18279 4267
rect 23397 4233 23431 4267
rect 25053 4233 25087 4267
rect 26157 4233 26191 4267
rect 1869 4165 1903 4199
rect 2421 4165 2455 4199
rect 3433 4165 3467 4199
rect 6285 4165 6319 4199
rect 7757 4165 7791 4199
rect 14289 4165 14323 4199
rect 23029 4165 23063 4199
rect 5549 4097 5583 4131
rect 8769 4097 8803 4131
rect 10057 4097 10091 4131
rect 24133 4097 24167 4131
rect 1476 4029 1510 4063
rect 2513 4029 2547 4063
rect 4169 4029 4203 4063
rect 6653 4029 6687 4063
rect 7364 4029 7398 4063
rect 9413 4029 9447 4063
rect 12265 4029 12299 4063
rect 12725 4029 12759 4063
rect 12909 4029 12943 4063
rect 14473 4029 14507 4063
rect 16313 4029 16347 4063
rect 16865 4029 16899 4063
rect 18981 4029 19015 4063
rect 19441 4029 19475 4063
rect 19993 4029 20027 4063
rect 20177 4029 20211 4063
rect 21833 4029 21867 4063
rect 22753 4029 22787 4063
rect 25672 4029 25706 4063
rect 2834 3961 2868 3995
rect 5273 3961 5307 3995
rect 5365 3961 5399 3995
rect 8401 3961 8435 3995
rect 8493 3961 8527 3995
rect 10333 3961 10367 3995
rect 10425 3961 10459 3995
rect 10977 3961 11011 3995
rect 20453 3961 20487 3995
rect 21281 3961 21315 3995
rect 22154 3961 22188 3995
rect 24225 3961 24259 3995
rect 24777 3961 24811 3995
rect 1547 3893 1581 3927
rect 3801 3893 3835 3927
rect 5089 3893 5123 3927
rect 7435 3893 7469 3927
rect 8217 3893 8251 3927
rect 12541 3893 12575 3927
rect 13829 3893 13863 3927
rect 14841 3893 14875 3927
rect 15577 3893 15611 3927
rect 16681 3893 16715 3927
rect 18889 3893 18923 3927
rect 20913 3893 20947 3927
rect 21649 3893 21683 3927
rect 23857 3893 23891 3927
rect 25743 3893 25777 3927
rect 3433 3689 3467 3723
rect 6561 3689 6595 3723
rect 9137 3689 9171 3723
rect 9413 3689 9447 3723
rect 12449 3689 12483 3723
rect 13277 3689 13311 3723
rect 13829 3689 13863 3723
rect 15761 3689 15795 3723
rect 19901 3689 19935 3723
rect 21097 3689 21131 3723
rect 2513 3621 2547 3655
rect 2605 3621 2639 3655
rect 3157 3621 3191 3655
rect 3893 3621 3927 3655
rect 4169 3621 4203 3655
rect 4270 3621 4304 3655
rect 6003 3621 6037 3655
rect 8217 3621 8251 3655
rect 8769 3621 8803 3655
rect 9781 3621 9815 3655
rect 9873 3621 9907 3655
rect 10425 3621 10459 3655
rect 14473 3621 14507 3655
rect 21741 3621 21775 3655
rect 21833 3621 21867 3655
rect 24133 3621 24167 3655
rect 24685 3621 24719 3655
rect 1409 3553 1443 3587
rect 5641 3553 5675 3587
rect 10609 3553 10643 3587
rect 11253 3553 11287 3587
rect 11713 3553 11747 3587
rect 12817 3553 12851 3587
rect 13093 3553 13127 3587
rect 15301 3553 15335 3587
rect 15577 3553 15611 3587
rect 16957 3553 16991 3587
rect 17049 3553 17083 3587
rect 17509 3553 17543 3587
rect 17877 3553 17911 3587
rect 18245 3553 18279 3587
rect 19349 3553 19383 3587
rect 21465 3553 21499 3587
rect 7573 3485 7607 3519
rect 8125 3485 8159 3519
rect 1685 3417 1719 3451
rect 4721 3417 4755 3451
rect 5181 3417 5215 3451
rect 7849 3417 7883 3451
rect 11805 3485 11839 3519
rect 16589 3485 16623 3519
rect 22017 3485 22051 3519
rect 24041 3485 24075 3519
rect 10701 3417 10735 3451
rect 12909 3417 12943 3451
rect 15393 3417 15427 3451
rect 18429 3417 18463 3451
rect 19533 3417 19567 3451
rect 1869 3349 1903 3383
rect 2329 3349 2363 3383
rect 10609 3349 10643 3383
rect 14841 3349 14875 3383
rect 18797 3349 18831 3383
rect 19165 3349 19199 3383
rect 20453 3349 20487 3383
rect 23765 3349 23799 3383
rect 1593 3145 1627 3179
rect 3249 3145 3283 3179
rect 3617 3145 3651 3179
rect 5089 3145 5123 3179
rect 6561 3145 6595 3179
rect 6975 3145 7009 3179
rect 7849 3145 7883 3179
rect 9229 3145 9263 3179
rect 9505 3145 9539 3179
rect 11253 3145 11287 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 21373 3145 21407 3179
rect 22017 3145 22051 3179
rect 23397 3145 23431 3179
rect 2145 3077 2179 3111
rect 4721 3077 4755 3111
rect 5549 3077 5583 3111
rect 6285 3077 6319 3111
rect 8125 3077 8159 3111
rect 11805 3077 11839 3111
rect 14565 3077 14599 3111
rect 14841 3077 14875 3111
rect 19901 3077 19935 3111
rect 2329 3009 2363 3043
rect 2973 3009 3007 3043
rect 8309 3009 8343 3043
rect 10149 3009 10183 3043
rect 10793 3009 10827 3043
rect 15485 3009 15519 3043
rect 17785 3009 17819 3043
rect 19625 3009 19659 3043
rect 20453 3009 20487 3043
rect 21741 3009 21775 3043
rect 24409 3009 24443 3043
rect 24685 3009 24719 3043
rect 3801 2941 3835 2975
rect 5733 2941 5767 2975
rect 6872 2941 6906 2975
rect 12449 2941 12483 2975
rect 12909 2941 12943 2975
rect 14749 2941 14783 2975
rect 15025 2941 15059 2975
rect 18429 2941 18463 2975
rect 18613 2941 18647 2975
rect 18981 2941 19015 2975
rect 19349 2941 19383 2975
rect 22201 2941 22235 2975
rect 22753 2941 22787 2975
rect 23765 2941 23799 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 2421 2873 2455 2907
rect 4122 2873 4156 2907
rect 7297 2873 7331 2907
rect 8630 2873 8664 2907
rect 9873 2873 9907 2907
rect 10241 2873 10275 2907
rect 12173 2873 12207 2907
rect 16129 2873 16163 2907
rect 16486 2873 16520 2907
rect 16589 2873 16623 2907
rect 17141 2873 17175 2907
rect 20774 2873 20808 2907
rect 5917 2805 5951 2839
rect 12541 2805 12575 2839
rect 13553 2805 13587 2839
rect 15853 2805 15887 2839
rect 17417 2805 17451 2839
rect 20269 2805 20303 2839
rect 22385 2805 22419 2839
rect 25421 2805 25455 2839
rect 1593 2601 1627 2635
rect 3433 2601 3467 2635
rect 3801 2601 3835 2635
rect 5089 2601 5123 2635
rect 7067 2601 7101 2635
rect 9229 2601 9263 2635
rect 16129 2601 16163 2635
rect 16589 2601 16623 2635
rect 17693 2601 17727 2635
rect 18153 2601 18187 2635
rect 18705 2601 18739 2635
rect 19533 2601 19567 2635
rect 22661 2601 22695 2635
rect 23765 2601 23799 2635
rect 26157 2601 26191 2635
rect 2237 2533 2271 2567
rect 2605 2533 2639 2567
rect 4261 2533 4295 2567
rect 7757 2533 7791 2567
rect 8262 2533 8296 2567
rect 10057 2533 10091 2567
rect 10425 2533 10459 2567
rect 10977 2533 11011 2567
rect 11345 2533 11379 2567
rect 12633 2533 12667 2567
rect 13829 2533 13863 2567
rect 15209 2533 15243 2567
rect 16865 2533 16899 2567
rect 21005 2533 21039 2567
rect 21373 2533 21407 2567
rect 21925 2533 21959 2567
rect 23673 2533 23707 2567
rect 24133 2533 24167 2567
rect 24225 2533 24259 2567
rect 1409 2465 1443 2499
rect 5825 2465 5859 2499
rect 6285 2465 6319 2499
rect 6996 2465 7030 2499
rect 7389 2465 7423 2499
rect 7941 2465 7975 2499
rect 8861 2465 8895 2499
rect 12725 2465 12759 2499
rect 14289 2465 14323 2499
rect 15577 2465 15611 2499
rect 18337 2465 18371 2499
rect 19901 2465 19935 2499
rect 20152 2465 20186 2499
rect 22845 2465 22879 2499
rect 2513 2397 2547 2431
rect 4169 2397 4203 2431
rect 5457 2397 5491 2431
rect 9597 2397 9631 2431
rect 10333 2397 10367 2431
rect 14197 2397 14231 2431
rect 16773 2397 16807 2431
rect 17141 2397 17175 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 3065 2329 3099 2363
rect 4721 2329 4755 2363
rect 12357 2329 12391 2363
rect 14933 2329 14967 2363
rect 19257 2329 19291 2363
rect 23029 2329 23063 2363
rect 25672 2465 25706 2499
rect 24409 2397 24443 2431
rect 1961 2261 1995 2295
rect 6009 2261 6043 2295
rect 14473 2261 14507 2295
rect 15761 2261 15795 2295
rect 20223 2261 20257 2295
rect 20637 2261 20671 2295
rect 23397 2261 23431 2295
rect 23673 2261 23707 2295
rect 25743 2261 25777 2295
<< metal1 >>
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1578 23848 1584 23860
rect 1539 23820 1584 23848
rect 1578 23808 1584 23820
rect 1636 23808 1642 23860
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 1443 23616 2084 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2056 23517 2084 23616
rect 23474 23604 23480 23656
rect 23532 23644 23538 23656
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 23532 23616 24593 23644
rect 23532 23604 23538 23616
rect 24581 23613 24593 23616
rect 24627 23644 24639 23647
rect 25133 23647 25191 23653
rect 25133 23644 25145 23647
rect 24627 23616 25145 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 25133 23613 25145 23616
rect 25179 23613 25191 23647
rect 25133 23607 25191 23613
rect 2041 23511 2099 23517
rect 2041 23477 2053 23511
rect 2087 23508 2099 23511
rect 2130 23508 2136 23520
rect 2087 23480 2136 23508
rect 2087 23477 2099 23480
rect 2041 23471 2099 23477
rect 2130 23468 2136 23480
rect 2188 23468 2194 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 24762 21672 24768 21684
rect 24723 21644 24768 21672
rect 24762 21632 24768 21644
rect 24820 21632 24826 21684
rect 1118 21428 1124 21480
rect 1176 21468 1182 21480
rect 1397 21471 1455 21477
rect 1397 21468 1409 21471
rect 1176 21440 1409 21468
rect 1176 21428 1182 21440
rect 1397 21437 1409 21440
rect 1443 21468 1455 21471
rect 1949 21471 2007 21477
rect 1949 21468 1961 21471
rect 1443 21440 1961 21468
rect 1443 21437 1455 21440
rect 1397 21431 1455 21437
rect 1949 21437 1961 21440
rect 1995 21437 2007 21471
rect 1949 21431 2007 21437
rect 24026 21428 24032 21480
rect 24084 21468 24090 21480
rect 24581 21471 24639 21477
rect 24581 21468 24593 21471
rect 24084 21440 24593 21468
rect 24084 21428 24090 21440
rect 24581 21437 24593 21440
rect 24627 21468 24639 21471
rect 25133 21471 25191 21477
rect 25133 21468 25145 21471
rect 24627 21440 25145 21468
rect 24627 21437 24639 21440
rect 24581 21431 24639 21437
rect 25133 21437 25145 21440
rect 25179 21437 25191 21471
rect 25133 21431 25191 21437
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1394 20380 1400 20392
rect 1452 20389 1458 20392
rect 1452 20383 1490 20389
rect 1342 20352 1400 20380
rect 1394 20340 1400 20352
rect 1478 20380 1490 20383
rect 1857 20383 1915 20389
rect 1857 20380 1869 20383
rect 1478 20352 1869 20380
rect 1478 20349 1490 20352
rect 1452 20343 1490 20349
rect 1857 20349 1869 20352
rect 1903 20349 1915 20383
rect 1857 20343 1915 20349
rect 1452 20340 1458 20343
rect 937 20247 995 20253
rect 937 20213 949 20247
rect 983 20244 995 20247
rect 1535 20247 1593 20253
rect 1535 20244 1547 20247
rect 983 20216 1547 20244
rect 983 20213 995 20216
rect 937 20207 995 20213
rect 1535 20213 1547 20216
rect 1581 20213 1593 20247
rect 1535 20207 1593 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1302 19864 1308 19916
rect 1360 19904 1366 19916
rect 1432 19907 1490 19913
rect 1432 19904 1444 19907
rect 1360 19876 1444 19904
rect 1360 19864 1366 19876
rect 1432 19873 1444 19876
rect 1478 19904 1490 19907
rect 2222 19904 2228 19916
rect 1478 19876 2228 19904
rect 1478 19873 1490 19876
rect 1432 19867 1490 19873
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 1302 19660 1308 19712
rect 1360 19700 1366 19712
rect 1535 19703 1593 19709
rect 1535 19700 1547 19703
rect 1360 19672 1547 19700
rect 1360 19660 1366 19672
rect 1535 19669 1547 19672
rect 1581 19669 1593 19703
rect 1535 19663 1593 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2222 19496 2228 19508
rect 2183 19468 2228 19496
rect 2222 19456 2228 19468
rect 2280 19456 2286 19508
rect 2038 19388 2044 19440
rect 2096 19428 2102 19440
rect 2547 19431 2605 19437
rect 2547 19428 2559 19431
rect 2096 19400 2559 19428
rect 2096 19388 2102 19400
rect 2547 19397 2559 19400
rect 2593 19397 2605 19431
rect 2547 19391 2605 19397
rect 1464 19295 1522 19301
rect 1464 19261 1476 19295
rect 1510 19292 1522 19295
rect 1854 19292 1860 19304
rect 1510 19264 1860 19292
rect 1510 19261 1522 19264
rect 1464 19255 1522 19261
rect 1854 19252 1860 19264
rect 1912 19252 1918 19304
rect 2476 19295 2534 19301
rect 2476 19261 2488 19295
rect 2522 19292 2534 19295
rect 2522 19264 3004 19292
rect 2522 19261 2534 19264
rect 2476 19255 2534 19261
rect 1535 19159 1593 19165
rect 1535 19125 1547 19159
rect 1581 19156 1593 19159
rect 1946 19156 1952 19168
rect 1581 19128 1952 19156
rect 1581 19125 1593 19128
rect 1535 19119 1593 19125
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 2976 19165 3004 19264
rect 2961 19159 3019 19165
rect 2961 19125 2973 19159
rect 3007 19156 3019 19159
rect 3234 19156 3240 19168
rect 3007 19128 3240 19156
rect 3007 19125 3019 19128
rect 2961 19119 3019 19125
rect 3234 19116 3240 19128
rect 3292 19116 3298 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1210 18776 1216 18828
rect 1268 18816 1274 18828
rect 1432 18819 1490 18825
rect 1432 18816 1444 18819
rect 1268 18788 1444 18816
rect 1268 18776 1274 18788
rect 1432 18785 1444 18788
rect 1478 18785 1490 18819
rect 1432 18779 1490 18785
rect 2222 18776 2228 18828
rect 2280 18816 2286 18828
rect 2444 18819 2502 18825
rect 2444 18816 2456 18819
rect 2280 18788 2456 18816
rect 2280 18776 2286 18788
rect 2444 18785 2456 18788
rect 2490 18785 2502 18819
rect 2444 18779 2502 18785
rect 1535 18615 1593 18621
rect 1535 18581 1547 18615
rect 1581 18612 1593 18615
rect 1762 18612 1768 18624
rect 1581 18584 1768 18612
rect 1581 18581 1593 18584
rect 1535 18575 1593 18581
rect 1762 18572 1768 18584
rect 1820 18572 1826 18624
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2547 18615 2605 18621
rect 2547 18612 2559 18615
rect 2372 18584 2559 18612
rect 2372 18572 2378 18584
rect 2547 18581 2559 18584
rect 2593 18581 2605 18615
rect 2547 18575 2605 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1118 18300 1124 18352
rect 1176 18340 1182 18352
rect 1394 18340 1400 18352
rect 1176 18312 1400 18340
rect 1176 18300 1182 18312
rect 1394 18300 1400 18312
rect 1452 18300 1458 18352
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 1447 18244 2329 18272
rect 934 18164 940 18216
rect 992 18204 998 18216
rect 1447 18213 1475 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 1432 18207 1490 18213
rect 1432 18204 1444 18207
rect 992 18176 1444 18204
rect 992 18164 998 18176
rect 1432 18173 1444 18176
rect 1478 18173 1490 18207
rect 1432 18167 1490 18173
rect 2222 18164 2228 18216
rect 2280 18204 2286 18216
rect 2593 18207 2651 18213
rect 2593 18204 2605 18207
rect 2280 18176 2605 18204
rect 2280 18164 2286 18176
rect 2593 18173 2605 18176
rect 2639 18173 2651 18207
rect 2593 18167 2651 18173
rect 3856 18207 3914 18213
rect 3856 18173 3868 18207
rect 3902 18204 3914 18207
rect 6892 18207 6950 18213
rect 3902 18176 4154 18204
rect 3902 18173 3914 18176
rect 3856 18167 3914 18173
rect 290 18096 296 18148
rect 348 18136 354 18148
rect 1210 18136 1216 18148
rect 348 18108 1216 18136
rect 348 18096 354 18108
rect 1210 18096 1216 18108
rect 1268 18136 1274 18148
rect 1857 18139 1915 18145
rect 1857 18136 1869 18139
rect 1268 18108 1869 18136
rect 1268 18096 1274 18108
rect 1857 18105 1869 18108
rect 1903 18105 1915 18139
rect 4126 18136 4154 18176
rect 6892 18173 6904 18207
rect 6938 18173 6950 18207
rect 6892 18167 6950 18173
rect 4338 18136 4344 18148
rect 4126 18108 4344 18136
rect 1857 18099 1915 18105
rect 4338 18096 4344 18108
rect 4396 18096 4402 18148
rect 6907 18136 6935 18167
rect 7282 18136 7288 18148
rect 6907 18108 7288 18136
rect 7282 18096 7288 18108
rect 7340 18096 7346 18148
rect 1118 18028 1124 18080
rect 1176 18068 1182 18080
rect 1535 18071 1593 18077
rect 1535 18068 1547 18071
rect 1176 18040 1547 18068
rect 1176 18028 1182 18040
rect 1535 18037 1547 18040
rect 1581 18037 1593 18071
rect 2774 18068 2780 18080
rect 2735 18040 2780 18068
rect 1535 18031 1593 18037
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 3927 18071 3985 18077
rect 3927 18068 3939 18071
rect 3476 18040 3939 18068
rect 3476 18028 3482 18040
rect 3927 18037 3939 18040
rect 3973 18037 3985 18071
rect 3927 18031 3985 18037
rect 6822 18028 6828 18080
rect 6880 18068 6886 18080
rect 6963 18071 7021 18077
rect 6963 18068 6975 18071
rect 6880 18040 6975 18068
rect 6880 18028 6886 18040
rect 6963 18037 6975 18040
rect 7009 18037 7021 18071
rect 6963 18031 7021 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1578 17864 1584 17876
rect 1539 17836 1584 17864
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 2314 17728 2320 17740
rect 1443 17700 2320 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 2568 17731 2626 17737
rect 2568 17697 2580 17731
rect 2614 17728 2626 17731
rect 3050 17728 3056 17740
rect 2614 17700 3056 17728
rect 2614 17697 2626 17700
rect 2568 17691 2626 17697
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 3970 17728 3976 17740
rect 3931 17700 3976 17728
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 5144 17731 5202 17737
rect 5144 17697 5156 17731
rect 5190 17728 5202 17731
rect 5258 17728 5264 17740
rect 5190 17700 5264 17728
rect 5190 17697 5202 17700
rect 5144 17691 5202 17697
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 6730 17728 6736 17740
rect 6691 17700 6736 17728
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 13446 17728 13452 17740
rect 13407 17700 13452 17728
rect 13446 17688 13452 17700
rect 13504 17688 13510 17740
rect 13906 17728 13912 17740
rect 13867 17700 13912 17728
rect 13906 17688 13912 17700
rect 13964 17688 13970 17740
rect 15562 17728 15568 17740
rect 15523 17700 15568 17728
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 24581 17731 24639 17737
rect 24581 17697 24593 17731
rect 24627 17728 24639 17731
rect 24670 17728 24676 17740
rect 24627 17700 24676 17728
rect 24627 17697 24639 17700
rect 24581 17691 24639 17697
rect 24670 17688 24676 17700
rect 24728 17688 24734 17740
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 11664 17632 12357 17660
rect 11664 17620 11670 17632
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 12345 17623 12403 17629
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 2639 17527 2697 17533
rect 2639 17493 2651 17527
rect 2685 17524 2697 17527
rect 2958 17524 2964 17536
rect 2685 17496 2964 17524
rect 2685 17493 2697 17496
rect 2639 17487 2697 17493
rect 2958 17484 2964 17496
rect 3016 17484 3022 17536
rect 3786 17484 3792 17536
rect 3844 17524 3850 17536
rect 4203 17527 4261 17533
rect 4203 17524 4215 17527
rect 3844 17496 4215 17524
rect 3844 17484 3850 17496
rect 4203 17493 4215 17496
rect 4249 17493 4261 17527
rect 4203 17487 4261 17493
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 5215 17527 5273 17533
rect 5215 17524 5227 17527
rect 5132 17496 5227 17524
rect 5132 17484 5138 17496
rect 5215 17493 5227 17496
rect 5261 17493 5273 17527
rect 5215 17487 5273 17493
rect 6917 17527 6975 17533
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7190 17524 7196 17536
rect 6963 17496 7196 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 15703 17527 15761 17533
rect 15703 17524 15715 17527
rect 15344 17496 15715 17524
rect 15344 17484 15350 17496
rect 15703 17493 15715 17496
rect 15749 17493 15761 17527
rect 15703 17487 15761 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 2314 17320 2320 17332
rect 2275 17292 2320 17320
rect 2314 17280 2320 17292
rect 2372 17280 2378 17332
rect 2547 17323 2605 17329
rect 2547 17289 2559 17323
rect 2593 17320 2605 17323
rect 8662 17320 8668 17332
rect 2593 17292 8668 17320
rect 2593 17289 2605 17292
rect 2547 17283 2605 17289
rect 8662 17280 8668 17292
rect 8720 17280 8726 17332
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 13446 17320 13452 17332
rect 11020 17292 13452 17320
rect 11020 17280 11026 17292
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 6362 17212 6368 17264
rect 6420 17252 6426 17264
rect 6963 17255 7021 17261
rect 6963 17252 6975 17255
rect 6420 17224 6975 17252
rect 6420 17212 6426 17224
rect 6963 17221 6975 17224
rect 7009 17221 7021 17255
rect 6963 17215 7021 17221
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 9217 17255 9275 17261
rect 9217 17252 9229 17255
rect 8812 17224 9229 17252
rect 8812 17212 8846 17224
rect 9217 17221 9229 17224
rect 9263 17221 9275 17255
rect 9217 17215 9275 17221
rect 10870 17212 10876 17264
rect 10928 17252 10934 17264
rect 11793 17255 11851 17261
rect 11793 17252 11805 17255
rect 10928 17224 11805 17252
rect 10928 17212 10934 17224
rect 11793 17221 11805 17224
rect 11839 17221 11851 17255
rect 11793 17215 11851 17221
rect 3973 17187 4031 17193
rect 3973 17184 3985 17187
rect 3503 17156 3985 17184
rect 106 17076 112 17128
rect 164 17116 170 17128
rect 1432 17119 1490 17125
rect 1432 17116 1444 17119
rect 164 17088 1444 17116
rect 164 17076 170 17088
rect 1432 17085 1444 17088
rect 1478 17116 1490 17119
rect 1857 17119 1915 17125
rect 1857 17116 1869 17119
rect 1478 17088 1869 17116
rect 1478 17085 1490 17088
rect 1432 17079 1490 17085
rect 1857 17085 1869 17088
rect 1903 17085 1915 17119
rect 1857 17079 1915 17085
rect 2476 17119 2534 17125
rect 2476 17085 2488 17119
rect 2522 17116 2534 17119
rect 2866 17116 2872 17128
rect 2522 17088 2872 17116
rect 2522 17085 2534 17088
rect 2476 17079 2534 17085
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 3503 17125 3531 17156
rect 3973 17153 3985 17156
rect 4019 17184 4031 17187
rect 4614 17184 4620 17196
rect 4019 17156 4620 17184
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 8818 17125 8846 17212
rect 11808 17184 11836 17215
rect 12986 17184 12992 17196
rect 11808 17156 12572 17184
rect 12947 17156 12992 17184
rect 3488 17119 3546 17125
rect 3488 17085 3500 17119
rect 3534 17085 3546 17119
rect 3488 17079 3546 17085
rect 4500 17119 4558 17125
rect 4500 17085 4512 17119
rect 4546 17116 4558 17119
rect 5512 17119 5570 17125
rect 4546 17088 4844 17116
rect 4546 17085 4558 17088
rect 4500 17079 4558 17085
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 3970 17048 3976 17060
rect 3200 17020 3976 17048
rect 3200 17008 3206 17020
rect 3970 17008 3976 17020
rect 4028 17048 4034 17060
rect 4249 17051 4307 17057
rect 4249 17048 4261 17051
rect 4028 17020 4261 17048
rect 4028 17008 4034 17020
rect 4249 17017 4261 17020
rect 4295 17017 4307 17051
rect 4249 17011 4307 17017
rect 4816 16992 4844 17088
rect 5512 17085 5524 17119
rect 5558 17116 5570 17119
rect 6892 17119 6950 17125
rect 5558 17088 6040 17116
rect 5558 17085 5570 17088
rect 5512 17079 5570 17085
rect 845 16983 903 16989
rect 845 16949 857 16983
rect 891 16980 903 16983
rect 1535 16983 1593 16989
rect 1535 16980 1547 16983
rect 891 16952 1547 16980
rect 891 16949 903 16952
rect 845 16943 903 16949
rect 1535 16949 1547 16952
rect 1581 16949 1593 16983
rect 1535 16943 1593 16949
rect 3050 16940 3056 16992
rect 3108 16980 3114 16992
rect 3237 16983 3295 16989
rect 3237 16980 3249 16983
rect 3108 16952 3249 16980
rect 3108 16940 3114 16952
rect 3237 16949 3249 16952
rect 3283 16949 3295 16983
rect 3237 16943 3295 16949
rect 3559 16983 3617 16989
rect 3559 16949 3571 16983
rect 3605 16980 3617 16983
rect 3694 16980 3700 16992
rect 3605 16952 3700 16980
rect 3605 16949 3617 16952
rect 3559 16943 3617 16949
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 4571 16983 4629 16989
rect 4571 16949 4583 16983
rect 4617 16980 4629 16983
rect 4706 16980 4712 16992
rect 4617 16952 4712 16980
rect 4617 16949 4629 16952
rect 4571 16943 4629 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4856 16952 4905 16980
rect 4856 16940 4862 16952
rect 4893 16949 4905 16952
rect 4939 16949 4951 16983
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 4893 16943 4951 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 6012 16989 6040 17088
rect 6892 17085 6904 17119
rect 6938 17116 6950 17119
rect 8803 17119 8861 17125
rect 6938 17088 7420 17116
rect 6938 17085 6950 17088
rect 6892 17079 6950 17085
rect 7392 16992 7420 17088
rect 8803 17085 8815 17119
rect 8849 17085 8861 17119
rect 8803 17079 8861 17085
rect 8895 17119 8953 17125
rect 8895 17085 8907 17119
rect 8941 17116 8953 17119
rect 9214 17116 9220 17128
rect 8941 17088 9220 17116
rect 8941 17085 8953 17088
rect 8895 17079 8953 17085
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 10848 17119 10906 17125
rect 10848 17085 10860 17119
rect 10894 17116 10906 17119
rect 11333 17119 11391 17125
rect 11333 17116 11345 17119
rect 10894 17088 11345 17116
rect 10894 17085 10906 17088
rect 10848 17079 10906 17085
rect 11333 17085 11345 17088
rect 11379 17116 11391 17119
rect 11790 17116 11796 17128
rect 11379 17088 11796 17116
rect 11379 17085 11391 17088
rect 11333 17079 11391 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11974 17076 11980 17128
rect 12032 17116 12038 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 12032 17088 12265 17116
rect 12032 17076 12038 17088
rect 12253 17085 12265 17088
rect 12299 17116 12311 17119
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12299 17088 12449 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12544 17116 12572 17156
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 15562 17184 15568 17196
rect 13872 17156 15568 17184
rect 13872 17144 13878 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12544 17088 12909 17116
rect 12437 17079 12495 17085
rect 12897 17085 12909 17088
rect 12943 17116 12955 17119
rect 12943 17088 13814 17116
rect 12943 17085 12955 17088
rect 12897 17079 12955 17085
rect 5583 16983 5641 16989
rect 5583 16980 5595 16983
rect 5408 16952 5595 16980
rect 5408 16940 5414 16952
rect 5583 16949 5595 16952
rect 5629 16949 5641 16983
rect 5583 16943 5641 16949
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 6178 16980 6184 16992
rect 6043 16952 6184 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6178 16940 6184 16952
rect 6236 16940 6242 16992
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 6730 16980 6736 16992
rect 6687 16952 6736 16980
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 7650 16980 7656 16992
rect 7611 16952 7656 16980
rect 7650 16940 7656 16952
rect 7708 16940 7714 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9769 16983 9827 16989
rect 9769 16980 9781 16983
rect 9180 16952 9781 16980
rect 9180 16940 9186 16952
rect 9769 16949 9781 16952
rect 9815 16949 9827 16983
rect 9769 16943 9827 16949
rect 10919 16983 10977 16989
rect 10919 16949 10931 16983
rect 10965 16980 10977 16983
rect 11054 16980 11060 16992
rect 10965 16952 11060 16980
rect 10965 16949 10977 16952
rect 10919 16943 10977 16949
rect 11054 16940 11060 16952
rect 11112 16940 11118 16992
rect 13786 16980 13814 17088
rect 14182 17076 14188 17128
rect 14240 17116 14246 17128
rect 14369 17119 14427 17125
rect 14369 17116 14381 17119
rect 14240 17088 14381 17116
rect 14240 17076 14246 17088
rect 14369 17085 14381 17088
rect 14415 17085 14427 17119
rect 14369 17079 14427 17085
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15013 17079 15071 17085
rect 14277 17051 14335 17057
rect 14277 17017 14289 17051
rect 14323 17048 14335 17051
rect 15028 17048 15056 17079
rect 15654 17076 15660 17128
rect 15712 17116 15718 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15712 17088 15945 17116
rect 15712 17076 15718 17088
rect 15933 17085 15945 17088
rect 15979 17116 15991 17119
rect 16393 17119 16451 17125
rect 16393 17116 16405 17119
rect 15979 17088 16405 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 16393 17085 16405 17088
rect 16439 17085 16451 17119
rect 16393 17079 16451 17085
rect 15838 17048 15844 17060
rect 14323 17020 15844 17048
rect 14323 17017 14335 17020
rect 14277 17011 14335 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 13906 16980 13912 16992
rect 13786 16952 13912 16980
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 16022 16940 16028 16992
rect 16080 16980 16086 16992
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 16080 16952 16129 16980
rect 16080 16940 16086 16952
rect 16117 16949 16129 16952
rect 16163 16949 16175 16983
rect 16117 16943 16175 16949
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 23753 16983 23811 16989
rect 23753 16980 23765 16983
rect 22980 16952 23765 16980
rect 22980 16940 22986 16952
rect 23753 16949 23765 16952
rect 23799 16949 23811 16983
rect 24578 16980 24584 16992
rect 24539 16952 24584 16980
rect 23753 16943 23811 16949
rect 24578 16940 24584 16952
rect 24636 16940 24642 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1026 16736 1032 16788
rect 1084 16776 1090 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1084 16748 1593 16776
rect 1084 16736 1090 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 7742 16776 7748 16788
rect 7703 16748 7748 16776
rect 1581 16739 1639 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16776 13691 16779
rect 13722 16776 13728 16788
rect 13679 16748 13728 16776
rect 13679 16745 13691 16748
rect 13633 16739 13691 16745
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 23707 16779 23765 16785
rect 23707 16745 23719 16779
rect 23753 16776 23765 16779
rect 24578 16776 24584 16788
rect 23753 16748 24584 16776
rect 23753 16745 23765 16748
rect 23707 16739 23765 16745
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 6178 16708 6184 16720
rect 1412 16680 6184 16708
rect 1412 16649 1440 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 1397 16643 1455 16649
rect 1397 16609 1409 16643
rect 1443 16640 1455 16643
rect 1578 16640 1584 16652
rect 1443 16612 1584 16640
rect 1443 16609 1455 16612
rect 1397 16603 1455 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2501 16643 2559 16649
rect 2501 16609 2513 16643
rect 2547 16640 2559 16643
rect 2590 16640 2596 16652
rect 2547 16612 2596 16640
rect 2547 16609 2559 16612
rect 2501 16603 2559 16609
rect 2590 16600 2596 16612
rect 2648 16600 2654 16652
rect 4132 16643 4190 16649
rect 4132 16609 4144 16643
rect 4178 16640 4190 16643
rect 4430 16640 4436 16652
rect 4178 16612 4436 16640
rect 4178 16609 4190 16612
rect 4132 16603 4190 16609
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 6270 16640 6276 16652
rect 5675 16612 6276 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 6270 16600 6276 16612
rect 6328 16600 6334 16652
rect 6708 16643 6766 16649
rect 6708 16609 6720 16643
rect 6754 16640 6766 16643
rect 7098 16640 7104 16652
rect 6754 16612 7104 16640
rect 6754 16609 6766 16612
rect 6708 16603 6766 16609
rect 7098 16600 7104 16612
rect 7156 16600 7162 16652
rect 7834 16640 7840 16652
rect 7795 16612 7840 16640
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 7650 16572 7656 16584
rect 7484 16544 7656 16572
rect 5994 16464 6000 16516
rect 6052 16504 6058 16516
rect 6779 16507 6837 16513
rect 6779 16504 6791 16507
rect 6052 16476 6791 16504
rect 6052 16464 6058 16476
rect 6779 16473 6791 16476
rect 6825 16473 6837 16507
rect 6779 16467 6837 16473
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 2639 16439 2697 16445
rect 2639 16436 2651 16439
rect 2556 16408 2651 16436
rect 2556 16396 2562 16408
rect 2639 16405 2651 16408
rect 2685 16405 2697 16439
rect 2639 16399 2697 16405
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 4203 16439 4261 16445
rect 4203 16436 4215 16439
rect 3384 16408 4215 16436
rect 3384 16396 3390 16408
rect 4203 16405 4215 16408
rect 4249 16405 4261 16439
rect 4203 16399 4261 16405
rect 5813 16439 5871 16445
rect 5813 16405 5825 16439
rect 5859 16436 5871 16439
rect 6086 16436 6092 16448
rect 5859 16408 6092 16436
rect 5859 16405 5871 16408
rect 5813 16399 5871 16405
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 7484 16445 7512 16544
rect 7650 16532 7656 16544
rect 7708 16572 7714 16584
rect 8128 16572 8156 16603
rect 8202 16572 8208 16584
rect 7708 16544 8208 16572
rect 7708 16532 7714 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 9692 16572 9720 16603
rect 9766 16600 9772 16652
rect 9824 16640 9830 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9824 16612 10149 16640
rect 9824 16600 9830 16612
rect 10137 16609 10149 16612
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 12710 16640 12716 16652
rect 12667 16612 12716 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 13630 16640 13636 16652
rect 13591 16612 13636 16640
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13964 16612 14105 16640
rect 13964 16600 13970 16612
rect 14093 16609 14105 16612
rect 14139 16640 14151 16643
rect 14274 16640 14280 16652
rect 14139 16612 14280 16640
rect 14139 16609 14151 16612
rect 14093 16603 14151 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15378 16640 15384 16652
rect 15335 16612 15384 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 15470 16600 15476 16652
rect 15528 16640 15534 16652
rect 15565 16643 15623 16649
rect 15565 16640 15577 16643
rect 15528 16612 15577 16640
rect 15528 16600 15534 16612
rect 15565 16609 15577 16612
rect 15611 16609 15623 16643
rect 16850 16640 16856 16652
rect 16811 16612 16856 16640
rect 15565 16603 15623 16609
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 23477 16643 23535 16649
rect 23477 16609 23489 16643
rect 23523 16640 23535 16643
rect 23566 16640 23572 16652
rect 23523 16612 23572 16640
rect 23523 16609 23535 16612
rect 23477 16603 23535 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 24648 16643 24706 16649
rect 24648 16609 24660 16643
rect 24694 16640 24706 16643
rect 24762 16640 24768 16652
rect 24694 16612 24768 16640
rect 24694 16609 24706 16612
rect 24648 16603 24706 16609
rect 24762 16600 24768 16612
rect 24820 16600 24826 16652
rect 10042 16572 10048 16584
rect 9692 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 14608 16544 15761 16572
rect 14608 16532 14614 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20864 16544 20913 16572
rect 20864 16532 20870 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 14182 16464 14188 16516
rect 14240 16504 14246 16516
rect 15381 16507 15439 16513
rect 15381 16504 15393 16507
rect 14240 16476 15393 16504
rect 14240 16464 14246 16476
rect 15381 16473 15393 16476
rect 15427 16504 15439 16507
rect 16666 16504 16672 16516
rect 15427 16476 16672 16504
rect 15427 16473 15439 16476
rect 15381 16467 15439 16473
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 24719 16507 24777 16513
rect 24719 16504 24731 16507
rect 23446 16476 24731 16504
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 6696 16408 7481 16436
rect 6696 16396 6702 16408
rect 7469 16405 7481 16408
rect 7515 16405 7527 16439
rect 10870 16436 10876 16448
rect 10831 16408 10876 16436
rect 7469 16399 7527 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 12250 16436 12256 16448
rect 12211 16408 12256 16436
rect 12250 16396 12256 16408
rect 12308 16436 12314 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12308 16408 13001 16436
rect 12308 16396 12314 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 17034 16436 17040 16448
rect 16995 16408 17040 16436
rect 12989 16399 13047 16405
rect 17034 16396 17040 16408
rect 17092 16396 17098 16448
rect 18598 16396 18604 16448
rect 18656 16436 18662 16448
rect 23446 16436 23474 16476
rect 24719 16473 24731 16476
rect 24765 16473 24777 16507
rect 24719 16467 24777 16473
rect 18656 16408 23474 16436
rect 18656 16396 18662 16408
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1486 16192 1492 16244
rect 1544 16232 1550 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1544 16204 1593 16232
rect 1544 16192 1550 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 4663 16235 4721 16241
rect 4663 16232 4675 16235
rect 2188 16204 4675 16232
rect 2188 16192 2194 16204
rect 4663 16201 4675 16204
rect 4709 16201 4721 16235
rect 4663 16195 4721 16201
rect 8757 16235 8815 16241
rect 8757 16201 8769 16235
rect 8803 16232 8815 16235
rect 11974 16232 11980 16244
rect 8803 16204 11980 16232
rect 8803 16201 8815 16204
rect 8757 16195 8815 16201
rect 2041 16167 2099 16173
rect 2041 16133 2053 16167
rect 2087 16164 2099 16167
rect 4154 16164 4160 16176
rect 2087 16136 4160 16164
rect 2087 16133 2099 16136
rect 2041 16127 2099 16133
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 2056 16028 2084 16127
rect 4154 16124 4160 16136
rect 4212 16124 4218 16176
rect 8772 16164 8800 16195
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 12124 16204 13737 16232
rect 12124 16192 12130 16204
rect 13725 16201 13737 16204
rect 13771 16232 13783 16235
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13771 16204 13829 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 13817 16195 13875 16201
rect 15378 16192 15384 16244
rect 15436 16232 15442 16244
rect 16114 16232 16120 16244
rect 15436 16204 16120 16232
rect 15436 16192 15442 16204
rect 16114 16192 16120 16204
rect 16172 16232 16178 16244
rect 16301 16235 16359 16241
rect 16301 16232 16313 16235
rect 16172 16204 16313 16232
rect 16172 16192 16178 16204
rect 16301 16201 16313 16204
rect 16347 16201 16359 16235
rect 16666 16232 16672 16244
rect 16627 16204 16672 16232
rect 16301 16195 16359 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 24581 16235 24639 16241
rect 24581 16201 24593 16235
rect 24627 16232 24639 16235
rect 24762 16232 24768 16244
rect 24627 16204 24768 16232
rect 24627 16201 24639 16204
rect 24581 16195 24639 16201
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25222 16232 25228 16244
rect 25183 16204 25228 16232
rect 25222 16192 25228 16204
rect 25280 16192 25286 16244
rect 8036 16136 8800 16164
rect 11885 16167 11943 16173
rect 6270 16096 6276 16108
rect 6231 16068 6276 16096
rect 6270 16056 6276 16068
rect 6328 16056 6334 16108
rect 1443 16000 2084 16028
rect 2547 16031 2605 16037
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2547 15997 2559 16031
rect 2593 15997 2605 16031
rect 2547 15991 2605 15997
rect 1486 15920 1492 15972
rect 1544 15960 1550 15972
rect 2562 15960 2590 15991
rect 2682 15988 2688 16040
rect 2740 16028 2746 16040
rect 2961 16031 3019 16037
rect 2961 16028 2973 16031
rect 2740 16000 2973 16028
rect 2740 15988 2746 16000
rect 2961 15997 2973 16000
rect 3007 15997 3019 16031
rect 2961 15991 3019 15997
rect 3580 16031 3638 16037
rect 3580 15997 3592 16031
rect 3626 16028 3638 16031
rect 3626 16000 4016 16028
rect 3626 15997 3638 16000
rect 3580 15991 3638 15997
rect 3988 15972 4016 16000
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4592 16031 4650 16037
rect 4592 16028 4604 16031
rect 4396 16000 4604 16028
rect 4396 15988 4402 16000
rect 4592 15997 4604 16000
rect 4638 16028 4650 16031
rect 4985 16031 5043 16037
rect 4985 16028 4997 16031
rect 4638 16000 4997 16028
rect 4638 15997 4650 16000
rect 4592 15991 4650 15997
rect 4985 15997 4997 16000
rect 5031 15997 5043 16031
rect 4985 15991 5043 15997
rect 5721 16031 5779 16037
rect 5721 15997 5733 16031
rect 5767 16028 5779 16031
rect 5767 16000 6592 16028
rect 5767 15997 5779 16000
rect 5721 15991 5779 15997
rect 3329 15963 3387 15969
rect 3329 15960 3341 15963
rect 1544 15932 3341 15960
rect 1544 15920 1550 15932
rect 3329 15929 3341 15932
rect 3375 15929 3387 15963
rect 3970 15960 3976 15972
rect 3931 15932 3976 15960
rect 3329 15923 3387 15929
rect 3970 15920 3976 15932
rect 4028 15920 4034 15972
rect 6564 15904 6592 16000
rect 7466 15988 7472 16040
rect 7524 16028 7530 16040
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 7524 16000 7941 16028
rect 7524 15988 7530 16000
rect 7929 15997 7941 16000
rect 7975 16028 7987 16031
rect 8036 16028 8064 16136
rect 11885 16133 11897 16167
rect 11931 16164 11943 16167
rect 12710 16164 12716 16176
rect 11931 16136 12716 16164
rect 11931 16133 11943 16136
rect 11885 16127 11943 16133
rect 12710 16124 12716 16136
rect 12768 16124 12774 16176
rect 17129 16167 17187 16173
rect 17129 16133 17141 16167
rect 17175 16164 17187 16167
rect 17586 16164 17592 16176
rect 17175 16136 17592 16164
rect 17175 16133 17187 16136
rect 17129 16127 17187 16133
rect 17586 16124 17592 16136
rect 17644 16124 17650 16176
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 23566 16164 23572 16176
rect 22060 16136 23572 16164
rect 22060 16124 22066 16136
rect 23566 16124 23572 16136
rect 23624 16164 23630 16176
rect 24121 16167 24179 16173
rect 24121 16164 24133 16167
rect 23624 16136 24133 16164
rect 23624 16124 23630 16136
rect 24121 16133 24133 16136
rect 24167 16133 24179 16167
rect 24121 16127 24179 16133
rect 8312 16068 9812 16096
rect 7975 16000 8064 16028
rect 8113 16031 8171 16037
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 8113 15997 8125 16031
rect 8159 16028 8171 16031
rect 8202 16028 8208 16040
rect 8159 16000 8208 16028
rect 8159 15997 8171 16000
rect 8113 15991 8171 15997
rect 8202 15988 8208 16000
rect 8260 16028 8266 16040
rect 8312 16028 8340 16068
rect 9784 16040 9812 16068
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 12308 16068 12541 16096
rect 12308 16056 12314 16068
rect 12529 16065 12541 16068
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 13587 16068 14780 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 8260 16000 8340 16028
rect 8260 15988 8266 16000
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8444 16000 9137 16028
rect 8444 15988 8450 16000
rect 9125 15997 9137 16000
rect 9171 16028 9183 16031
rect 9217 16031 9275 16037
rect 9217 16028 9229 16031
rect 9171 16000 9229 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 9217 15997 9229 16000
rect 9263 15997 9275 16031
rect 9766 16028 9772 16040
rect 9727 16000 9772 16028
rect 9217 15991 9275 15997
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10781 16031 10839 16037
rect 10781 16028 10793 16031
rect 10735 16000 10793 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10781 15997 10793 16000
rect 10827 15997 10839 16031
rect 10781 15991 10839 15997
rect 7561 15963 7619 15969
rect 7561 15929 7573 15963
rect 7607 15960 7619 15963
rect 7834 15960 7840 15972
rect 7607 15932 7840 15960
rect 7607 15929 7619 15932
rect 7561 15923 7619 15929
rect 7834 15920 7840 15932
rect 7892 15960 7898 15972
rect 8294 15960 8300 15972
rect 7892 15932 8300 15960
rect 7892 15920 7898 15932
rect 8294 15920 8300 15932
rect 8352 15960 8358 15972
rect 10704 15960 10732 15991
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 10928 16000 11253 16028
rect 10928 15988 10934 16000
rect 11241 15997 11253 16000
rect 11287 15997 11299 16031
rect 11241 15991 11299 15997
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 11514 15960 11520 15972
rect 8352 15932 10732 15960
rect 11475 15932 11520 15960
rect 8352 15920 8358 15932
rect 11514 15920 11520 15932
rect 11572 15920 11578 15972
rect 12452 15960 12480 15991
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12676 16000 12725 16028
rect 12676 15988 12682 16000
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 13556 16028 13584 16059
rect 12713 15991 12771 15997
rect 12820 16000 13584 16028
rect 13725 16031 13783 16037
rect 12820 15960 12848 16000
rect 13725 15997 13737 16031
rect 13771 16028 13783 16031
rect 14036 16031 14094 16037
rect 14036 16028 14048 16031
rect 13771 16000 14048 16028
rect 13771 15997 13783 16000
rect 13725 15991 13783 15997
rect 14036 15997 14048 16000
rect 14082 15997 14094 16031
rect 14036 15991 14094 15997
rect 12452 15932 12848 15960
rect 12894 15920 12900 15972
rect 12952 15960 12958 15972
rect 14139 15963 14197 15969
rect 14139 15960 14151 15963
rect 12952 15932 14151 15960
rect 12952 15920 12958 15932
rect 14139 15929 14151 15932
rect 14185 15929 14197 15963
rect 14752 15960 14780 16068
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 15252 16068 15301 16096
rect 15252 16056 15258 16068
rect 15289 16065 15301 16068
rect 15335 16096 15347 16099
rect 15335 16068 16988 16096
rect 15335 16065 15347 16068
rect 15289 16059 15347 16065
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 16028 14887 16031
rect 15838 16028 15844 16040
rect 14875 16000 15844 16028
rect 14875 15997 14887 16000
rect 14829 15991 14887 15997
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 16960 16037 16988 16068
rect 22738 16056 22744 16108
rect 22796 16096 22802 16108
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22796 16068 23029 16096
rect 22796 16056 22802 16068
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 16945 16031 17003 16037
rect 16945 15997 16957 16031
rect 16991 16028 17003 16031
rect 17773 16031 17831 16037
rect 17773 16028 17785 16031
rect 16991 16000 17785 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17773 15997 17785 16000
rect 17819 15997 17831 16031
rect 18046 16028 18052 16040
rect 17959 16000 18052 16028
rect 17773 15991 17831 15997
rect 18046 15988 18052 16000
rect 18104 16028 18110 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18104 16000 18521 16028
rect 18104 15988 18110 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 22608 16031 22666 16037
rect 22608 15997 22620 16031
rect 22654 16028 22666 16031
rect 22756 16028 22784 16056
rect 22654 16000 22784 16028
rect 24740 16031 24798 16037
rect 22654 15997 22666 16000
rect 22608 15991 22666 15997
rect 24740 15997 24752 16031
rect 24786 16028 24798 16031
rect 25222 16028 25228 16040
rect 24786 16000 25228 16028
rect 24786 15997 24798 16000
rect 24740 15991 24798 15997
rect 25222 15988 25228 16000
rect 25280 15988 25286 16040
rect 18414 15960 18420 15972
rect 14752 15932 18420 15960
rect 14139 15923 14197 15929
rect 18414 15920 18420 15932
rect 18472 15920 18478 15972
rect 22695 15963 22753 15969
rect 22695 15929 22707 15963
rect 22741 15960 22753 15963
rect 23106 15960 23112 15972
rect 22741 15932 23112 15960
rect 22741 15929 22753 15932
rect 22695 15923 22753 15929
rect 23106 15920 23112 15932
rect 23164 15920 23170 15972
rect 2406 15852 2412 15904
rect 2464 15892 2470 15904
rect 2639 15895 2697 15901
rect 2639 15892 2651 15895
rect 2464 15864 2651 15892
rect 2464 15852 2470 15864
rect 2639 15861 2651 15864
rect 2685 15861 2697 15895
rect 2639 15855 2697 15861
rect 3651 15895 3709 15901
rect 3651 15861 3663 15895
rect 3697 15892 3709 15895
rect 3878 15892 3884 15904
rect 3697 15864 3884 15892
rect 3697 15861 3709 15864
rect 3651 15855 3709 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4430 15892 4436 15904
rect 4391 15864 4436 15892
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 5905 15895 5963 15901
rect 5905 15892 5917 15895
rect 5592 15864 5917 15892
rect 5592 15852 5598 15864
rect 5905 15861 5917 15864
rect 5951 15861 5963 15895
rect 6546 15892 6552 15904
rect 6507 15864 6552 15892
rect 5905 15855 5963 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 8018 15892 8024 15904
rect 7975 15864 8024 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 8018 15852 8024 15864
rect 8076 15852 8082 15904
rect 9306 15892 9312 15904
rect 9267 15864 9312 15892
rect 9306 15852 9312 15864
rect 9364 15852 9370 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 10100 15864 10241 15892
rect 10100 15852 10106 15864
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 10229 15855 10287 15861
rect 12253 15895 12311 15901
rect 12253 15861 12265 15895
rect 12299 15892 12311 15895
rect 12434 15892 12440 15904
rect 12299 15864 12440 15892
rect 12299 15861 12311 15864
rect 12253 15855 12311 15861
rect 12434 15852 12440 15864
rect 12492 15852 12498 15904
rect 13265 15895 13323 15901
rect 13265 15861 13277 15895
rect 13311 15892 13323 15895
rect 13538 15892 13544 15904
rect 13311 15864 13544 15892
rect 13311 15861 13323 15864
rect 13265 15855 13323 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15470 15892 15476 15904
rect 15243 15864 15476 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17405 15895 17463 15901
rect 17405 15892 17417 15895
rect 16908 15864 17417 15892
rect 16908 15852 16914 15864
rect 17405 15861 17417 15864
rect 17451 15861 17463 15895
rect 17405 15855 17463 15861
rect 18138 15852 18144 15904
rect 18196 15892 18202 15904
rect 18233 15895 18291 15901
rect 18233 15892 18245 15895
rect 18196 15864 18245 15892
rect 18196 15852 18202 15864
rect 18233 15861 18245 15864
rect 18279 15861 18291 15895
rect 18233 15855 18291 15861
rect 21085 15895 21143 15901
rect 21085 15861 21097 15895
rect 21131 15892 21143 15895
rect 21726 15892 21732 15904
rect 21131 15864 21732 15892
rect 21131 15861 21143 15864
rect 21085 15855 21143 15861
rect 21726 15852 21732 15864
rect 21784 15852 21790 15904
rect 22462 15852 22468 15904
rect 22520 15892 22526 15904
rect 23661 15895 23719 15901
rect 23661 15892 23673 15895
rect 22520 15864 23673 15892
rect 22520 15852 22526 15864
rect 23661 15861 23673 15864
rect 23707 15861 23719 15895
rect 23661 15855 23719 15861
rect 24811 15895 24869 15901
rect 24811 15861 24823 15895
rect 24857 15892 24869 15895
rect 24946 15892 24952 15904
rect 24857 15864 24952 15892
rect 24857 15861 24869 15864
rect 24811 15855 24869 15861
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 7561 15691 7619 15697
rect 2096 15660 4154 15688
rect 2096 15648 2102 15660
rect 14 15580 20 15632
rect 72 15620 78 15632
rect 2682 15620 2688 15632
rect 72 15592 2688 15620
rect 72 15580 78 15592
rect 2682 15580 2688 15592
rect 2740 15580 2746 15632
rect 4126 15620 4154 15660
rect 7561 15657 7573 15691
rect 7607 15688 7619 15691
rect 7926 15688 7932 15700
rect 7607 15660 7932 15688
rect 7607 15657 7619 15660
rect 7561 15651 7619 15657
rect 7576 15620 7604 15651
rect 7926 15648 7932 15660
rect 7984 15688 7990 15700
rect 13630 15688 13636 15700
rect 7984 15660 13636 15688
rect 7984 15648 7990 15660
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 4126 15592 7604 15620
rect 9309 15623 9367 15629
rect 2038 15552 2044 15564
rect 1999 15524 2044 15552
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 2777 15555 2835 15561
rect 2777 15552 2789 15555
rect 2271 15524 2789 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 2777 15521 2789 15524
rect 2823 15552 2835 15555
rect 2866 15552 2872 15564
rect 2823 15524 2872 15552
rect 2823 15521 2835 15524
rect 2777 15515 2835 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 4132 15555 4190 15561
rect 4132 15521 4144 15555
rect 4178 15552 4190 15555
rect 4246 15552 4252 15564
rect 4178 15524 4252 15552
rect 4178 15521 4190 15524
rect 4132 15515 4190 15521
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4890 15512 4896 15564
rect 4948 15552 4954 15564
rect 5112 15555 5170 15561
rect 5112 15552 5124 15555
rect 4948 15524 5124 15552
rect 4948 15512 4954 15524
rect 5112 15521 5124 15524
rect 5158 15521 5170 15555
rect 5112 15515 5170 15521
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 6564 15561 6592 15592
rect 9309 15589 9321 15623
rect 9355 15620 9367 15623
rect 9766 15620 9772 15632
rect 9355 15592 9772 15620
rect 9355 15589 9367 15592
rect 9309 15583 9367 15589
rect 9766 15580 9772 15592
rect 9824 15620 9830 15632
rect 9953 15623 10011 15629
rect 9953 15620 9965 15623
rect 9824 15592 9965 15620
rect 9824 15580 9830 15592
rect 9953 15589 9965 15592
rect 9999 15620 10011 15623
rect 14274 15620 14280 15632
rect 9999 15592 11100 15620
rect 14187 15592 14280 15620
rect 9999 15589 10011 15592
rect 9953 15583 10011 15589
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 6512 15524 6561 15552
rect 6512 15512 6518 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6549 15515 6607 15521
rect 6638 15512 6644 15564
rect 6696 15552 6702 15564
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6696 15524 6745 15552
rect 6696 15512 6702 15524
rect 6733 15521 6745 15524
rect 6779 15521 6791 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 6733 15515 6791 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 8386 15552 8392 15564
rect 8347 15524 8392 15552
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 10962 15552 10968 15564
rect 10919 15524 10968 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11072 15561 11100 15592
rect 14274 15580 14280 15592
rect 14332 15620 14338 15632
rect 18230 15620 18236 15632
rect 14332 15592 18236 15620
rect 14332 15580 14338 15592
rect 18230 15580 18236 15592
rect 18288 15580 18294 15632
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11698 15552 11704 15564
rect 11103 15524 11704 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15552 12219 15555
rect 12342 15552 12348 15564
rect 12207 15524 12348 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 12492 15524 12537 15552
rect 12492 15512 12498 15524
rect 13078 15512 13084 15564
rect 13136 15552 13142 15564
rect 13760 15555 13818 15561
rect 13760 15552 13772 15555
rect 13136 15524 13772 15552
rect 13136 15512 13142 15524
rect 13760 15521 13772 15524
rect 13806 15521 13818 15555
rect 13760 15515 13818 15521
rect 15289 15555 15347 15561
rect 15289 15521 15301 15555
rect 15335 15552 15347 15555
rect 15378 15552 15384 15564
rect 15335 15524 15384 15552
rect 15335 15521 15347 15524
rect 15289 15515 15347 15521
rect 15378 15512 15384 15524
rect 15436 15512 15442 15564
rect 15565 15555 15623 15561
rect 15565 15521 15577 15555
rect 15611 15521 15623 15555
rect 17218 15552 17224 15564
rect 17179 15524 17224 15552
rect 15565 15515 15623 15521
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 3050 15484 3056 15496
rect 2562 15456 3056 15484
rect 1486 15376 1492 15428
rect 1544 15416 1550 15428
rect 2562 15416 2590 15456
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 7006 15484 7012 15496
rect 6967 15456 7012 15484
rect 7006 15444 7012 15456
rect 7064 15444 7070 15496
rect 8570 15484 8576 15496
rect 8531 15456 8576 15484
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 12621 15487 12679 15493
rect 12621 15484 12633 15487
rect 11296 15456 12633 15484
rect 11296 15444 11302 15456
rect 12621 15453 12633 15456
rect 12667 15453 12679 15487
rect 12621 15447 12679 15453
rect 15105 15487 15163 15493
rect 15105 15453 15117 15487
rect 15151 15484 15163 15487
rect 15580 15484 15608 15515
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 18414 15552 18420 15564
rect 18375 15524 18420 15552
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 20968 15555 21026 15561
rect 20968 15521 20980 15555
rect 21014 15552 21026 15555
rect 22094 15552 22100 15564
rect 21014 15524 22100 15552
rect 21014 15521 21026 15524
rect 20968 15515 21026 15521
rect 22094 15512 22100 15524
rect 22152 15512 22158 15564
rect 23290 15512 23296 15564
rect 23348 15552 23354 15564
rect 23696 15555 23754 15561
rect 23696 15552 23708 15555
rect 23348 15524 23708 15552
rect 23348 15512 23354 15524
rect 23696 15521 23708 15524
rect 23742 15521 23754 15555
rect 23696 15515 23754 15521
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 15151 15456 16865 15484
rect 15151 15453 15163 15456
rect 15105 15447 15163 15453
rect 16853 15453 16865 15456
rect 16899 15484 16911 15487
rect 17770 15484 17776 15496
rect 16899 15456 17776 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19429 15487 19487 15493
rect 19429 15484 19441 15487
rect 19392 15456 19441 15484
rect 19392 15444 19398 15456
rect 19429 15453 19441 15456
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 21634 15444 21640 15496
rect 21692 15484 21698 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21692 15456 21925 15484
rect 21692 15444 21698 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 24673 15487 24731 15493
rect 24673 15453 24685 15487
rect 24719 15484 24731 15487
rect 25314 15484 25320 15496
rect 24719 15456 25320 15484
rect 24719 15453 24731 15456
rect 24673 15447 24731 15453
rect 25314 15444 25320 15456
rect 25372 15444 25378 15496
rect 1544 15388 2590 15416
rect 1544 15376 1550 15388
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 5215 15419 5273 15425
rect 5215 15416 5227 15419
rect 4120 15388 5227 15416
rect 4120 15376 4126 15388
rect 5215 15385 5227 15388
rect 5261 15385 5273 15419
rect 12250 15416 12256 15428
rect 12211 15388 12256 15416
rect 5215 15379 5273 15385
rect 12250 15376 12256 15388
rect 12308 15376 12314 15428
rect 13863 15419 13921 15425
rect 13863 15385 13875 15419
rect 13909 15416 13921 15419
rect 14274 15416 14280 15428
rect 13909 15388 14280 15416
rect 13909 15385 13921 15388
rect 13863 15379 13921 15385
rect 14274 15376 14280 15388
rect 14332 15376 14338 15428
rect 14366 15376 14372 15428
rect 14424 15416 14430 15428
rect 15194 15416 15200 15428
rect 14424 15388 15200 15416
rect 14424 15376 14430 15388
rect 15194 15376 15200 15388
rect 15252 15416 15258 15428
rect 15381 15419 15439 15425
rect 15381 15416 15393 15419
rect 15252 15388 15393 15416
rect 15252 15376 15258 15388
rect 15381 15385 15393 15388
rect 15427 15385 15439 15419
rect 15381 15379 15439 15385
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 4203 15351 4261 15357
rect 4203 15348 4215 15351
rect 3108 15320 4215 15348
rect 3108 15308 3114 15320
rect 4203 15317 4215 15320
rect 4249 15317 4261 15351
rect 5534 15348 5540 15360
rect 5495 15320 5540 15348
rect 4203 15311 4261 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 15562 15308 15568 15360
rect 15620 15348 15626 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 15620 15320 16313 15348
rect 15620 15308 15626 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16301 15311 16359 15317
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 18782 15348 18788 15360
rect 18647 15320 18788 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 21039 15351 21097 15357
rect 21039 15317 21051 15351
rect 21085 15348 21097 15351
rect 21174 15348 21180 15360
rect 21085 15320 21180 15348
rect 21085 15317 21097 15320
rect 21039 15311 21097 15317
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 23799 15351 23857 15357
rect 23799 15317 23811 15351
rect 23845 15348 23857 15351
rect 24762 15348 24768 15360
rect 23845 15320 24768 15348
rect 23845 15317 23857 15320
rect 23799 15311 23857 15317
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 2961 15147 3019 15153
rect 2961 15144 2973 15147
rect 2924 15116 2973 15144
rect 2924 15104 2930 15116
rect 2961 15113 2973 15116
rect 3007 15113 3019 15147
rect 2961 15107 3019 15113
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 6454 15144 6460 15156
rect 6411 15116 6460 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 10229 15147 10287 15153
rect 10229 15113 10241 15147
rect 10275 15144 10287 15147
rect 10962 15144 10968 15156
rect 10275 15116 10968 15144
rect 10275 15113 10287 15116
rect 10229 15107 10287 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 14700 15116 22293 15144
rect 14700 15104 14706 15116
rect 7558 15076 7564 15088
rect 2240 15048 7564 15076
rect 2240 14949 2268 15048
rect 7558 15036 7564 15048
rect 7616 15076 7622 15088
rect 8849 15079 8907 15085
rect 8849 15076 8861 15079
rect 7616 15048 8861 15076
rect 7616 15036 7622 15048
rect 8849 15045 8861 15048
rect 8895 15076 8907 15079
rect 10042 15076 10048 15088
rect 8895 15048 10048 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 2884 14980 5672 15008
rect 2884 14952 2912 14980
rect 1857 14943 1915 14949
rect 1857 14909 1869 14943
rect 1903 14940 1915 14943
rect 2225 14943 2283 14949
rect 2225 14940 2237 14943
rect 1903 14912 2237 14940
rect 1903 14909 1915 14912
rect 1857 14903 1915 14909
rect 2225 14909 2237 14912
rect 2271 14909 2283 14943
rect 2225 14903 2283 14909
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14940 2559 14943
rect 2866 14940 2872 14952
rect 2547 14912 2872 14940
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 3988 14949 4016 14980
rect 5644 14952 5672 14980
rect 6454 14968 6460 15020
rect 6512 15008 6518 15020
rect 7466 15008 7472 15020
rect 6512 14980 7472 15008
rect 6512 14968 6518 14980
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14940 3479 14943
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 3467 14912 3525 14940
rect 3467 14909 3479 14912
rect 3421 14903 3479 14909
rect 3513 14909 3525 14912
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14909 4031 14943
rect 3973 14903 4031 14909
rect 3528 14872 3556 14903
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 5353 14943 5411 14949
rect 5353 14940 5365 14943
rect 5224 14912 5365 14940
rect 5224 14900 5230 14912
rect 5353 14909 5365 14912
rect 5399 14909 5411 14943
rect 5626 14940 5632 14952
rect 5587 14912 5632 14940
rect 5353 14903 5411 14909
rect 5368 14872 5396 14903
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 7745 14943 7803 14949
rect 7745 14909 7757 14943
rect 7791 14909 7803 14943
rect 7926 14940 7932 14952
rect 7887 14912 7932 14940
rect 7745 14903 7803 14909
rect 6178 14872 6184 14884
rect 3528 14844 5304 14872
rect 5368 14844 6184 14872
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 3602 14804 3608 14816
rect 3563 14776 3608 14804
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4246 14764 4252 14816
rect 4304 14804 4310 14816
rect 4525 14807 4583 14813
rect 4525 14804 4537 14807
rect 4304 14776 4537 14804
rect 4304 14764 4310 14776
rect 4525 14773 4537 14776
rect 4571 14773 4583 14807
rect 4890 14804 4896 14816
rect 4851 14776 4896 14804
rect 4525 14767 4583 14773
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 5169 14807 5227 14813
rect 5169 14804 5181 14807
rect 5040 14776 5181 14804
rect 5040 14764 5046 14776
rect 5169 14773 5181 14776
rect 5215 14773 5227 14807
rect 5276 14804 5304 14844
rect 6178 14832 6184 14844
rect 6236 14832 6242 14884
rect 7377 14875 7435 14881
rect 7377 14841 7389 14875
rect 7423 14872 7435 14875
rect 7760 14872 7788 14903
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8864 14940 8892 15039
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 10134 15036 10140 15088
rect 10192 15076 10198 15088
rect 17773 15079 17831 15085
rect 17773 15076 17785 15079
rect 10192 15048 17785 15076
rect 10192 15036 10198 15048
rect 17773 15045 17785 15048
rect 17819 15045 17831 15079
rect 17773 15039 17831 15045
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 10367 14980 10640 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8864 14912 9045 14940
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 9033 14903 9091 14909
rect 9140 14912 9505 14940
rect 8110 14872 8116 14884
rect 7423 14844 8116 14872
rect 7423 14841 7435 14844
rect 7377 14835 7435 14841
rect 8110 14832 8116 14844
rect 8168 14872 8174 14884
rect 8573 14875 8631 14881
rect 8573 14872 8585 14875
rect 8168 14844 8585 14872
rect 8168 14832 8174 14844
rect 8573 14841 8585 14844
rect 8619 14872 8631 14875
rect 9140 14872 9168 14912
rect 9493 14909 9505 14912
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 8619 14844 9168 14872
rect 9508 14872 9536 14903
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10612 14949 10640 14980
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 16025 15011 16083 15017
rect 16025 15008 16037 15011
rect 14792 14980 16037 15008
rect 14792 14968 14798 14980
rect 16025 14977 16037 14980
rect 16071 14977 16083 15011
rect 16025 14971 16083 14977
rect 10597 14943 10655 14949
rect 10100 14912 10548 14940
rect 10100 14900 10106 14912
rect 10321 14875 10379 14881
rect 10321 14872 10333 14875
rect 9508 14844 10333 14872
rect 8619 14841 8631 14844
rect 8573 14835 8631 14841
rect 6454 14804 6460 14816
rect 5276 14776 6460 14804
rect 5169 14767 5227 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 7524 14776 7573 14804
rect 7524 14764 7530 14776
rect 7561 14773 7573 14776
rect 7607 14773 7619 14807
rect 7561 14767 7619 14773
rect 9030 14764 9036 14816
rect 9088 14804 9094 14816
rect 9140 14804 9168 14844
rect 10321 14841 10333 14844
rect 10367 14872 10379 14875
rect 10413 14875 10471 14881
rect 10413 14872 10425 14875
rect 10367 14844 10425 14872
rect 10367 14841 10379 14844
rect 10321 14835 10379 14841
rect 10413 14841 10425 14844
rect 10459 14841 10471 14875
rect 10413 14835 10471 14841
rect 9088 14776 9168 14804
rect 9309 14807 9367 14813
rect 9088 14764 9094 14776
rect 9309 14773 9321 14807
rect 9355 14804 9367 14807
rect 9398 14804 9404 14816
rect 9355 14776 9404 14804
rect 9355 14773 9367 14776
rect 9309 14767 9367 14773
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10137 14807 10195 14813
rect 10137 14804 10149 14807
rect 9732 14776 10149 14804
rect 9732 14764 9738 14776
rect 10137 14773 10149 14776
rect 10183 14804 10195 14807
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10183 14776 10241 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 10229 14773 10241 14776
rect 10275 14773 10287 14807
rect 10520 14804 10548 14912
rect 10597 14909 10609 14943
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 11057 14943 11115 14949
rect 11057 14940 11069 14943
rect 11020 14912 11069 14940
rect 11020 14900 11026 14912
rect 11057 14909 11069 14912
rect 11103 14909 11115 14943
rect 11057 14903 11115 14909
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14940 11943 14943
rect 12253 14943 12311 14949
rect 12253 14940 12265 14943
rect 11931 14912 12265 14940
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12253 14909 12265 14912
rect 12299 14940 12311 14943
rect 12434 14940 12440 14952
rect 12299 14912 12440 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12434 14900 12440 14912
rect 12492 14940 12498 14952
rect 12802 14940 12808 14952
rect 12492 14912 12808 14940
rect 12492 14900 12498 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13924 14912 14105 14940
rect 13170 14872 13176 14884
rect 13131 14844 13176 14872
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 13924 14816 13952 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 15562 14940 15568 14952
rect 15523 14912 15568 14940
rect 14093 14903 14151 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14940 15715 14943
rect 15746 14940 15752 14952
rect 15703 14912 15752 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 15746 14900 15752 14912
rect 15804 14900 15810 14952
rect 15841 14943 15899 14949
rect 15841 14909 15853 14943
rect 15887 14940 15899 14943
rect 17788 14940 17816 15039
rect 18966 15036 18972 15088
rect 19024 15076 19030 15088
rect 19797 15079 19855 15085
rect 19797 15076 19809 15079
rect 19024 15048 19809 15076
rect 19024 15036 19030 15048
rect 19797 15045 19809 15048
rect 19843 15045 19855 15079
rect 19797 15039 19855 15045
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 15887 14912 16988 14940
rect 17788 14912 18061 14940
rect 15887 14909 15899 14912
rect 15841 14903 15899 14909
rect 14737 14875 14795 14881
rect 14737 14841 14749 14875
rect 14783 14872 14795 14875
rect 14826 14872 14832 14884
rect 14783 14844 14832 14872
rect 14783 14841 14795 14844
rect 14737 14835 14795 14841
rect 14826 14832 14832 14844
rect 14884 14832 14890 14884
rect 15105 14875 15163 14881
rect 15105 14841 15117 14875
rect 15151 14872 15163 14875
rect 15856 14872 15884 14903
rect 15151 14844 15884 14872
rect 15151 14841 15163 14844
rect 15105 14835 15163 14841
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 10520 14776 10701 14804
rect 10229 14767 10287 14773
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 13449 14807 13507 14813
rect 13449 14804 13461 14807
rect 13136 14776 13461 14804
rect 13136 14764 13142 14776
rect 13449 14773 13461 14776
rect 13495 14773 13507 14807
rect 13906 14804 13912 14816
rect 13867 14776 13912 14804
rect 13449 14767 13507 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 15473 14807 15531 14813
rect 15473 14773 15485 14807
rect 15519 14804 15531 14807
rect 15746 14804 15752 14816
rect 15519 14776 15752 14804
rect 15519 14773 15531 14776
rect 15473 14767 15531 14773
rect 15746 14764 15752 14776
rect 15804 14804 15810 14816
rect 16666 14804 16672 14816
rect 15804 14776 16672 14804
rect 15804 14764 15810 14776
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 16960 14813 16988 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18049 14903 18107 14909
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18288 14912 18521 14940
rect 18288 14900 18294 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 19613 14943 19671 14949
rect 19613 14909 19625 14943
rect 19659 14909 19671 14943
rect 19613 14903 19671 14909
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 19628 14872 19656 14903
rect 20346 14900 20352 14952
rect 20404 14940 20410 14952
rect 20844 14943 20902 14949
rect 20844 14940 20856 14943
rect 20404 14912 20856 14940
rect 20404 14900 20410 14912
rect 20844 14909 20856 14912
rect 20890 14909 20902 14943
rect 20844 14903 20902 14909
rect 20947 14943 21005 14949
rect 20947 14909 20959 14943
rect 20993 14940 21005 14943
rect 21542 14940 21548 14952
rect 20993 14912 21548 14940
rect 20993 14909 21005 14912
rect 20947 14903 21005 14909
rect 20073 14875 20131 14881
rect 20073 14872 20085 14875
rect 18380 14844 20085 14872
rect 18380 14832 18386 14844
rect 20073 14841 20085 14844
rect 20119 14841 20131 14875
rect 20859 14872 20887 14903
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 21887 14949 21915 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22281 15107 22339 15113
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 24765 15147 24823 15153
rect 24765 15144 24777 15147
rect 24268 15116 24777 15144
rect 24268 15104 24274 15116
rect 24765 15113 24777 15116
rect 24811 15113 24823 15147
rect 24765 15107 24823 15113
rect 21872 14943 21930 14949
rect 21872 14909 21884 14943
rect 21918 14940 21930 14943
rect 24581 14943 24639 14949
rect 24581 14940 24593 14943
rect 21918 14912 24593 14940
rect 21918 14909 21930 14912
rect 21872 14903 21930 14909
rect 24581 14909 24593 14912
rect 24627 14940 24639 14943
rect 25133 14943 25191 14949
rect 25133 14940 25145 14943
rect 24627 14912 25145 14940
rect 24627 14909 24639 14912
rect 24581 14903 24639 14909
rect 25133 14909 25145 14912
rect 25179 14909 25191 14943
rect 25133 14903 25191 14909
rect 21269 14875 21327 14881
rect 21269 14872 21281 14875
rect 20859 14844 21281 14872
rect 20073 14835 20131 14841
rect 21269 14841 21281 14844
rect 21315 14841 21327 14875
rect 21269 14835 21327 14841
rect 21450 14832 21456 14884
rect 21508 14872 21514 14884
rect 21959 14875 22017 14881
rect 21959 14872 21971 14875
rect 21508 14844 21971 14872
rect 21508 14832 21514 14844
rect 21959 14841 21971 14844
rect 22005 14841 22017 14875
rect 21959 14835 22017 14841
rect 16945 14807 17003 14813
rect 16945 14773 16957 14807
rect 16991 14804 17003 14807
rect 17218 14804 17224 14816
rect 16991 14776 17224 14804
rect 16991 14773 17003 14776
rect 16945 14767 17003 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 17862 14764 17868 14816
rect 17920 14804 17926 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 17920 14776 18153 14804
rect 17920 14764 17926 14776
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18141 14767 18199 14773
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18472 14776 19073 14804
rect 18472 14764 18478 14776
rect 19061 14773 19073 14776
rect 19107 14773 19119 14807
rect 19061 14767 19119 14773
rect 21729 14807 21787 14813
rect 21729 14773 21741 14807
rect 21775 14804 21787 14807
rect 22094 14804 22100 14816
rect 21775 14776 22100 14804
rect 21775 14773 21787 14776
rect 21729 14767 21787 14773
rect 22094 14764 22100 14776
rect 22152 14764 22158 14816
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 23845 14807 23903 14813
rect 23845 14804 23857 14807
rect 23348 14776 23857 14804
rect 23348 14764 23354 14776
rect 23845 14773 23857 14776
rect 23891 14773 23903 14807
rect 23845 14767 23903 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1210 14560 1216 14612
rect 1268 14600 1274 14612
rect 1857 14603 1915 14609
rect 1857 14600 1869 14603
rect 1268 14572 1869 14600
rect 1268 14560 1274 14572
rect 1857 14569 1869 14572
rect 1903 14600 1915 14603
rect 1946 14600 1952 14612
rect 1903 14572 1952 14600
rect 1903 14569 1915 14572
rect 1857 14563 1915 14569
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2332 14572 2820 14600
rect 2332 14541 2360 14572
rect 937 14535 995 14541
rect 937 14501 949 14535
rect 983 14532 995 14535
rect 2317 14535 2375 14541
rect 2317 14532 2329 14535
rect 983 14504 2329 14532
rect 983 14501 995 14504
rect 937 14495 995 14501
rect 2317 14501 2329 14504
rect 2363 14501 2375 14535
rect 2317 14495 2375 14501
rect 2409 14535 2467 14541
rect 2409 14501 2421 14535
rect 2455 14532 2467 14535
rect 2590 14532 2596 14544
rect 2455 14504 2596 14532
rect 2455 14501 2467 14504
rect 2409 14495 2467 14501
rect 2590 14492 2596 14504
rect 2648 14492 2654 14544
rect 2792 14532 2820 14572
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 2924 14572 3525 14600
rect 2924 14560 2930 14572
rect 3513 14569 3525 14572
rect 3559 14569 3571 14603
rect 5166 14600 5172 14612
rect 5127 14572 5172 14600
rect 3513 14563 3571 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5442 14600 5448 14612
rect 5403 14572 5448 14600
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 6457 14603 6515 14609
rect 6457 14569 6469 14603
rect 6503 14600 6515 14603
rect 6638 14600 6644 14612
rect 6503 14572 6644 14600
rect 6503 14569 6515 14572
rect 6457 14563 6515 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7745 14603 7803 14609
rect 7745 14569 7757 14603
rect 7791 14600 7803 14603
rect 7926 14600 7932 14612
rect 7791 14572 7932 14600
rect 7791 14569 7803 14572
rect 7745 14563 7803 14569
rect 7926 14560 7932 14572
rect 7984 14600 7990 14612
rect 8386 14600 8392 14612
rect 7984 14572 8392 14600
rect 7984 14560 7990 14572
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 10962 14600 10968 14612
rect 10827 14572 10968 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 12308 14572 12633 14600
rect 12308 14560 12314 14572
rect 12621 14569 12633 14572
rect 12667 14569 12679 14603
rect 16393 14603 16451 14609
rect 12621 14563 12679 14569
rect 13786 14572 16344 14600
rect 9030 14532 9036 14544
rect 2792 14504 3556 14532
rect 3528 14476 3556 14504
rect 8128 14504 9036 14532
rect 8128 14476 8156 14504
rect 9030 14492 9036 14504
rect 9088 14492 9094 14544
rect 9858 14532 9864 14544
rect 9819 14504 9864 14532
rect 9858 14492 9864 14504
rect 9916 14492 9922 14544
rect 11422 14532 11428 14544
rect 11383 14504 11428 14532
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 12342 14532 12348 14544
rect 12303 14504 12348 14532
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 13786 14532 13814 14572
rect 12820 14504 13814 14532
rect 3510 14424 3516 14476
rect 3568 14424 3574 14476
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4154 14464 4160 14476
rect 4111 14436 4160 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 5534 14464 5540 14476
rect 5495 14436 5540 14464
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 5905 14467 5963 14473
rect 5905 14464 5917 14467
rect 5684 14436 5917 14464
rect 5684 14424 5690 14436
rect 5905 14433 5917 14436
rect 5951 14464 5963 14467
rect 8110 14464 8116 14476
rect 5951 14436 6960 14464
rect 8023 14436 8116 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 5166 14356 5172 14408
rect 5224 14396 5230 14408
rect 5644 14396 5672 14424
rect 5224 14368 5672 14396
rect 5224 14356 5230 14368
rect 2866 14288 2872 14340
rect 2924 14328 2930 14340
rect 3050 14328 3056 14340
rect 2924 14300 3056 14328
rect 2924 14288 2930 14300
rect 3050 14288 3056 14300
rect 3108 14288 3114 14340
rect 4295 14263 4353 14269
rect 4295 14229 4307 14263
rect 4341 14260 4353 14263
rect 4522 14260 4528 14272
rect 4341 14232 4528 14260
rect 4341 14229 4353 14232
rect 4295 14223 4353 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 4614 14220 4620 14272
rect 4672 14260 4678 14272
rect 6932 14269 6960 14436
rect 8110 14424 8116 14436
rect 8168 14424 8174 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 12360 14464 12388 14492
rect 12820 14473 12848 14504
rect 14826 14492 14832 14544
rect 14884 14532 14890 14544
rect 16114 14532 16120 14544
rect 14884 14504 16120 14532
rect 14884 14492 14890 14504
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12360 14436 12817 14464
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14464 13139 14467
rect 13170 14464 13176 14476
rect 13127 14436 13176 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 13170 14424 13176 14436
rect 13228 14464 13234 14476
rect 13354 14464 13360 14476
rect 13228 14436 13360 14464
rect 13228 14424 13234 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 15304 14473 15332 14504
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16316 14532 16344 14572
rect 16393 14569 16405 14603
rect 16439 14600 16451 14603
rect 16482 14600 16488 14612
rect 16439 14572 16488 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 16482 14560 16488 14572
rect 16540 14600 16546 14612
rect 18046 14600 18052 14612
rect 16540 14572 18052 14600
rect 16540 14560 16546 14572
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 23707 14603 23765 14609
rect 23707 14569 23719 14603
rect 23753 14600 23765 14603
rect 24026 14600 24032 14612
rect 23753 14572 24032 14600
rect 23753 14569 23765 14572
rect 23707 14563 23765 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 18322 14532 18328 14544
rect 16316 14504 18328 14532
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 15378 14424 15384 14476
rect 15436 14424 15442 14476
rect 15470 14424 15476 14476
rect 15528 14464 15534 14476
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15528 14436 15577 14464
rect 15528 14424 15534 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 17380 14467 17438 14473
rect 17380 14433 17392 14467
rect 17426 14464 17438 14467
rect 17494 14464 17500 14476
rect 17426 14436 17500 14464
rect 17426 14433 17438 14436
rect 17380 14427 17438 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 18874 14464 18880 14476
rect 18835 14436 18880 14464
rect 18874 14424 18880 14436
rect 18932 14424 18938 14476
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 20936 14467 20994 14473
rect 20936 14464 20948 14467
rect 20680 14436 20948 14464
rect 20680 14424 20686 14436
rect 20936 14433 20948 14436
rect 20982 14433 20994 14467
rect 20936 14427 20994 14433
rect 21980 14467 22038 14473
rect 21980 14433 21992 14467
rect 22026 14464 22038 14467
rect 22278 14464 22284 14476
rect 22026 14436 22284 14464
rect 22026 14433 22038 14436
rect 21980 14427 22038 14433
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 23636 14467 23694 14473
rect 23636 14433 23648 14467
rect 23682 14464 23694 14467
rect 23750 14464 23756 14476
rect 23682 14436 23756 14464
rect 23682 14433 23694 14436
rect 23636 14427 23694 14433
rect 23750 14424 23756 14436
rect 23808 14424 23814 14476
rect 24581 14467 24639 14473
rect 24581 14433 24593 14467
rect 24627 14464 24639 14467
rect 24670 14464 24676 14476
rect 24627 14436 24676 14464
rect 24627 14433 24639 14436
rect 24581 14427 24639 14433
rect 24670 14424 24676 14436
rect 24728 14424 24734 14476
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8938 14396 8944 14408
rect 8619 14368 8944 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8938 14356 8944 14368
rect 8996 14356 9002 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14396 10471 14399
rect 10962 14396 10968 14408
rect 10459 14368 10968 14396
rect 10459 14365 10471 14368
rect 10413 14359 10471 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 11330 14396 11336 14408
rect 11291 14368 11336 14396
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 11974 14396 11980 14408
rect 11935 14368 11980 14396
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 12250 14356 12256 14408
rect 12308 14396 12314 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 12308 14368 13277 14396
rect 12308 14356 12314 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 15396 14396 15424 14424
rect 13265 14359 13323 14365
rect 15304 14368 15424 14396
rect 16025 14399 16083 14405
rect 12710 14288 12716 14340
rect 12768 14328 12774 14340
rect 12897 14331 12955 14337
rect 12897 14328 12909 14331
rect 12768 14300 12909 14328
rect 12768 14288 12774 14300
rect 12897 14297 12909 14300
rect 12943 14297 12955 14331
rect 12897 14291 12955 14297
rect 4709 14263 4767 14269
rect 4709 14260 4721 14263
rect 4672 14232 4721 14260
rect 4672 14220 4678 14232
rect 4709 14229 4721 14232
rect 4755 14229 4767 14263
rect 4709 14223 4767 14229
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7282 14260 7288 14272
rect 6963 14232 7288 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11698 14260 11704 14272
rect 11195 14232 11704 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12526 14220 12532 14272
rect 12584 14260 12590 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 12584 14232 13829 14260
rect 12584 14220 12590 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 14366 14220 14372 14272
rect 14424 14260 14430 14272
rect 14645 14263 14703 14269
rect 14645 14260 14657 14263
rect 14424 14232 14657 14260
rect 14424 14220 14430 14232
rect 14645 14229 14657 14232
rect 14691 14229 14703 14263
rect 14645 14223 14703 14229
rect 15105 14263 15163 14269
rect 15105 14229 15117 14263
rect 15151 14260 15163 14263
rect 15304 14260 15332 14368
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16390 14396 16396 14408
rect 16071 14368 16396 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16390 14356 16396 14368
rect 16448 14356 16454 14408
rect 15381 14331 15439 14337
rect 15381 14297 15393 14331
rect 15427 14328 15439 14331
rect 15930 14328 15936 14340
rect 15427 14300 15936 14328
rect 15427 14297 15439 14300
rect 15381 14291 15439 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 20530 14288 20536 14340
rect 20588 14328 20594 14340
rect 22051 14331 22109 14337
rect 22051 14328 22063 14331
rect 20588 14300 22063 14328
rect 20588 14288 20594 14300
rect 22051 14297 22063 14300
rect 22097 14297 22109 14331
rect 22051 14291 22109 14297
rect 16206 14260 16212 14272
rect 15151 14232 16212 14260
rect 15151 14229 15163 14232
rect 15105 14223 15163 14229
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 16761 14263 16819 14269
rect 16761 14229 16773 14263
rect 16807 14260 16819 14263
rect 17310 14260 17316 14272
rect 16807 14232 17316 14260
rect 16807 14229 16819 14232
rect 16761 14223 16819 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17451 14263 17509 14269
rect 17451 14229 17463 14263
rect 17497 14260 17509 14263
rect 17954 14260 17960 14272
rect 17497 14232 17960 14260
rect 17497 14229 17509 14232
rect 17451 14223 17509 14229
rect 17954 14220 17960 14232
rect 18012 14220 18018 14272
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18230 14260 18236 14272
rect 18187 14232 18236 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18230 14220 18236 14232
rect 18288 14220 18294 14272
rect 18598 14260 18604 14272
rect 18559 14232 18604 14260
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19426 14260 19432 14272
rect 19387 14232 19432 14260
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 20898 14220 20904 14272
rect 20956 14260 20962 14272
rect 21039 14263 21097 14269
rect 21039 14260 21051 14263
rect 20956 14232 21051 14260
rect 20956 14220 20962 14232
rect 21039 14229 21051 14232
rect 21085 14229 21097 14263
rect 21039 14223 21097 14229
rect 24719 14263 24777 14269
rect 24719 14229 24731 14263
rect 24765 14260 24777 14263
rect 24854 14260 24860 14272
rect 24765 14232 24860 14260
rect 24765 14229 24777 14232
rect 24719 14223 24777 14229
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1670 14056 1676 14068
rect 1627 14028 1676 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2041 14059 2099 14065
rect 2041 14025 2053 14059
rect 2087 14056 2099 14059
rect 2130 14056 2136 14068
rect 2087 14028 2136 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2056 13852 2084 14019
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 4893 14059 4951 14065
rect 4893 14025 4905 14059
rect 4939 14056 4951 14059
rect 5166 14056 5172 14068
rect 4939 14028 5172 14056
rect 4939 14025 4951 14028
rect 4893 14019 4951 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 7929 14059 7987 14065
rect 7929 14025 7941 14059
rect 7975 14056 7987 14059
rect 8110 14056 8116 14068
rect 7975 14028 8116 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9674 14016 9680 14068
rect 9732 14016 9738 14068
rect 11333 14059 11391 14065
rect 11333 14025 11345 14059
rect 11379 14056 11391 14059
rect 11422 14056 11428 14068
rect 11379 14028 11428 14056
rect 11379 14025 11391 14028
rect 11333 14019 11391 14025
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 12253 14059 12311 14065
rect 12253 14025 12265 14059
rect 12299 14056 12311 14059
rect 12342 14056 12348 14068
rect 12299 14028 12348 14056
rect 12299 14025 12311 14028
rect 12253 14019 12311 14025
rect 12342 14016 12348 14028
rect 12400 14016 12406 14068
rect 12802 14016 12808 14068
rect 12860 14056 12866 14068
rect 13170 14056 13176 14068
rect 12860 14028 13176 14056
rect 12860 14016 12866 14028
rect 13170 14016 13176 14028
rect 13228 14016 13234 14068
rect 18874 14056 18880 14068
rect 18835 14028 18880 14056
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 24489 14059 24547 14065
rect 24489 14025 24501 14059
rect 24535 14056 24547 14059
rect 24670 14056 24676 14068
rect 24535 14028 24676 14056
rect 24535 14025 24547 14028
rect 24489 14019 24547 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 5626 13988 5632 14000
rect 5368 13960 5632 13988
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2958 13920 2964 13932
rect 2188 13892 2964 13920
rect 2188 13880 2194 13892
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3513 13923 3571 13929
rect 3513 13889 3525 13923
rect 3559 13920 3571 13923
rect 4338 13920 4344 13932
rect 3559 13892 4344 13920
rect 3559 13889 3571 13892
rect 3513 13883 3571 13889
rect 4338 13880 4344 13892
rect 4396 13920 4402 13932
rect 5368 13929 5396 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 6178 13948 6184 14000
rect 6236 13988 6242 14000
rect 9692 13988 9720 14016
rect 6236 13960 9720 13988
rect 6236 13948 6242 13960
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 15896 13960 16221 13988
rect 15896 13948 15902 13960
rect 16209 13957 16221 13960
rect 16255 13988 16267 13991
rect 16850 13988 16856 14000
rect 16255 13960 16856 13988
rect 16255 13957 16267 13960
rect 16209 13951 16267 13957
rect 16850 13948 16856 13960
rect 16908 13948 16914 14000
rect 16942 13948 16948 14000
rect 17000 13988 17006 14000
rect 18233 13991 18291 13997
rect 18233 13988 18245 13991
rect 17000 13960 18245 13988
rect 17000 13948 17006 13960
rect 18233 13957 18245 13960
rect 18279 13957 18291 13991
rect 18233 13951 18291 13957
rect 20346 13948 20352 14000
rect 20404 13988 20410 14000
rect 20404 13960 23474 13988
rect 20404 13948 20410 13960
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 4396 13892 5365 13920
rect 4396 13880 4402 13892
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 5592 13892 6101 13920
rect 5592 13880 5598 13892
rect 6089 13889 6101 13892
rect 6135 13920 6147 13923
rect 7650 13920 7656 13932
rect 6135 13892 7656 13920
rect 6135 13889 6147 13892
rect 6089 13883 6147 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9950 13920 9956 13932
rect 9723 13892 9956 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9950 13880 9956 13892
rect 10008 13920 10014 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10008 13892 10885 13920
rect 10008 13880 10014 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 11388 13892 11621 13920
rect 11388 13880 11394 13892
rect 11609 13889 11621 13892
rect 11655 13889 11667 13923
rect 11609 13883 11667 13889
rect 11974 13880 11980 13932
rect 12032 13920 12038 13932
rect 12526 13920 12532 13932
rect 12032 13892 12532 13920
rect 12032 13880 12038 13892
rect 12526 13880 12532 13892
rect 12584 13880 12590 13932
rect 12802 13920 12808 13932
rect 12763 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 17310 13920 17316 13932
rect 16132 13892 17316 13920
rect 1443 13824 2084 13852
rect 2409 13855 2467 13861
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2409 13821 2421 13855
rect 2455 13852 2467 13855
rect 2590 13852 2596 13864
rect 2455 13824 2596 13852
rect 2455 13821 2467 13824
rect 2409 13815 2467 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13852 6607 13855
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6595 13824 6837 13852
rect 6595 13821 6607 13824
rect 6549 13815 6607 13821
rect 6825 13821 6837 13824
rect 6871 13852 6883 13855
rect 7282 13852 7288 13864
rect 6871 13824 6905 13852
rect 7243 13824 7288 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 2682 13744 2688 13796
rect 2740 13784 2746 13796
rect 2869 13787 2927 13793
rect 2869 13784 2881 13787
rect 2740 13756 2881 13784
rect 2740 13744 2746 13756
rect 2869 13753 2881 13756
rect 2915 13753 2927 13787
rect 2869 13747 2927 13753
rect 2961 13787 3019 13793
rect 2961 13753 2973 13787
rect 3007 13784 3019 13787
rect 3142 13784 3148 13796
rect 3007 13756 3148 13784
rect 3007 13753 3019 13756
rect 2961 13747 3019 13753
rect 3142 13744 3148 13756
rect 3200 13784 3206 13796
rect 3789 13787 3847 13793
rect 3789 13784 3801 13787
rect 3200 13756 3801 13784
rect 3200 13744 3206 13756
rect 3789 13753 3801 13756
rect 3835 13753 3847 13787
rect 3789 13747 3847 13753
rect 3970 13744 3976 13796
rect 4028 13784 4034 13796
rect 4614 13784 4620 13796
rect 4028 13756 4620 13784
rect 4028 13744 4034 13756
rect 4614 13744 4620 13756
rect 4672 13784 4678 13796
rect 5077 13787 5135 13793
rect 5077 13784 5089 13787
rect 4672 13756 5089 13784
rect 4672 13744 4678 13756
rect 5077 13753 5089 13756
rect 5123 13753 5135 13787
rect 5077 13747 5135 13753
rect 5166 13744 5172 13796
rect 5224 13784 5230 13796
rect 5224 13756 5269 13784
rect 5224 13744 5230 13756
rect 6638 13744 6644 13796
rect 6696 13784 6702 13796
rect 6840 13784 6868 13815
rect 7282 13812 7288 13824
rect 7340 13812 7346 13864
rect 7926 13852 7932 13864
rect 7852 13824 7932 13852
rect 7852 13784 7880 13824
rect 7926 13812 7932 13824
rect 7984 13812 7990 13864
rect 8754 13861 8760 13864
rect 8716 13855 8760 13861
rect 8716 13852 8728 13855
rect 8667 13824 8728 13852
rect 8716 13821 8728 13824
rect 8716 13815 8760 13821
rect 8747 13812 8760 13815
rect 8812 13812 8818 13864
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 8904 13824 9505 13852
rect 8904 13812 8910 13824
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13412 13824 13829 13852
rect 13412 13812 13418 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 13817 13815 13875 13821
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14458 13852 14464 13864
rect 14415 13824 14464 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15746 13852 15752 13864
rect 15335 13824 15752 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 16132 13861 16160 13892
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 23446 13920 23474 13960
rect 23934 13948 23940 14000
rect 23992 13988 23998 14000
rect 24765 13991 24823 13997
rect 24765 13988 24777 13991
rect 23992 13960 24777 13988
rect 23992 13948 23998 13960
rect 24765 13957 24777 13960
rect 24811 13957 24823 13991
rect 24765 13951 24823 13957
rect 25133 13923 25191 13929
rect 25133 13920 25145 13923
rect 23446 13892 25145 13920
rect 16117 13855 16175 13861
rect 16117 13821 16129 13855
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 16393 13855 16451 13861
rect 16393 13821 16405 13855
rect 16439 13852 16451 13855
rect 16482 13852 16488 13864
rect 16439 13824 16488 13852
rect 16439 13821 16451 13824
rect 16393 13815 16451 13821
rect 16482 13812 16488 13824
rect 16540 13852 16546 13864
rect 16758 13852 16764 13864
rect 16540 13824 16764 13852
rect 16540 13812 16546 13824
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17828 13824 18061 13852
rect 17828 13812 17834 13824
rect 18049 13821 18061 13824
rect 18095 13852 18107 13855
rect 18509 13855 18567 13861
rect 18509 13852 18521 13855
rect 18095 13824 18521 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18509 13821 18521 13824
rect 18555 13821 18567 13855
rect 19426 13852 19432 13864
rect 19387 13824 19432 13852
rect 18509 13815 18567 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20438 13812 20444 13864
rect 20496 13852 20502 13864
rect 24596 13861 24624 13892
rect 25133 13889 25145 13892
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 20752 13855 20810 13861
rect 20752 13852 20764 13855
rect 20496 13824 20764 13852
rect 20496 13812 20502 13824
rect 20752 13821 20764 13824
rect 20798 13852 20810 13855
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 20798 13824 21189 13852
rect 20798 13821 20810 13824
rect 20752 13815 20810 13821
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 21177 13815 21235 13821
rect 22624 13855 22682 13861
rect 22624 13821 22636 13855
rect 22670 13852 22682 13855
rect 24581 13855 24639 13861
rect 22670 13824 22876 13852
rect 22670 13821 22682 13824
rect 22624 13815 22682 13821
rect 6696 13756 7880 13784
rect 8747 13784 8775 13812
rect 10039 13787 10097 13793
rect 8747 13756 9260 13784
rect 6696 13744 6702 13756
rect 198 13676 204 13728
rect 256 13716 262 13728
rect 3234 13716 3240 13728
rect 256 13688 3240 13716
rect 256 13676 262 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4154 13676 4160 13728
rect 4212 13716 4218 13728
rect 6914 13716 6920 13728
rect 4212 13688 4257 13716
rect 6875 13688 6920 13716
rect 4212 13676 4218 13688
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 7834 13716 7840 13728
rect 7708 13688 7840 13716
rect 7708 13676 7714 13688
rect 7834 13676 7840 13688
rect 7892 13716 7898 13728
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7892 13688 8217 13716
rect 7892 13676 7898 13688
rect 8205 13685 8217 13688
rect 8251 13716 8263 13719
rect 8294 13716 8300 13728
rect 8251 13688 8300 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8803 13719 8861 13725
rect 8803 13685 8815 13719
rect 8849 13716 8861 13719
rect 9030 13716 9036 13728
rect 8849 13688 9036 13716
rect 8849 13685 8861 13688
rect 8803 13679 8861 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 9232 13725 9260 13756
rect 10039 13753 10051 13787
rect 10085 13784 10097 13787
rect 10686 13784 10692 13796
rect 10085 13756 10692 13784
rect 10085 13753 10097 13756
rect 10039 13747 10097 13753
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 12598 13787 12656 13793
rect 12598 13784 12610 13787
rect 12452 13756 12610 13784
rect 12452 13728 12480 13756
rect 12598 13753 12610 13756
rect 12644 13753 12656 13787
rect 14690 13787 14748 13793
rect 14690 13784 14702 13787
rect 12598 13747 12656 13753
rect 14200 13756 14702 13784
rect 9217 13719 9275 13725
rect 9217 13685 9229 13719
rect 9263 13716 9275 13719
rect 9490 13716 9496 13728
rect 9263 13688 9496 13716
rect 9263 13685 9275 13688
rect 9217 13679 9275 13685
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 10597 13719 10655 13725
rect 10597 13685 10609 13719
rect 10643 13716 10655 13719
rect 10778 13716 10784 13728
rect 10643 13688 10784 13716
rect 10643 13685 10655 13688
rect 10597 13679 10655 13685
rect 10778 13676 10784 13688
rect 10836 13676 10842 13728
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 13262 13716 13268 13728
rect 12768 13688 13268 13716
rect 12768 13676 12774 13688
rect 13262 13676 13268 13688
rect 13320 13716 13326 13728
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 13320 13688 13461 13716
rect 13320 13676 13326 13688
rect 13449 13685 13461 13688
rect 13495 13685 13507 13719
rect 13449 13679 13507 13685
rect 13998 13676 14004 13728
rect 14056 13716 14062 13728
rect 14200 13725 14228 13756
rect 14690 13753 14702 13756
rect 14736 13753 14748 13787
rect 14690 13747 14748 13753
rect 15470 13744 15476 13796
rect 15528 13784 15534 13796
rect 15565 13787 15623 13793
rect 15565 13784 15577 13787
rect 15528 13756 15577 13784
rect 15528 13744 15534 13756
rect 15565 13753 15577 13756
rect 15611 13753 15623 13787
rect 15565 13747 15623 13753
rect 20622 13744 20628 13796
rect 20680 13784 20686 13796
rect 21545 13787 21603 13793
rect 21545 13784 21557 13787
rect 20680 13756 21557 13784
rect 20680 13744 20686 13756
rect 21545 13753 21557 13756
rect 21591 13753 21603 13787
rect 21545 13747 21603 13753
rect 14185 13719 14243 13725
rect 14185 13716 14197 13719
rect 14056 13688 14197 13716
rect 14056 13676 14062 13688
rect 14185 13685 14197 13688
rect 14231 13685 14243 13719
rect 15930 13716 15936 13728
rect 15891 13688 15936 13716
rect 14185 13679 14243 13685
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16574 13716 16580 13728
rect 16535 13688 16580 13716
rect 16574 13676 16580 13688
rect 16632 13676 16638 13728
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17034 13716 17040 13728
rect 16908 13688 17040 13716
rect 16908 13676 16914 13688
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 17402 13716 17408 13728
rect 17363 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 19426 13716 19432 13728
rect 19387 13688 19432 13716
rect 19426 13676 19432 13688
rect 19484 13676 19490 13728
rect 19978 13676 19984 13728
rect 20036 13716 20042 13728
rect 20855 13719 20913 13725
rect 20855 13716 20867 13719
rect 20036 13688 20867 13716
rect 20036 13676 20042 13688
rect 20855 13685 20867 13688
rect 20901 13685 20913 13719
rect 20855 13679 20913 13685
rect 22005 13719 22063 13725
rect 22005 13685 22017 13719
rect 22051 13716 22063 13719
rect 22278 13716 22284 13728
rect 22051 13688 22284 13716
rect 22051 13685 22063 13688
rect 22005 13679 22063 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22554 13676 22560 13728
rect 22612 13716 22618 13728
rect 22695 13719 22753 13725
rect 22695 13716 22707 13719
rect 22612 13688 22707 13716
rect 22612 13676 22618 13688
rect 22695 13685 22707 13688
rect 22741 13685 22753 13719
rect 22848 13716 22876 13824
rect 24581 13821 24593 13855
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 23014 13716 23020 13728
rect 22848 13688 23020 13716
rect 22695 13679 22753 13685
rect 23014 13676 23020 13688
rect 23072 13676 23078 13728
rect 23750 13676 23756 13728
rect 23808 13716 23814 13728
rect 23845 13719 23903 13725
rect 23845 13716 23857 13719
rect 23808 13688 23857 13716
rect 23808 13676 23814 13688
rect 23845 13685 23857 13688
rect 23891 13685 23903 13719
rect 23845 13679 23903 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1302 13472 1308 13524
rect 1360 13512 1366 13524
rect 1673 13515 1731 13521
rect 1673 13512 1685 13515
rect 1360 13484 1685 13512
rect 1360 13472 1366 13484
rect 1673 13481 1685 13484
rect 1719 13481 1731 13515
rect 2038 13512 2044 13524
rect 1999 13484 2044 13512
rect 1673 13475 1731 13481
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 2498 13512 2504 13524
rect 2424 13484 2504 13512
rect 2056 13376 2084 13472
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 2056 13348 2237 13376
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 2424 13308 2452 13484
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 3142 13512 3148 13524
rect 3103 13484 3148 13512
rect 3142 13472 3148 13484
rect 3200 13472 3206 13524
rect 3510 13512 3516 13524
rect 3471 13484 3516 13512
rect 3510 13472 3516 13484
rect 3568 13472 3574 13524
rect 4893 13515 4951 13521
rect 4893 13481 4905 13515
rect 4939 13512 4951 13515
rect 5166 13512 5172 13524
rect 4939 13484 5172 13512
rect 4939 13481 4951 13484
rect 4893 13475 4951 13481
rect 5166 13472 5172 13484
rect 5224 13512 5230 13524
rect 5905 13515 5963 13521
rect 5905 13512 5917 13515
rect 5224 13484 5917 13512
rect 5224 13472 5230 13484
rect 5905 13481 5917 13484
rect 5951 13481 5963 13515
rect 5905 13475 5963 13481
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 9858 13512 9864 13524
rect 8803 13484 9864 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 11238 13512 11244 13524
rect 10054 13484 11244 13512
rect 2587 13447 2645 13453
rect 2587 13413 2599 13447
rect 2633 13444 2645 13447
rect 3234 13444 3240 13456
rect 2633 13416 3240 13444
rect 2633 13413 2645 13416
rect 2587 13407 2645 13413
rect 3234 13404 3240 13416
rect 3292 13444 3298 13456
rect 5306 13447 5364 13453
rect 5306 13444 5318 13447
rect 3292 13416 5318 13444
rect 3292 13404 3298 13416
rect 5306 13413 5318 13416
rect 5352 13413 5364 13447
rect 5306 13407 5364 13413
rect 8199 13447 8257 13453
rect 8199 13413 8211 13447
rect 8245 13444 8257 13447
rect 8846 13444 8852 13456
rect 8245 13416 8852 13444
rect 8245 13413 8257 13416
rect 8199 13407 8257 13413
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 3878 13376 3884 13388
rect 2556 13348 3884 13376
rect 2556 13336 2562 13348
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4982 13376 4988 13388
rect 4943 13348 4988 13376
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5166 13336 5172 13388
rect 5224 13376 5230 13388
rect 5321 13376 5349 13407
rect 8846 13404 8852 13416
rect 8904 13404 8910 13456
rect 9493 13447 9551 13453
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 9582 13444 9588 13456
rect 9539 13416 9588 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 9766 13404 9772 13456
rect 9824 13444 9830 13456
rect 10054 13444 10082 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 12069 13515 12127 13521
rect 12069 13481 12081 13515
rect 12115 13512 12127 13515
rect 12434 13512 12440 13524
rect 12115 13484 12440 13512
rect 12115 13481 12127 13484
rect 12069 13475 12127 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 13998 13512 14004 13524
rect 13959 13484 14004 13512
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 14642 13512 14648 13524
rect 14424 13484 14648 13512
rect 14424 13472 14430 13484
rect 14642 13472 14648 13484
rect 14700 13472 14706 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 17034 13512 17040 13524
rect 16264 13484 17040 13512
rect 16264 13472 16270 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17494 13512 17500 13524
rect 17368 13484 17500 13512
rect 17368 13472 17374 13484
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18564 13484 19334 13512
rect 18564 13472 18570 13484
rect 9824 13416 10082 13444
rect 9824 13404 9830 13416
rect 10686 13404 10692 13456
rect 10744 13444 10750 13456
rect 11511 13447 11569 13453
rect 11511 13444 11523 13447
rect 10744 13416 11523 13444
rect 10744 13404 10750 13416
rect 11511 13413 11523 13416
rect 11557 13444 11569 13447
rect 12158 13444 12164 13456
rect 11557 13416 12164 13444
rect 11557 13413 11569 13416
rect 11511 13407 11569 13413
rect 12158 13404 12164 13416
rect 12216 13404 12222 13456
rect 14016 13444 14044 13472
rect 15610 13447 15668 13453
rect 15610 13444 15622 13447
rect 14016 13416 15622 13444
rect 15610 13413 15622 13416
rect 15656 13413 15668 13447
rect 15610 13407 15668 13413
rect 16390 13404 16396 13456
rect 16448 13444 16454 13456
rect 18046 13444 18052 13456
rect 16448 13416 18052 13444
rect 16448 13404 16454 13416
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18785 13447 18843 13453
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 18874 13444 18880 13456
rect 18831 13416 18880 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 18874 13404 18880 13416
rect 18932 13404 18938 13456
rect 19306 13444 19334 13484
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 24765 13515 24823 13521
rect 24765 13512 24777 13515
rect 24176 13484 24777 13512
rect 24176 13472 24182 13484
rect 24765 13481 24777 13484
rect 24811 13481 24823 13515
rect 24765 13475 24823 13481
rect 20070 13444 20076 13456
rect 19306 13416 20076 13444
rect 20070 13404 20076 13416
rect 20128 13444 20134 13456
rect 27614 13444 27620 13456
rect 20128 13416 27620 13444
rect 20128 13404 20134 13416
rect 27614 13404 27620 13416
rect 27672 13404 27678 13456
rect 6892 13379 6950 13385
rect 6892 13376 6904 13379
rect 5224 13348 5349 13376
rect 5597 13348 6904 13376
rect 5224 13336 5230 13348
rect 3142 13308 3148 13320
rect 2424 13280 3148 13308
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 3510 13268 3516 13320
rect 3568 13308 3574 13320
rect 4246 13308 4252 13320
rect 3568 13280 4252 13308
rect 3568 13268 3574 13280
rect 4246 13268 4252 13280
rect 4304 13308 4310 13320
rect 5597 13308 5625 13348
rect 6892 13345 6904 13348
rect 6938 13376 6950 13379
rect 7098 13376 7104 13388
rect 6938 13348 7104 13376
rect 6938 13345 6950 13348
rect 6892 13339 6950 13345
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13376 7895 13379
rect 7926 13376 7932 13388
rect 7883 13348 7932 13376
rect 7883 13345 7895 13348
rect 7837 13339 7895 13345
rect 7926 13336 7932 13348
rect 7984 13376 7990 13388
rect 9306 13376 9312 13388
rect 7984 13348 9312 13376
rect 7984 13336 7990 13348
rect 9306 13336 9312 13348
rect 9364 13336 9370 13388
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12124 13348 12909 13376
rect 12124 13336 12130 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 13170 13376 13176 13388
rect 13131 13348 13176 13376
rect 12897 13339 12955 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 14826 13376 14832 13388
rect 14148 13348 14832 13376
rect 14148 13336 14154 13348
rect 14826 13336 14832 13348
rect 14884 13376 14890 13388
rect 15289 13379 15347 13385
rect 15289 13376 15301 13379
rect 14884 13348 15301 13376
rect 14884 13336 14890 13348
rect 15289 13345 15301 13348
rect 15335 13345 15347 13379
rect 15289 13339 15347 13345
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 16724 13348 16988 13376
rect 16724 13336 16730 13348
rect 10134 13308 10140 13320
rect 4304 13280 5625 13308
rect 10095 13280 10140 13308
rect 4304 13268 4310 13280
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 11146 13308 11152 13320
rect 10560 13280 11152 13308
rect 10560 13268 10566 13280
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 11296 13280 13369 13308
rect 11296 13268 11302 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 14458 13308 14464 13320
rect 14371 13280 14464 13308
rect 13357 13271 13415 13277
rect 14458 13268 14464 13280
rect 14516 13308 14522 13320
rect 14516 13280 16896 13308
rect 14516 13268 14522 13280
rect 3694 13200 3700 13252
rect 3752 13240 3758 13252
rect 3878 13240 3884 13252
rect 3752 13212 3884 13240
rect 3752 13200 3758 13212
rect 3878 13200 3884 13212
rect 3936 13200 3942 13252
rect 12989 13243 13047 13249
rect 12989 13209 13001 13243
rect 13035 13240 13047 13243
rect 13262 13240 13268 13252
rect 13035 13212 13268 13240
rect 13035 13209 13047 13212
rect 12989 13203 13047 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14918 13240 14924 13252
rect 14332 13212 14924 13240
rect 14332 13200 14338 13212
rect 14918 13200 14924 13212
rect 14976 13240 14982 13252
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 14976 13212 15025 13240
rect 14976 13200 14982 13212
rect 15013 13209 15025 13212
rect 15059 13209 15071 13243
rect 15013 13203 15071 13209
rect 15838 13200 15844 13252
rect 15896 13240 15902 13252
rect 15896 13212 16528 13240
rect 15896 13200 15902 13212
rect 16500 13184 16528 13212
rect 2682 13132 2688 13184
rect 2740 13172 2746 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 2740 13144 3801 13172
rect 2740 13132 2746 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 6963 13175 7021 13181
rect 6963 13141 6975 13175
rect 7009 13172 7021 13175
rect 8110 13172 8116 13184
rect 7009 13144 8116 13172
rect 7009 13141 7021 13144
rect 6963 13135 7021 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 10778 13172 10784 13184
rect 10735 13144 10784 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11330 13132 11336 13184
rect 11388 13172 11394 13184
rect 13906 13172 13912 13184
rect 11388 13144 13912 13172
rect 11388 13132 11394 13144
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 16206 13172 16212 13184
rect 16167 13144 16212 13172
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 16482 13172 16488 13184
rect 16443 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 16868 13172 16896 13280
rect 16960 13240 16988 13348
rect 17034 13336 17040 13388
rect 17092 13376 17098 13388
rect 17310 13376 17316 13388
rect 17092 13348 17137 13376
rect 17271 13348 17316 13376
rect 17092 13336 17098 13348
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 20772 13348 21005 13376
rect 20772 13336 20778 13348
rect 20993 13345 21005 13348
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 22465 13379 22523 13385
rect 22465 13345 22477 13379
rect 22511 13376 22523 13379
rect 22646 13376 22652 13388
rect 22511 13348 22652 13376
rect 22511 13345 22523 13348
rect 22465 13339 22523 13345
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 23636 13379 23694 13385
rect 23636 13345 23648 13379
rect 23682 13376 23694 13379
rect 23934 13376 23940 13388
rect 23682 13348 23940 13376
rect 23682 13345 23694 13348
rect 23636 13339 23694 13345
rect 23934 13336 23940 13348
rect 23992 13336 23998 13388
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 24268 13348 24593 13376
rect 24268 13336 24274 13348
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 17770 13308 17776 13320
rect 17731 13280 17776 13308
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13308 18751 13311
rect 19978 13308 19984 13320
rect 18739 13280 19984 13308
rect 18739 13277 18751 13280
rect 18693 13271 18751 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22738 13308 22744 13320
rect 22244 13280 22744 13308
rect 22244 13268 22250 13280
rect 22738 13268 22744 13280
rect 22796 13268 22802 13320
rect 17034 13240 17040 13252
rect 16960 13212 17040 13240
rect 17034 13200 17040 13212
rect 17092 13240 17098 13252
rect 17129 13243 17187 13249
rect 17129 13240 17141 13243
rect 17092 13212 17141 13240
rect 17092 13200 17098 13212
rect 17129 13209 17141 13212
rect 17175 13209 17187 13243
rect 19242 13240 19248 13252
rect 19203 13212 19248 13240
rect 17129 13203 17187 13209
rect 19242 13200 19248 13212
rect 19300 13240 19306 13252
rect 20165 13243 20223 13249
rect 20165 13240 20177 13243
rect 19300 13212 20177 13240
rect 19300 13200 19306 13212
rect 20165 13209 20177 13212
rect 20211 13209 20223 13243
rect 21818 13240 21824 13252
rect 20165 13203 20223 13209
rect 21238 13212 21824 13240
rect 21238 13172 21266 13212
rect 21818 13200 21824 13212
rect 21876 13200 21882 13252
rect 21358 13172 21364 13184
rect 16868 13144 21266 13172
rect 21319 13144 21364 13172
rect 21358 13132 21364 13144
rect 21416 13132 21422 13184
rect 22695 13175 22753 13181
rect 22695 13141 22707 13175
rect 22741 13172 22753 13175
rect 22830 13172 22836 13184
rect 22741 13144 22836 13172
rect 22741 13141 22753 13144
rect 22695 13135 22753 13141
rect 22830 13132 22836 13144
rect 22888 13132 22894 13184
rect 23707 13175 23765 13181
rect 23707 13141 23719 13175
rect 23753 13172 23765 13175
rect 23842 13172 23848 13184
rect 23753 13144 23848 13172
rect 23753 13141 23765 13144
rect 23707 13135 23765 13141
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2038 12928 2044 12980
rect 2096 12968 2102 12980
rect 2222 12968 2228 12980
rect 2096 12940 2228 12968
rect 2096 12928 2102 12940
rect 2222 12928 2228 12940
rect 2280 12928 2286 12980
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3234 12968 3240 12980
rect 3191 12940 3240 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 4154 12968 4160 12980
rect 3436 12940 4160 12968
rect 2590 12860 2596 12912
rect 2648 12900 2654 12912
rect 3436 12909 3464 12940
rect 4154 12928 4160 12940
rect 4212 12928 4218 12980
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 4982 12968 4988 12980
rect 4755 12940 4988 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5077 12971 5135 12977
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5166 12968 5172 12980
rect 5123 12940 5172 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5166 12928 5172 12940
rect 5224 12968 5230 12980
rect 5994 12968 6000 12980
rect 5224 12940 6000 12968
rect 5224 12928 5230 12940
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 7098 12968 7104 12980
rect 7059 12940 7104 12968
rect 7098 12928 7104 12940
rect 7156 12928 7162 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7469 12971 7527 12977
rect 7469 12968 7481 12971
rect 7248 12940 7481 12968
rect 7248 12928 7254 12940
rect 7469 12937 7481 12940
rect 7515 12937 7527 12971
rect 7469 12931 7527 12937
rect 8846 12928 8852 12980
rect 8904 12928 8910 12980
rect 10502 12968 10508 12980
rect 10463 12940 10508 12968
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 14884 12940 14933 12968
rect 14884 12928 14890 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 17126 12928 17132 12980
rect 17184 12968 17190 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 17184 12940 17785 12968
rect 17184 12928 17190 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 18509 12971 18567 12977
rect 18509 12937 18521 12971
rect 18555 12968 18567 12971
rect 18598 12968 18604 12980
rect 18555 12940 18604 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 19705 12971 19763 12977
rect 18800 12940 19656 12968
rect 3421 12903 3479 12909
rect 3421 12900 3433 12903
rect 2648 12872 3433 12900
rect 2648 12860 2654 12872
rect 3421 12869 3433 12872
rect 3467 12869 3479 12903
rect 5350 12900 5356 12912
rect 3421 12863 3479 12869
rect 3712 12872 5356 12900
rect 3712 12844 3740 12872
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 8294 12900 8300 12912
rect 8159 12872 8300 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 8294 12860 8300 12872
rect 8352 12900 8358 12912
rect 8864 12900 8892 12928
rect 9493 12903 9551 12909
rect 9493 12900 9505 12903
rect 8352 12872 9505 12900
rect 8352 12860 8358 12872
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 2133 12835 2191 12841
rect 2133 12832 2145 12835
rect 1360 12804 2145 12832
rect 1360 12792 1366 12804
rect 2133 12801 2145 12804
rect 2179 12801 2191 12835
rect 3694 12832 3700 12844
rect 3607 12804 3700 12832
rect 2133 12795 2191 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 3970 12832 3976 12844
rect 3931 12804 3976 12832
rect 3970 12792 3976 12804
rect 4028 12792 4034 12844
rect 5534 12832 5540 12844
rect 5495 12804 5540 12832
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7064 12804 8217 12832
rect 7064 12792 7070 12804
rect 8205 12801 8217 12804
rect 8251 12832 8263 12835
rect 8846 12832 8852 12844
rect 8251 12804 8852 12832
rect 8251 12801 8263 12804
rect 8205 12795 8263 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 7260 12767 7318 12773
rect 7260 12733 7272 12767
rect 7306 12764 7318 12767
rect 7469 12767 7527 12773
rect 7469 12764 7481 12767
rect 7306 12736 7481 12764
rect 7306 12733 7318 12736
rect 7260 12727 7318 12733
rect 7469 12733 7481 12736
rect 7515 12764 7527 12767
rect 7515 12736 7788 12764
rect 7515 12733 7527 12736
rect 7469 12727 7527 12733
rect 1949 12699 2007 12705
rect 1949 12665 1961 12699
rect 1995 12696 2007 12699
rect 2130 12696 2136 12708
rect 1995 12668 2136 12696
rect 1995 12665 2007 12668
rect 1949 12659 2007 12665
rect 2130 12656 2136 12668
rect 2188 12696 2194 12708
rect 2225 12699 2283 12705
rect 2225 12696 2237 12699
rect 2188 12668 2237 12696
rect 2188 12656 2194 12668
rect 2225 12665 2237 12668
rect 2271 12665 2283 12699
rect 2225 12659 2283 12665
rect 2777 12699 2835 12705
rect 2777 12665 2789 12699
rect 2823 12696 2835 12699
rect 3789 12699 3847 12705
rect 2823 12668 3648 12696
rect 2823 12665 2835 12668
rect 2777 12659 2835 12665
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 3234 12628 3240 12640
rect 2924 12600 3240 12628
rect 2924 12588 2930 12600
rect 3234 12588 3240 12600
rect 3292 12588 3298 12640
rect 3620 12628 3648 12668
rect 3789 12665 3801 12699
rect 3835 12696 3847 12699
rect 4154 12696 4160 12708
rect 3835 12668 4160 12696
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 4154 12656 4160 12668
rect 4212 12656 4218 12708
rect 5261 12699 5319 12705
rect 5261 12696 5273 12699
rect 4908 12668 5273 12696
rect 4908 12628 4936 12668
rect 5261 12665 5273 12668
rect 5307 12665 5319 12699
rect 5261 12659 5319 12665
rect 3620 12600 4936 12628
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5276 12628 5304 12659
rect 5350 12656 5356 12708
rect 5408 12696 5414 12708
rect 7098 12696 7104 12708
rect 5408 12668 5453 12696
rect 6196 12668 7104 12696
rect 5408 12656 5414 12668
rect 6196 12637 6224 12668
rect 7098 12656 7104 12668
rect 7156 12656 7162 12708
rect 6181 12631 6239 12637
rect 6181 12628 6193 12631
rect 5224 12600 6193 12628
rect 5224 12588 5230 12600
rect 6181 12597 6193 12600
rect 6227 12597 6239 12631
rect 6181 12591 6239 12597
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 7006 12628 7012 12640
rect 6696 12600 7012 12628
rect 6696 12588 6702 12600
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7331 12631 7389 12637
rect 7331 12597 7343 12631
rect 7377 12628 7389 12631
rect 7558 12628 7564 12640
rect 7377 12600 7564 12628
rect 7377 12597 7389 12600
rect 7331 12591 7389 12597
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 7760 12637 7788 12736
rect 8567 12699 8625 12705
rect 8567 12665 8579 12699
rect 8613 12696 8625 12699
rect 8956 12696 8984 12872
rect 9493 12869 9505 12872
rect 9539 12900 9551 12903
rect 10686 12900 10692 12912
rect 9539 12872 10692 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 10686 12860 10692 12872
rect 10744 12860 10750 12912
rect 11701 12903 11759 12909
rect 11701 12869 11713 12903
rect 11747 12900 11759 12903
rect 12158 12900 12164 12912
rect 11747 12872 12164 12900
rect 11747 12869 11759 12872
rect 11701 12863 11759 12869
rect 12158 12860 12164 12872
rect 12216 12900 12222 12912
rect 13998 12900 14004 12912
rect 12216 12872 14004 12900
rect 12216 12860 12222 12872
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 16209 12903 16267 12909
rect 16209 12869 16221 12903
rect 16255 12900 16267 12903
rect 16390 12900 16396 12912
rect 16255 12872 16396 12900
rect 16255 12869 16267 12872
rect 16209 12863 16267 12869
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 16666 12860 16672 12912
rect 16724 12900 16730 12912
rect 16850 12900 16856 12912
rect 16724 12872 16856 12900
rect 16724 12860 16730 12872
rect 16850 12860 16856 12872
rect 16908 12860 16914 12912
rect 18230 12860 18236 12912
rect 18288 12900 18294 12912
rect 18800 12900 18828 12940
rect 19242 12900 19248 12912
rect 18288 12872 18828 12900
rect 19203 12872 19248 12900
rect 18288 12860 18294 12872
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 19628 12900 19656 12940
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 19978 12968 19984 12980
rect 19751 12940 19984 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 20220 12940 21465 12968
rect 20220 12928 20226 12940
rect 21453 12937 21465 12940
rect 21499 12968 21511 12971
rect 21545 12971 21603 12977
rect 21545 12968 21557 12971
rect 21499 12940 21557 12968
rect 21499 12937 21511 12940
rect 21453 12931 21511 12937
rect 21545 12937 21557 12940
rect 21591 12937 21603 12971
rect 21545 12931 21603 12937
rect 22830 12928 22836 12980
rect 22888 12968 22894 12980
rect 23014 12968 23020 12980
rect 22888 12940 23020 12968
rect 22888 12928 22894 12940
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24397 12971 24455 12977
rect 24397 12968 24409 12971
rect 24268 12940 24409 12968
rect 24268 12928 24274 12940
rect 24397 12937 24409 12940
rect 24443 12937 24455 12971
rect 24397 12931 24455 12937
rect 21177 12903 21235 12909
rect 21177 12900 21189 12903
rect 19628 12872 21189 12900
rect 21177 12869 21189 12872
rect 21223 12869 21235 12903
rect 21177 12863 21235 12869
rect 10962 12832 10968 12844
rect 10923 12804 10968 12832
rect 10962 12792 10968 12804
rect 11020 12832 11026 12844
rect 12667 12835 12725 12841
rect 11020 12804 12607 12832
rect 11020 12792 11026 12804
rect 12579 12773 12607 12804
rect 12667 12801 12679 12835
rect 12713 12832 12725 12835
rect 18506 12832 18512 12844
rect 12713 12804 18512 12832
rect 12713 12801 12725 12804
rect 12667 12795 12725 12801
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 19260 12832 19288 12860
rect 20257 12835 20315 12841
rect 20257 12832 20269 12835
rect 19260 12804 20269 12832
rect 20257 12801 20269 12804
rect 20303 12801 20315 12835
rect 20622 12832 20628 12844
rect 20583 12804 20628 12832
rect 20257 12795 20315 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21192 12832 21220 12863
rect 23658 12860 23664 12912
rect 23716 12900 23722 12912
rect 24765 12903 24823 12909
rect 24765 12900 24777 12903
rect 23716 12872 24777 12900
rect 23716 12860 23722 12872
rect 24765 12869 24777 12872
rect 24811 12869 24823 12903
rect 24765 12863 24823 12869
rect 21192 12804 22232 12832
rect 12564 12767 12622 12773
rect 12564 12733 12576 12767
rect 12610 12764 12622 12767
rect 12802 12764 12808 12776
rect 12610 12736 12808 12764
rect 12610 12733 12622 12736
rect 12564 12727 12622 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13538 12764 13544 12776
rect 13499 12736 13544 12764
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 15470 12764 15476 12776
rect 14884 12736 15476 12764
rect 14884 12724 14890 12736
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 22204 12773 22232 12804
rect 21453 12767 21511 12773
rect 21453 12733 21465 12767
rect 21499 12764 21511 12767
rect 21729 12767 21787 12773
rect 21729 12764 21741 12767
rect 21499 12736 21741 12764
rect 21499 12733 21511 12736
rect 21453 12727 21511 12733
rect 21729 12733 21741 12736
rect 21775 12733 21787 12767
rect 21729 12727 21787 12733
rect 22189 12767 22247 12773
rect 22189 12733 22201 12767
rect 22235 12733 22247 12767
rect 24581 12767 24639 12773
rect 24581 12764 24593 12767
rect 22189 12727 22247 12733
rect 23446 12736 24593 12764
rect 8613 12668 8984 12696
rect 10137 12699 10195 12705
rect 8613 12665 8625 12668
rect 8567 12659 8625 12665
rect 10137 12665 10149 12699
rect 10183 12696 10195 12699
rect 10686 12696 10692 12708
rect 10183 12668 10692 12696
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 13903 12699 13961 12705
rect 10836 12668 10881 12696
rect 10836 12656 10842 12668
rect 13903 12665 13915 12699
rect 13949 12696 13961 12699
rect 13998 12696 14004 12708
rect 13949 12668 14004 12696
rect 13949 12665 13961 12668
rect 13903 12659 13961 12665
rect 13998 12656 14004 12668
rect 14056 12696 14062 12708
rect 15289 12699 15347 12705
rect 15289 12696 15301 12699
rect 14056 12668 15301 12696
rect 14056 12656 14062 12668
rect 15289 12665 15301 12668
rect 15335 12665 15347 12699
rect 15289 12659 15347 12665
rect 15378 12656 15384 12708
rect 15436 12696 15442 12708
rect 15657 12699 15715 12705
rect 15657 12696 15669 12699
rect 15436 12668 15669 12696
rect 15436 12656 15442 12668
rect 15657 12665 15669 12668
rect 15703 12665 15715 12699
rect 15657 12659 15715 12665
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 15804 12668 15849 12696
rect 15804 12656 15810 12668
rect 16850 12656 16856 12708
rect 16908 12696 16914 12708
rect 17310 12696 17316 12708
rect 16908 12668 17316 12696
rect 16908 12656 16914 12668
rect 17310 12656 17316 12668
rect 17368 12696 17374 12708
rect 17405 12699 17463 12705
rect 17405 12696 17417 12699
rect 17368 12668 17417 12696
rect 17368 12656 17374 12668
rect 17405 12665 17417 12668
rect 17451 12665 17463 12699
rect 17405 12659 17463 12665
rect 17954 12656 17960 12708
rect 18012 12696 18018 12708
rect 18690 12696 18696 12708
rect 18012 12668 18696 12696
rect 18012 12656 18018 12668
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 18785 12699 18843 12705
rect 18785 12665 18797 12699
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 20349 12699 20407 12705
rect 20349 12665 20361 12699
rect 20395 12665 20407 12699
rect 20349 12659 20407 12665
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8478 12628 8484 12640
rect 7791 12600 8484 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9125 12631 9183 12637
rect 9125 12597 9137 12631
rect 9171 12628 9183 12631
rect 9306 12628 9312 12640
rect 9171 12600 9312 12628
rect 9171 12597 9183 12600
rect 9125 12591 9183 12597
rect 9306 12588 9312 12600
rect 9364 12588 9370 12640
rect 12066 12588 12072 12640
rect 12124 12628 12130 12640
rect 12161 12631 12219 12637
rect 12161 12628 12173 12631
rect 12124 12600 12173 12628
rect 12124 12588 12130 12600
rect 12161 12597 12173 12600
rect 12207 12597 12219 12631
rect 12161 12591 12219 12597
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 12989 12631 13047 12637
rect 12989 12628 13001 12631
rect 12676 12600 13001 12628
rect 12676 12588 12682 12600
rect 12989 12597 13001 12600
rect 13035 12628 13047 12631
rect 13170 12628 13176 12640
rect 13035 12600 13176 12628
rect 13035 12597 13047 12600
rect 12989 12591 13047 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 13320 12600 13369 12628
rect 13320 12588 13326 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 13357 12591 13415 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 15764 12628 15792 12656
rect 16577 12631 16635 12637
rect 16577 12628 16589 12631
rect 15764 12600 16589 12628
rect 16577 12597 16589 12600
rect 16623 12597 16635 12631
rect 17034 12628 17040 12640
rect 16995 12600 17040 12628
rect 16577 12591 16635 12597
rect 17034 12588 17040 12600
rect 17092 12588 17098 12640
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 18800 12628 18828 12659
rect 18656 12600 18828 12628
rect 18656 12588 18662 12600
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19518 12628 19524 12640
rect 19208 12600 19524 12628
rect 19208 12588 19214 12600
rect 19518 12588 19524 12600
rect 19576 12628 19582 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19576 12600 19993 12628
rect 19576 12588 19582 12600
rect 19981 12597 19993 12600
rect 20027 12628 20039 12631
rect 20364 12628 20392 12659
rect 20438 12656 20444 12708
rect 20496 12696 20502 12708
rect 23446 12696 23474 12736
rect 24581 12733 24593 12736
rect 24627 12764 24639 12767
rect 25133 12767 25191 12773
rect 25133 12764 25145 12767
rect 24627 12736 25145 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 25133 12733 25145 12736
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 20496 12668 23474 12696
rect 20496 12656 20502 12668
rect 21818 12628 21824 12640
rect 20027 12600 20392 12628
rect 21779 12600 21824 12628
rect 20027 12597 20039 12600
rect 19981 12591 20039 12597
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 22741 12631 22799 12637
rect 22741 12628 22753 12631
rect 22704 12600 22753 12628
rect 22704 12588 22710 12600
rect 22741 12597 22753 12600
rect 22787 12597 22799 12631
rect 23934 12628 23940 12640
rect 23847 12600 23940 12628
rect 22741 12591 22799 12597
rect 23934 12588 23940 12600
rect 23992 12628 23998 12640
rect 24210 12628 24216 12640
rect 23992 12600 24216 12628
rect 23992 12588 23998 12600
rect 24210 12588 24216 12600
rect 24268 12588 24274 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1673 12427 1731 12433
rect 1673 12393 1685 12427
rect 1719 12424 1731 12427
rect 1854 12424 1860 12436
rect 1719 12396 1860 12424
rect 1719 12393 1731 12396
rect 1673 12387 1731 12393
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 2004 12396 2053 12424
rect 2004 12384 2010 12396
rect 2041 12393 2053 12396
rect 2087 12424 2099 12427
rect 2314 12424 2320 12436
rect 2087 12396 2320 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 3510 12384 3516 12436
rect 3568 12384 3574 12436
rect 3694 12424 3700 12436
rect 3655 12396 3700 12424
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 7926 12424 7932 12436
rect 7887 12396 7932 12424
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8904 12396 9045 12424
rect 8904 12384 8910 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 9306 12384 9312 12436
rect 9364 12424 9370 12436
rect 9364 12396 10640 12424
rect 9364 12384 9370 12396
rect 2130 12316 2136 12368
rect 2188 12356 2194 12368
rect 2409 12359 2467 12365
rect 2409 12356 2421 12359
rect 2188 12328 2421 12356
rect 2188 12316 2194 12328
rect 2409 12325 2421 12328
rect 2455 12325 2467 12359
rect 2409 12319 2467 12325
rect 3528 12288 3556 12384
rect 5899 12359 5957 12365
rect 5899 12325 5911 12359
rect 5945 12356 5957 12359
rect 5994 12356 6000 12368
rect 5945 12328 6000 12356
rect 5945 12325 5957 12328
rect 5899 12319 5957 12325
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 7558 12316 7564 12368
rect 7616 12356 7622 12368
rect 8113 12359 8171 12365
rect 8113 12356 8125 12359
rect 7616 12328 8125 12356
rect 7616 12316 7622 12328
rect 8113 12325 8125 12328
rect 8159 12325 8171 12359
rect 8113 12319 8171 12325
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 9324 12356 9352 12384
rect 8260 12328 9352 12356
rect 8260 12316 8266 12328
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10612 12365 10640 12396
rect 10962 12384 10968 12436
rect 11020 12424 11026 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11020 12396 11805 12424
rect 11020 12384 11026 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 13357 12427 13415 12433
rect 13357 12393 13369 12427
rect 13403 12424 13415 12427
rect 14277 12427 14335 12433
rect 13403 12396 13768 12424
rect 13403 12393 13415 12396
rect 13357 12387 13415 12393
rect 10505 12359 10563 12365
rect 10505 12356 10517 12359
rect 10192 12328 10517 12356
rect 10192 12316 10198 12328
rect 10505 12325 10517 12328
rect 10551 12325 10563 12359
rect 10505 12319 10563 12325
rect 10597 12359 10655 12365
rect 10597 12325 10609 12359
rect 10643 12356 10655 12359
rect 11422 12356 11428 12368
rect 10643 12328 11428 12356
rect 10643 12325 10655 12328
rect 10597 12319 10655 12325
rect 11422 12316 11428 12328
rect 11480 12316 11486 12368
rect 13740 12356 13768 12396
rect 14277 12393 14289 12427
rect 14323 12424 14335 12427
rect 17862 12424 17868 12436
rect 14323 12396 17868 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 13998 12356 14004 12368
rect 13740 12328 14004 12356
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 3694 12288 3700 12300
rect 3528 12260 3700 12288
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4982 12288 4988 12300
rect 4111 12260 4988 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12288 5319 12291
rect 5350 12288 5356 12300
rect 5307 12260 5356 12288
rect 5307 12257 5319 12260
rect 5261 12251 5319 12257
rect 5350 12248 5356 12260
rect 5408 12288 5414 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 5408 12260 6469 12288
rect 5408 12248 5414 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 8846 12288 8852 12300
rect 8803 12260 8852 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 8846 12248 8852 12260
rect 8904 12288 8910 12300
rect 9582 12288 9588 12300
rect 8904 12260 9588 12288
rect 8904 12248 8910 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 11882 12248 11888 12300
rect 11940 12288 11946 12300
rect 12012 12291 12070 12297
rect 12012 12288 12024 12291
rect 11940 12260 12024 12288
rect 11940 12248 11946 12260
rect 12012 12257 12024 12260
rect 12058 12257 12070 12291
rect 12012 12251 12070 12257
rect 13538 12248 13544 12300
rect 13596 12288 13602 12300
rect 14292 12288 14320 12387
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18693 12427 18751 12433
rect 18693 12393 18705 12427
rect 18739 12424 18751 12427
rect 18874 12424 18880 12436
rect 18739 12396 18880 12424
rect 18739 12393 18751 12396
rect 18693 12387 18751 12393
rect 18874 12384 18880 12396
rect 18932 12424 18938 12436
rect 18969 12427 19027 12433
rect 18969 12424 18981 12427
rect 18932 12396 18981 12424
rect 18932 12384 18938 12396
rect 18969 12393 18981 12396
rect 19015 12393 19027 12427
rect 20714 12424 20720 12436
rect 20675 12396 20720 12424
rect 18969 12387 19027 12393
rect 20714 12384 20720 12396
rect 20772 12384 20778 12436
rect 14458 12316 14464 12368
rect 14516 12356 14522 12368
rect 15378 12356 15384 12368
rect 14516 12328 15384 12356
rect 14516 12316 14522 12328
rect 15378 12316 15384 12328
rect 15436 12356 15442 12368
rect 15473 12359 15531 12365
rect 15473 12356 15485 12359
rect 15436 12328 15485 12356
rect 15436 12316 15442 12328
rect 15473 12325 15485 12328
rect 15519 12325 15531 12359
rect 15473 12319 15531 12325
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16390 12356 16396 12368
rect 16071 12328 16396 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16390 12316 16396 12328
rect 16448 12316 16454 12368
rect 17954 12316 17960 12368
rect 18012 12356 18018 12368
rect 18094 12359 18152 12365
rect 18094 12356 18106 12359
rect 18012 12328 18106 12356
rect 18012 12316 18018 12328
rect 18094 12325 18106 12328
rect 18140 12325 18152 12359
rect 18094 12319 18152 12325
rect 13596 12260 14320 12288
rect 13596 12248 13602 12260
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 19886 12297 19892 12300
rect 19337 12291 19395 12297
rect 19337 12288 19349 12291
rect 18748 12260 19349 12288
rect 18748 12248 18754 12260
rect 19337 12257 19349 12260
rect 19383 12257 19395 12291
rect 19864 12291 19892 12297
rect 19864 12288 19876 12291
rect 19799 12260 19876 12288
rect 19337 12251 19395 12257
rect 19864 12257 19876 12260
rect 19944 12288 19950 12300
rect 20070 12288 20076 12300
rect 19944 12260 20076 12288
rect 19864 12251 19892 12257
rect 19886 12248 19892 12251
rect 19944 12248 19950 12260
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21269 12291 21327 12297
rect 21269 12288 21281 12291
rect 21140 12260 21281 12288
rect 21140 12248 21146 12260
rect 21269 12257 21281 12260
rect 21315 12257 21327 12291
rect 23566 12288 23572 12300
rect 23527 12260 23572 12288
rect 21269 12251 21327 12257
rect 23566 12248 23572 12260
rect 23624 12248 23630 12300
rect 25041 12291 25099 12297
rect 25041 12257 25053 12291
rect 25087 12288 25099 12291
rect 25130 12288 25136 12300
rect 25087 12260 25136 12288
rect 25087 12257 25099 12260
rect 25041 12251 25099 12257
rect 25130 12248 25136 12260
rect 25188 12248 25194 12300
rect 2314 12220 2320 12232
rect 2275 12192 2320 12220
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 5534 12220 5540 12232
rect 5447 12192 5540 12220
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 6914 12220 6920 12232
rect 5592 12192 6920 12220
rect 5592 12180 5598 12192
rect 6914 12180 6920 12192
rect 6972 12180 6978 12232
rect 10686 12180 10692 12232
rect 10744 12220 10750 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10744 12192 10793 12220
rect 10744 12180 10750 12192
rect 10781 12189 10793 12192
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 12897 12223 12955 12229
rect 12897 12189 12909 12223
rect 12943 12220 12955 12223
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12943 12192 13001 12220
rect 12943 12189 12955 12192
rect 12897 12183 12955 12189
rect 12989 12189 13001 12192
rect 13035 12220 13047 12223
rect 13722 12220 13728 12232
rect 13035 12192 13728 12220
rect 13035 12189 13047 12192
rect 12989 12183 13047 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12220 15439 12223
rect 15470 12220 15476 12232
rect 15427 12192 15476 12220
rect 15427 12189 15439 12192
rect 15381 12183 15439 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 16574 12220 16580 12232
rect 15580 12192 16580 12220
rect 4246 12152 4252 12164
rect 4207 12124 4252 12152
rect 4246 12112 4252 12124
rect 4304 12112 4310 12164
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 9674 12152 9680 12164
rect 6788 12124 9680 12152
rect 6788 12112 6794 12124
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 9950 12112 9956 12164
rect 10008 12152 10014 12164
rect 12434 12152 12440 12164
rect 10008 12124 12440 12152
rect 10008 12112 10014 12124
rect 12434 12112 12440 12124
rect 12492 12112 12498 12164
rect 13078 12112 13084 12164
rect 13136 12152 13142 12164
rect 15580 12152 15608 12192
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17276 12192 17785 12220
rect 17276 12180 17282 12192
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 23532 12192 23577 12220
rect 23532 12180 23538 12192
rect 13136 12124 15608 12152
rect 13136 12112 13142 12124
rect 6564 12084 6592 12112
rect 8386 12084 8392 12096
rect 6564 12056 8392 12084
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 12115 12087 12173 12093
rect 12115 12053 12127 12087
rect 12161 12084 12173 12087
rect 12342 12084 12348 12096
rect 12161 12056 12348 12084
rect 12161 12053 12173 12056
rect 12115 12047 12173 12053
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13906 12084 13912 12096
rect 13867 12056 13912 12084
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15286 12084 15292 12096
rect 15151 12056 15292 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 16298 12084 16304 12096
rect 15804 12056 16304 12084
rect 15804 12044 15810 12056
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 19935 12087 19993 12093
rect 19935 12053 19947 12087
rect 19981 12084 19993 12087
rect 20898 12084 20904 12096
rect 19981 12056 20904 12084
rect 19981 12053 19993 12056
rect 19935 12047 19993 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 21450 12084 21456 12096
rect 21411 12056 21456 12084
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 25038 12044 25044 12096
rect 25096 12084 25102 12096
rect 25179 12087 25237 12093
rect 25179 12084 25191 12087
rect 25096 12056 25191 12084
rect 25096 12044 25102 12056
rect 25179 12053 25191 12056
rect 25225 12053 25237 12087
rect 25179 12047 25237 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2188 11852 2881 11880
rect 2188 11840 2194 11852
rect 2869 11849 2881 11852
rect 2915 11880 2927 11883
rect 3145 11883 3203 11889
rect 3145 11880 3157 11883
rect 2915 11852 3157 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3145 11849 3157 11852
rect 3191 11880 3203 11883
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3191 11852 3525 11880
rect 3191 11849 3203 11852
rect 3145 11843 3203 11849
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 3513 11843 3571 11849
rect 5261 11883 5319 11889
rect 5261 11849 5273 11883
rect 5307 11880 5319 11883
rect 5534 11880 5540 11892
rect 5307 11852 5540 11880
rect 5307 11849 5319 11852
rect 5261 11843 5319 11849
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 1857 11611 1915 11617
rect 1857 11577 1869 11611
rect 1903 11608 1915 11611
rect 2270 11611 2328 11617
rect 2270 11608 2282 11611
rect 1903 11580 2282 11608
rect 1903 11577 1915 11580
rect 1857 11571 1915 11577
rect 2270 11577 2282 11580
rect 2316 11608 2328 11611
rect 2958 11608 2964 11620
rect 2316 11580 2964 11608
rect 2316 11577 2328 11580
rect 2270 11571 2328 11577
rect 2958 11568 2964 11580
rect 3016 11568 3022 11620
rect 3528 11608 3556 11843
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 5994 11880 6000 11892
rect 5675 11852 6000 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6270 11880 6276 11892
rect 6231 11852 6276 11880
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8202 11880 8208 11892
rect 8159 11852 8208 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10229 11883 10287 11889
rect 10229 11880 10241 11883
rect 10192 11852 10241 11880
rect 10192 11840 10198 11852
rect 10229 11849 10241 11852
rect 10275 11849 10287 11883
rect 11422 11880 11428 11892
rect 11383 11852 11428 11880
rect 10229 11843 10287 11849
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 13446 11880 13452 11892
rect 13359 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11880 13510 11892
rect 13998 11880 14004 11892
rect 13504 11852 14004 11880
rect 13504 11840 13510 11852
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 15488 11852 17509 11880
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 6362 11812 6368 11824
rect 4212 11784 6368 11812
rect 4212 11772 4218 11784
rect 6362 11772 6368 11784
rect 6420 11812 6426 11824
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 6420 11784 6561 11812
rect 6420 11772 6426 11784
rect 6549 11781 6561 11784
rect 6595 11781 6607 11815
rect 6549 11775 6607 11781
rect 6822 11772 6828 11824
rect 6880 11812 6886 11824
rect 6880 11784 6960 11812
rect 6880 11772 6886 11784
rect 3786 11744 3792 11756
rect 3747 11716 3792 11744
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4065 11747 4123 11753
rect 4065 11744 4077 11747
rect 4028 11716 4077 11744
rect 4028 11704 4034 11716
rect 4065 11713 4077 11716
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 4430 11744 4436 11756
rect 4304 11716 4436 11744
rect 4304 11704 4310 11716
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 6932 11753 6960 11784
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 9364 11784 11008 11812
rect 9364 11772 9370 11784
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 7156 11716 7205 11744
rect 7156 11704 7162 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 10134 11744 10140 11756
rect 9088 11716 10140 11744
rect 9088 11704 9094 11716
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10192 11716 10517 11744
rect 10192 11704 10198 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 10744 11716 10793 11744
rect 10744 11704 10750 11716
rect 10781 11713 10793 11716
rect 10827 11713 10839 11747
rect 10980 11744 11008 11784
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 13538 11812 13544 11824
rect 11756 11784 13544 11812
rect 11756 11772 11762 11784
rect 13538 11772 13544 11784
rect 13596 11772 13602 11824
rect 14016 11812 14044 11840
rect 15488 11812 15516 11852
rect 17497 11849 17509 11852
rect 17543 11880 17555 11883
rect 17773 11883 17831 11889
rect 17773 11880 17785 11883
rect 17543 11852 17785 11880
rect 17543 11849 17555 11852
rect 17497 11843 17555 11849
rect 17773 11849 17785 11852
rect 17819 11880 17831 11883
rect 17954 11880 17960 11892
rect 17819 11852 17960 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 19150 11880 19156 11892
rect 19111 11852 19156 11880
rect 19150 11840 19156 11852
rect 19208 11840 19214 11892
rect 19426 11880 19432 11892
rect 19387 11852 19432 11880
rect 19426 11840 19432 11852
rect 19484 11880 19490 11892
rect 20162 11880 20168 11892
rect 19484 11852 20168 11880
rect 19484 11840 19490 11852
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 21082 11880 21088 11892
rect 21043 11852 21088 11880
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 21358 11880 21364 11892
rect 21319 11852 21364 11880
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23566 11880 23572 11892
rect 23523 11852 23572 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 23566 11840 23572 11852
rect 23624 11840 23630 11892
rect 25406 11880 25412 11892
rect 25367 11852 25412 11880
rect 25406 11840 25412 11852
rect 25464 11840 25470 11892
rect 14016 11784 15516 11812
rect 15562 11772 15568 11824
rect 15620 11812 15626 11824
rect 17402 11812 17408 11824
rect 15620 11784 17408 11812
rect 15620 11772 15626 11784
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 19886 11812 19892 11824
rect 19847 11784 19892 11812
rect 19886 11772 19892 11784
rect 19944 11772 19950 11824
rect 20622 11812 20628 11824
rect 20583 11784 20628 11812
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 21542 11772 21548 11824
rect 21600 11812 21606 11824
rect 21600 11784 21680 11812
rect 21600 11772 21606 11784
rect 12250 11744 12256 11756
rect 10980 11716 12256 11744
rect 10781 11707 10839 11713
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12529 11747 12587 11753
rect 12529 11713 12541 11747
rect 12575 11744 12587 11747
rect 12802 11744 12808 11756
rect 12575 11716 12808 11744
rect 12575 11713 12587 11716
rect 12529 11707 12587 11713
rect 12802 11704 12808 11716
rect 12860 11744 12866 11756
rect 13262 11744 13268 11756
rect 12860 11716 13268 11744
rect 12860 11704 12866 11716
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11744 15071 11747
rect 15286 11744 15292 11756
rect 15059 11716 15292 11744
rect 15059 11713 15071 11716
rect 15013 11707 15071 11713
rect 15286 11704 15292 11716
rect 15344 11744 15350 11756
rect 16022 11744 16028 11756
rect 15344 11716 16028 11744
rect 15344 11704 15350 11716
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16390 11744 16396 11756
rect 16351 11716 16396 11744
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 20073 11747 20131 11753
rect 20073 11744 20085 11747
rect 19392 11716 20085 11744
rect 19392 11704 19398 11716
rect 20073 11713 20085 11716
rect 20119 11744 20131 11747
rect 20254 11744 20260 11756
rect 20119 11716 20260 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20254 11704 20260 11716
rect 20312 11704 20318 11756
rect 21652 11753 21680 11784
rect 21637 11747 21695 11753
rect 21637 11713 21649 11747
rect 21683 11713 21695 11747
rect 21910 11744 21916 11756
rect 21871 11716 21916 11744
rect 21637 11707 21695 11713
rect 21910 11704 21916 11716
rect 21968 11704 21974 11756
rect 5788 11679 5846 11685
rect 5788 11645 5800 11679
rect 5834 11676 5846 11679
rect 6270 11676 6276 11688
rect 5834 11648 6276 11676
rect 5834 11645 5846 11648
rect 5788 11639 5846 11645
rect 6270 11636 6276 11648
rect 6328 11636 6334 11688
rect 8754 11676 8760 11688
rect 8667 11648 8760 11676
rect 8754 11636 8760 11648
rect 8812 11676 8818 11688
rect 8941 11679 8999 11685
rect 8941 11676 8953 11679
rect 8812 11648 8953 11676
rect 8812 11636 8818 11648
rect 8941 11645 8953 11648
rect 8987 11645 8999 11679
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 8941 11639 8999 11645
rect 12176 11648 12449 11676
rect 3881 11611 3939 11617
rect 3881 11608 3893 11611
rect 3528 11580 3893 11608
rect 3881 11577 3893 11580
rect 3927 11577 3939 11611
rect 3881 11571 3939 11577
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 7009 11611 7067 11617
rect 7009 11608 7021 11611
rect 6420 11580 7021 11608
rect 6420 11568 6426 11580
rect 7009 11577 7021 11580
rect 7055 11577 7067 11611
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 7009 11571 7067 11577
rect 9876 11580 10609 11608
rect 9876 11552 9904 11580
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 10597 11571 10655 11577
rect 937 11543 995 11549
rect 937 11509 949 11543
rect 983 11540 995 11543
rect 1210 11540 1216 11552
rect 983 11512 1216 11540
rect 983 11509 995 11512
rect 937 11503 995 11509
rect 1210 11500 1216 11512
rect 1268 11500 1274 11552
rect 4801 11543 4859 11549
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 4982 11540 4988 11552
rect 4847 11512 4988 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 5859 11543 5917 11549
rect 5859 11509 5871 11543
rect 5905 11540 5917 11543
rect 6454 11540 6460 11552
rect 5905 11512 6460 11540
rect 5905 11509 5917 11512
rect 5859 11503 5917 11509
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 9030 11500 9036 11552
rect 9088 11540 9094 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 9088 11512 9137 11540
rect 9088 11500 9094 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 9125 11503 9183 11509
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10778 11540 10784 11552
rect 10100 11512 10784 11540
rect 10100 11500 10106 11512
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 12176 11549 12204 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 12713 11679 12771 11685
rect 12713 11676 12725 11679
rect 12676 11648 12725 11676
rect 12676 11636 12682 11648
rect 12713 11645 12725 11648
rect 12759 11645 12771 11679
rect 12713 11639 12771 11645
rect 15746 11636 15752 11688
rect 15804 11636 15810 11688
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11676 18291 11679
rect 18874 11676 18880 11688
rect 18279 11648 18880 11676
rect 18279 11645 18291 11648
rect 18233 11639 18291 11645
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 23109 11679 23167 11685
rect 23109 11645 23121 11679
rect 23155 11676 23167 11679
rect 23750 11676 23756 11688
rect 23155 11648 23756 11676
rect 23155 11645 23167 11648
rect 23109 11639 23167 11645
rect 23750 11636 23756 11648
rect 23808 11636 23814 11688
rect 25222 11676 25228 11688
rect 25183 11648 25228 11676
rect 25222 11636 25228 11648
rect 25280 11676 25286 11688
rect 25777 11679 25835 11685
rect 25777 11676 25789 11679
rect 25280 11648 25789 11676
rect 25280 11636 25286 11648
rect 25777 11645 25789 11648
rect 25823 11645 25835 11679
rect 25777 11639 25835 11645
rect 14366 11608 14372 11620
rect 14327 11580 14372 11608
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 14461 11611 14519 11617
rect 14461 11577 14473 11611
rect 14507 11577 14519 11611
rect 15764 11608 15792 11636
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 15764 11580 15945 11608
rect 14461 11571 14519 11577
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 16025 11611 16083 11617
rect 16025 11577 16037 11611
rect 16071 11608 16083 11611
rect 16206 11608 16212 11620
rect 16071 11580 16212 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11848 11512 12173 11540
rect 11848 11500 11854 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12161 11503 12219 11509
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12308 11512 12909 11540
rect 12308 11500 12314 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 13998 11500 14004 11552
rect 14056 11540 14062 11552
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 14056 11512 14197 11540
rect 14056 11500 14062 11512
rect 14185 11509 14197 11512
rect 14231 11540 14243 11543
rect 14476 11540 14504 11571
rect 14231 11512 14504 11540
rect 15749 11543 15807 11549
rect 14231 11509 14243 11512
rect 14185 11503 14243 11509
rect 15749 11509 15761 11543
rect 15795 11540 15807 11543
rect 16040 11540 16068 11571
rect 16206 11568 16212 11580
rect 16264 11568 16270 11620
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 18554 11611 18612 11617
rect 18554 11608 18566 11611
rect 18012 11580 18566 11608
rect 18012 11568 18018 11580
rect 18554 11577 18566 11580
rect 18600 11608 18612 11611
rect 19518 11608 19524 11620
rect 18600 11580 19524 11608
rect 18600 11577 18612 11580
rect 18554 11571 18612 11577
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 21729 11611 21787 11617
rect 20220 11580 20265 11608
rect 20220 11568 20226 11580
rect 21729 11577 21741 11611
rect 21775 11577 21787 11611
rect 25130 11608 25136 11620
rect 25043 11580 25136 11608
rect 21729 11571 21787 11577
rect 15795 11512 16068 11540
rect 17129 11543 17187 11549
rect 15795 11509 15807 11512
rect 15749 11503 15807 11509
rect 17129 11509 17141 11543
rect 17175 11540 17187 11543
rect 17218 11540 17224 11552
rect 17175 11512 17224 11540
rect 17175 11509 17187 11512
rect 17129 11503 17187 11509
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 21358 11500 21364 11552
rect 21416 11540 21422 11552
rect 21744 11540 21772 11571
rect 25130 11568 25136 11580
rect 25188 11608 25194 11620
rect 27614 11608 27620 11620
rect 25188 11580 27620 11608
rect 25188 11568 25194 11580
rect 27614 11568 27620 11580
rect 27672 11568 27678 11620
rect 24118 11540 24124 11552
rect 21416 11512 21772 11540
rect 24079 11512 24124 11540
rect 21416 11500 21422 11512
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 2314 11336 2320 11348
rect 1443 11308 2320 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5074 11336 5080 11348
rect 5031 11308 5080 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6362 11336 6368 11348
rect 6323 11308 6368 11336
rect 6362 11296 6368 11308
rect 6420 11296 6426 11348
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7558 11296 7564 11348
rect 7616 11336 7622 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7616 11308 7665 11336
rect 7616 11296 7622 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10192 11308 10241 11336
rect 10192 11296 10198 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 10229 11299 10287 11305
rect 11514 11296 11520 11348
rect 11572 11336 11578 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 11572 11308 12817 11336
rect 11572 11296 11578 11308
rect 12805 11305 12817 11308
rect 12851 11336 12863 11339
rect 12897 11339 12955 11345
rect 12897 11336 12909 11339
rect 12851 11308 12909 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 12897 11305 12909 11308
rect 12943 11305 12955 11339
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 12897 11299 12955 11305
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 14366 11336 14372 11348
rect 13786 11308 14372 11336
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 2593 11271 2651 11277
rect 2593 11268 2605 11271
rect 1820 11240 2605 11268
rect 1820 11228 1826 11240
rect 2593 11237 2605 11240
rect 2639 11237 2651 11271
rect 2593 11231 2651 11237
rect 3145 11271 3203 11277
rect 3145 11237 3157 11271
rect 3191 11268 3203 11271
rect 3970 11268 3976 11280
rect 3191 11240 3976 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 5807 11271 5865 11277
rect 5807 11268 5819 11271
rect 4212 11240 5819 11268
rect 4212 11228 4218 11240
rect 5807 11237 5819 11240
rect 5853 11268 5865 11271
rect 5994 11268 6000 11280
rect 5853 11240 6000 11268
rect 5853 11237 5865 11240
rect 5807 11231 5865 11237
rect 5994 11228 6000 11240
rect 6052 11228 6058 11280
rect 8199 11271 8257 11277
rect 8199 11237 8211 11271
rect 8245 11268 8257 11271
rect 8294 11268 8300 11280
rect 8245 11240 8300 11268
rect 8245 11237 8257 11240
rect 8199 11231 8257 11237
rect 8294 11228 8300 11240
rect 8352 11228 8358 11280
rect 10042 11228 10048 11280
rect 10100 11268 10106 11280
rect 10597 11271 10655 11277
rect 10597 11268 10609 11271
rect 10100 11240 10609 11268
rect 10100 11228 10106 11240
rect 10597 11237 10609 11240
rect 10643 11237 10655 11271
rect 10597 11231 10655 11237
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4614 11200 4620 11212
rect 4111 11172 4620 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5442 11200 5448 11212
rect 5403 11172 5448 11200
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 7800 11172 7849 11200
rect 7800 11160 7806 11172
rect 7837 11169 7849 11172
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 11974 11160 11980 11212
rect 12032 11200 12038 11212
rect 12104 11203 12162 11209
rect 12104 11200 12116 11203
rect 12032 11172 12116 11200
rect 12032 11160 12038 11172
rect 12104 11169 12116 11172
rect 12150 11169 12162 11203
rect 12104 11163 12162 11169
rect 12207 11203 12265 11209
rect 12207 11169 12219 11203
rect 12253 11200 12265 11203
rect 13786 11200 13814 11308
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 15105 11339 15163 11345
rect 15105 11305 15117 11339
rect 15151 11336 15163 11339
rect 15470 11336 15476 11348
rect 15151 11308 15476 11336
rect 15151 11305 15163 11308
rect 15105 11299 15163 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 17218 11336 17224 11348
rect 17179 11308 17224 11336
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 20254 11336 20260 11348
rect 20215 11308 20260 11336
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 22005 11339 22063 11345
rect 22005 11336 22017 11339
rect 21600 11308 22017 11336
rect 21600 11296 21606 11308
rect 22005 11305 22017 11308
rect 22051 11305 22063 11339
rect 22005 11299 22063 11305
rect 13906 11228 13912 11280
rect 13964 11268 13970 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 13964 11240 15669 11268
rect 13964 11228 13970 11240
rect 15657 11237 15669 11240
rect 15703 11237 15715 11271
rect 15657 11231 15715 11237
rect 17494 11228 17500 11280
rect 17552 11268 17558 11280
rect 17552 11240 18000 11268
rect 17552 11228 17558 11240
rect 12253 11172 13814 11200
rect 17405 11203 17463 11209
rect 12253 11169 12265 11172
rect 12207 11163 12265 11169
rect 17405 11169 17417 11203
rect 17451 11169 17463 11203
rect 17405 11163 17463 11169
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2501 11135 2559 11141
rect 2501 11132 2513 11135
rect 2372 11104 2513 11132
rect 2372 11092 2378 11104
rect 2501 11101 2513 11104
rect 2547 11132 2559 11135
rect 3418 11132 3424 11144
rect 2547 11104 3424 11132
rect 2547 11101 2559 11104
rect 2501 11095 2559 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 10502 11132 10508 11144
rect 6512 11104 10508 11132
rect 6512 11092 6518 11104
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10686 11092 10692 11144
rect 10744 11132 10750 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 10744 11104 10793 11132
rect 10744 11092 10750 11104
rect 10781 11101 10793 11104
rect 10827 11101 10839 11135
rect 10781 11095 10839 11101
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12851 11104 13093 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 13630 11092 13636 11144
rect 13688 11132 13694 11144
rect 15562 11132 15568 11144
rect 13688 11104 13814 11132
rect 15523 11104 15568 11132
rect 13688 11092 13694 11104
rect 382 11024 388 11076
rect 440 11064 446 11076
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 440 11036 4261 11064
rect 440 11024 446 11036
rect 4249 11033 4261 11036
rect 4295 11033 4307 11067
rect 4249 11027 4307 11033
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 9766 11064 9772 11076
rect 6420 11036 9772 11064
rect 6420 11024 6426 11036
rect 9766 11024 9772 11036
rect 9824 11024 9830 11076
rect 13786 11064 13814 11104
rect 15562 11092 15568 11104
rect 15620 11092 15626 11144
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 17420 11132 17448 11163
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 17862 11200 17868 11212
rect 17644 11172 17868 11200
rect 17644 11160 17650 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 17972 11209 18000 11240
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 21177 11271 21235 11277
rect 21177 11268 21189 11271
rect 20772 11240 21189 11268
rect 20772 11228 20778 11240
rect 21177 11237 21189 11240
rect 21223 11237 21235 11271
rect 21177 11231 21235 11237
rect 21729 11271 21787 11277
rect 21729 11237 21741 11271
rect 21775 11268 21787 11271
rect 21910 11268 21916 11280
rect 21775 11240 21916 11268
rect 21775 11237 21787 11240
rect 21729 11231 21787 11237
rect 21910 11228 21916 11240
rect 21968 11228 21974 11280
rect 17957 11203 18015 11209
rect 17957 11169 17969 11203
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11200 18567 11203
rect 18966 11200 18972 11212
rect 18555 11172 18972 11200
rect 18555 11169 18567 11172
rect 18509 11163 18567 11169
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 19864 11203 19922 11209
rect 19864 11169 19876 11203
rect 19910 11200 19922 11203
rect 20438 11200 20444 11212
rect 19910 11172 20444 11200
rect 19910 11169 19922 11172
rect 19864 11163 19922 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 22002 11160 22008 11212
rect 22060 11200 22066 11212
rect 22592 11203 22650 11209
rect 22592 11200 22604 11203
rect 22060 11172 22604 11200
rect 22060 11160 22066 11172
rect 22592 11169 22604 11172
rect 22638 11169 22650 11203
rect 22592 11163 22650 11169
rect 23106 11160 23112 11212
rect 23164 11200 23170 11212
rect 23845 11203 23903 11209
rect 23845 11200 23857 11203
rect 23164 11172 23857 11200
rect 23164 11160 23170 11172
rect 23845 11169 23857 11172
rect 23891 11169 23903 11203
rect 23845 11163 23903 11169
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11200 25375 11203
rect 25406 11200 25412 11212
rect 25363 11172 25412 11200
rect 25363 11169 25375 11172
rect 25317 11163 25375 11169
rect 25406 11160 25412 11172
rect 25464 11160 25470 11212
rect 18138 11132 18144 11144
rect 17420 11104 18144 11132
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20956 11104 21097 11132
rect 20956 11092 20962 11104
rect 21085 11101 21097 11104
rect 21131 11132 21143 11135
rect 22462 11132 22468 11144
rect 21131 11104 22468 11132
rect 21131 11101 21143 11104
rect 21085 11095 21143 11101
rect 22462 11092 22468 11104
rect 22520 11092 22526 11144
rect 23290 11092 23296 11144
rect 23348 11132 23354 11144
rect 23753 11135 23811 11141
rect 23753 11132 23765 11135
rect 23348 11104 23765 11132
rect 23348 11092 23354 11104
rect 23753 11101 23765 11104
rect 23799 11132 23811 11135
rect 24026 11132 24032 11144
rect 23799 11104 24032 11132
rect 23799 11101 23811 11104
rect 23753 11095 23811 11101
rect 24026 11092 24032 11104
rect 24084 11092 24090 11144
rect 13786 11036 15792 11064
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 1857 10999 1915 11005
rect 1857 10996 1869 10999
rect 1820 10968 1869 10996
rect 1820 10956 1826 10968
rect 1857 10965 1869 10968
rect 1903 10965 1915 10999
rect 1857 10959 1915 10965
rect 6086 10956 6092 11008
rect 6144 10996 6150 11008
rect 6914 10996 6920 11008
rect 6144 10968 6920 10996
rect 6144 10956 6150 10968
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 8757 10999 8815 11005
rect 8757 10965 8769 10999
rect 8803 10996 8815 10999
rect 9953 10999 10011 11005
rect 9953 10996 9965 10999
rect 8803 10968 9965 10996
rect 8803 10965 8815 10968
rect 8757 10959 8815 10965
rect 9953 10965 9965 10968
rect 9999 10996 10011 10999
rect 10042 10996 10048 11008
rect 9999 10968 10048 10996
rect 9999 10965 10011 10968
rect 9953 10959 10011 10965
rect 10042 10956 10048 10968
rect 10100 10956 10106 11008
rect 12621 10999 12679 11005
rect 12621 10965 12633 10999
rect 12667 10996 12679 10999
rect 12802 10996 12808 11008
rect 12667 10968 12808 10996
rect 12667 10965 12679 10968
rect 12621 10959 12679 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 13722 10956 13728 11008
rect 13780 10996 13786 11008
rect 14001 10999 14059 11005
rect 14001 10996 14013 10999
rect 13780 10968 14013 10996
rect 13780 10956 13786 10968
rect 14001 10965 14013 10968
rect 14047 10996 14059 10999
rect 14090 10996 14096 11008
rect 14047 10968 14096 10996
rect 14047 10965 14059 10968
rect 14001 10959 14059 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 15764 10996 15792 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 25455 11067 25513 11073
rect 25455 11064 25467 11067
rect 15896 11036 25467 11064
rect 15896 11024 15902 11036
rect 25455 11033 25467 11036
rect 25501 11033 25513 11067
rect 25455 11027 25513 11033
rect 17954 10996 17960 11008
rect 15764 10968 17960 10996
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 18874 10996 18880 11008
rect 18835 10968 18880 10996
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 19334 10996 19340 11008
rect 19295 10968 19340 10996
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 19935 10999 19993 11005
rect 19935 10965 19947 10999
rect 19981 10996 19993 10999
rect 20162 10996 20168 11008
rect 19981 10968 20168 10996
rect 19981 10965 19993 10968
rect 19935 10959 19993 10965
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 20254 10956 20260 11008
rect 20312 10996 20318 11008
rect 22695 10999 22753 11005
rect 22695 10996 22707 10999
rect 20312 10968 22707 10996
rect 20312 10956 20318 10968
rect 22695 10965 22707 10968
rect 22741 10965 22753 10999
rect 22695 10959 22753 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2958 10792 2964 10804
rect 2919 10764 2964 10792
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 5442 10752 5448 10804
rect 5500 10792 5506 10804
rect 6273 10795 6331 10801
rect 6273 10792 6285 10795
rect 5500 10764 6285 10792
rect 5500 10752 5506 10764
rect 6273 10761 6285 10764
rect 6319 10761 6331 10795
rect 6273 10755 6331 10761
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8294 10792 8300 10804
rect 7975 10764 8300 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8294 10752 8300 10764
rect 8352 10792 8358 10804
rect 9309 10795 9367 10801
rect 9309 10792 9321 10795
rect 8352 10764 9321 10792
rect 8352 10752 8358 10764
rect 9309 10761 9321 10764
rect 9355 10761 9367 10795
rect 9309 10755 9367 10761
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 11241 10795 11299 10801
rect 11241 10792 11253 10795
rect 10560 10764 11253 10792
rect 10560 10752 10566 10764
rect 11241 10761 11253 10764
rect 11287 10761 11299 10795
rect 13998 10792 14004 10804
rect 13959 10764 14004 10792
rect 11241 10755 11299 10761
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 15930 10792 15936 10804
rect 15344 10764 15936 10792
rect 15344 10752 15350 10764
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 17494 10792 17500 10804
rect 17455 10764 17500 10792
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 17865 10795 17923 10801
rect 17865 10792 17877 10795
rect 17736 10764 17877 10792
rect 17736 10752 17742 10764
rect 17865 10761 17877 10764
rect 17911 10792 17923 10795
rect 18138 10792 18144 10804
rect 17911 10764 18144 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 19518 10752 19524 10804
rect 19576 10792 19582 10804
rect 19613 10795 19671 10801
rect 19613 10792 19625 10795
rect 19576 10764 19625 10792
rect 19576 10752 19582 10764
rect 19613 10761 19625 10764
rect 19659 10761 19671 10795
rect 20714 10792 20720 10804
rect 20675 10764 20720 10792
rect 19613 10755 19671 10761
rect 20714 10752 20720 10764
rect 20772 10792 20778 10804
rect 20993 10795 21051 10801
rect 20993 10792 21005 10795
rect 20772 10764 21005 10792
rect 20772 10752 20778 10764
rect 20993 10761 21005 10764
rect 21039 10761 21051 10795
rect 20993 10755 21051 10761
rect 21082 10752 21088 10804
rect 21140 10792 21146 10804
rect 21361 10795 21419 10801
rect 21361 10792 21373 10795
rect 21140 10764 21373 10792
rect 21140 10752 21146 10764
rect 21361 10761 21373 10764
rect 21407 10761 21419 10795
rect 21361 10755 21419 10761
rect 4798 10684 4804 10736
rect 4856 10724 4862 10736
rect 6963 10727 7021 10733
rect 4856 10696 6224 10724
rect 4856 10684 4862 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 1854 10656 1860 10668
rect 1719 10628 1860 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2590 10656 2596 10668
rect 2363 10628 2596 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2590 10616 2596 10628
rect 2648 10616 2654 10668
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10656 3203 10659
rect 3602 10656 3608 10668
rect 3191 10628 3608 10656
rect 3191 10625 3203 10628
rect 3145 10619 3203 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5074 10656 5080 10668
rect 5031 10628 5080 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5074 10616 5080 10628
rect 5132 10616 5138 10668
rect 5166 10616 5172 10668
rect 5224 10656 5230 10668
rect 5261 10659 5319 10665
rect 5261 10656 5273 10659
rect 5224 10628 5273 10656
rect 5224 10616 5230 10628
rect 5261 10625 5273 10628
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 6196 10600 6224 10696
rect 6963 10693 6975 10727
rect 7009 10724 7021 10727
rect 13630 10724 13636 10736
rect 7009 10696 13636 10724
rect 7009 10693 7021 10696
rect 6963 10687 7021 10693
rect 13630 10684 13636 10696
rect 13688 10684 13694 10736
rect 14642 10684 14648 10736
rect 14700 10724 14706 10736
rect 15746 10724 15752 10736
rect 14700 10696 15752 10724
rect 14700 10684 14706 10696
rect 15746 10684 15752 10696
rect 15804 10684 15810 10736
rect 16022 10724 16028 10736
rect 15983 10696 16028 10724
rect 16022 10684 16028 10696
rect 16080 10684 16086 10736
rect 16390 10684 16396 10736
rect 16448 10724 16454 10736
rect 18693 10727 18751 10733
rect 18693 10724 18705 10727
rect 16448 10696 18705 10724
rect 16448 10684 16454 10696
rect 18693 10693 18705 10696
rect 18739 10693 18751 10727
rect 18693 10687 18751 10693
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 8113 10659 8171 10665
rect 8113 10656 8125 10659
rect 8076 10628 8125 10656
rect 8076 10616 8082 10628
rect 8113 10625 8125 10628
rect 8159 10656 8171 10659
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 8159 10628 9689 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 10192 10628 10241 10656
rect 10192 10616 10198 10628
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 11974 10616 11980 10668
rect 12032 10656 12038 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 12032 10628 12081 10656
rect 12032 10616 12038 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13081 10659 13139 10665
rect 13081 10656 13093 10659
rect 13044 10628 13093 10656
rect 13044 10616 13050 10628
rect 13081 10625 13093 10628
rect 13127 10656 13139 10659
rect 14277 10659 14335 10665
rect 14277 10656 14289 10659
rect 13127 10628 14289 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 14277 10625 14289 10628
rect 14323 10625 14335 10659
rect 14277 10619 14335 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15562 10656 15568 10668
rect 15335 10628 15568 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 15562 10616 15568 10628
rect 15620 10656 15626 10668
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 15620 10628 16957 10656
rect 15620 10616 15626 10628
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 19334 10656 19340 10668
rect 18187 10628 19340 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 19334 10616 19340 10628
rect 19392 10616 19398 10668
rect 4065 10591 4123 10597
rect 4065 10588 4077 10591
rect 2608 10560 4077 10588
rect 1762 10520 1768 10532
rect 1723 10492 1768 10520
rect 1762 10480 1768 10492
rect 1820 10480 1826 10532
rect 1780 10452 1808 10480
rect 2608 10461 2636 10560
rect 4065 10557 4077 10560
rect 4111 10588 4123 10591
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4111 10560 4721 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 2958 10480 2964 10532
rect 3016 10520 3022 10532
rect 3466 10523 3524 10529
rect 3466 10520 3478 10523
rect 3016 10492 3478 10520
rect 3016 10480 3022 10492
rect 3466 10489 3478 10492
rect 3512 10520 3524 10523
rect 4154 10520 4160 10532
rect 3512 10492 4160 10520
rect 3512 10489 3524 10492
rect 3466 10483 3524 10489
rect 4154 10480 4160 10492
rect 4212 10480 4218 10532
rect 2593 10455 2651 10461
rect 2593 10452 2605 10455
rect 1780 10424 2605 10452
rect 2593 10421 2605 10424
rect 2639 10421 2651 10455
rect 2593 10415 2651 10421
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4614 10452 4620 10464
rect 4479 10424 4620 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4724 10452 4752 10551
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6860 10591 6918 10597
rect 6860 10588 6872 10591
rect 6236 10560 6872 10588
rect 6236 10548 6242 10560
rect 6860 10557 6872 10560
rect 6906 10588 6918 10591
rect 7285 10591 7343 10597
rect 7285 10588 7297 10591
rect 6906 10560 7297 10588
rect 6906 10557 6918 10560
rect 6860 10551 6918 10557
rect 7285 10557 7297 10560
rect 7331 10557 7343 10591
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 7285 10551 7343 10557
rect 19260 10560 19809 10588
rect 5077 10523 5135 10529
rect 5077 10489 5089 10523
rect 5123 10489 5135 10523
rect 5994 10520 6000 10532
rect 5907 10492 6000 10520
rect 5077 10483 5135 10489
rect 5092 10452 5120 10483
rect 5994 10480 6000 10492
rect 6052 10520 6058 10532
rect 8294 10520 8300 10532
rect 6052 10492 8300 10520
rect 6052 10480 6058 10492
rect 8294 10480 8300 10492
rect 8352 10520 8358 10532
rect 8434 10523 8492 10529
rect 8434 10520 8446 10523
rect 8352 10492 8446 10520
rect 8352 10480 8358 10492
rect 8434 10489 8446 10492
rect 8480 10489 8492 10523
rect 9950 10520 9956 10532
rect 9911 10492 9956 10520
rect 8434 10483 8492 10489
rect 9950 10480 9956 10492
rect 10008 10480 10014 10532
rect 10042 10480 10048 10532
rect 10100 10520 10106 10532
rect 10965 10523 11023 10529
rect 10100 10492 10193 10520
rect 10100 10480 10106 10492
rect 10965 10489 10977 10523
rect 11011 10520 11023 10523
rect 11330 10520 11336 10532
rect 11011 10492 11336 10520
rect 11011 10489 11023 10492
rect 10965 10483 11023 10489
rect 4724 10424 5120 10452
rect 8202 10412 8208 10464
rect 8260 10452 8266 10464
rect 9033 10455 9091 10461
rect 9033 10452 9045 10455
rect 8260 10424 9045 10452
rect 8260 10412 8266 10424
rect 9033 10421 9045 10424
rect 9079 10421 9091 10455
rect 10060 10452 10088 10480
rect 10980 10452 11008 10483
rect 11330 10480 11336 10492
rect 11388 10480 11394 10532
rect 15102 10480 15108 10532
rect 15160 10520 15166 10532
rect 15473 10523 15531 10529
rect 15473 10520 15485 10523
rect 15160 10492 15485 10520
rect 15160 10480 15166 10492
rect 15473 10489 15485 10492
rect 15519 10489 15531 10523
rect 15473 10483 15531 10489
rect 15565 10523 15623 10529
rect 15565 10489 15577 10523
rect 15611 10520 15623 10523
rect 16485 10523 16543 10529
rect 16485 10520 16497 10523
rect 15611 10492 16497 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 16485 10489 16497 10492
rect 16531 10520 16543 10523
rect 18233 10523 18291 10529
rect 18233 10520 18245 10523
rect 16531 10492 18245 10520
rect 16531 10489 16543 10492
rect 16485 10483 16543 10489
rect 18233 10489 18245 10492
rect 18279 10489 18291 10523
rect 19058 10520 19064 10532
rect 18233 10483 18291 10489
rect 18616 10492 19064 10520
rect 10060 10424 11008 10452
rect 12989 10455 13047 10461
rect 9033 10415 9091 10421
rect 12989 10421 13001 10455
rect 13035 10452 13047 10455
rect 13446 10452 13452 10464
rect 13035 10424 13452 10452
rect 13035 10421 13047 10424
rect 12989 10415 13047 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14148 10424 14933 10452
rect 14148 10412 14154 10424
rect 14921 10421 14933 10424
rect 14967 10452 14979 10455
rect 15580 10452 15608 10483
rect 14967 10424 15608 10452
rect 16853 10455 16911 10461
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 18616 10452 18644 10492
rect 19058 10480 19064 10492
rect 19116 10480 19122 10532
rect 16899 10424 18644 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 19260 10461 19288 10560
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 19797 10551 19855 10557
rect 19518 10480 19524 10532
rect 19576 10520 19582 10532
rect 20118 10523 20176 10529
rect 20118 10520 20130 10523
rect 19576 10492 20130 10520
rect 19576 10480 19582 10492
rect 20118 10489 20130 10492
rect 20164 10520 20176 10523
rect 21082 10520 21088 10532
rect 20164 10492 21088 10520
rect 20164 10489 20176 10492
rect 20118 10483 20176 10489
rect 21082 10480 21088 10492
rect 21140 10480 21146 10532
rect 21376 10520 21404 10755
rect 22462 10752 22468 10804
rect 22520 10792 22526 10804
rect 22557 10795 22615 10801
rect 22557 10792 22569 10795
rect 22520 10764 22569 10792
rect 22520 10752 22526 10764
rect 22557 10761 22569 10764
rect 22603 10761 22615 10795
rect 23106 10792 23112 10804
rect 23067 10764 23112 10792
rect 22557 10755 22615 10761
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 24946 10792 24952 10804
rect 23532 10764 23577 10792
rect 24907 10764 24952 10792
rect 23532 10752 23538 10764
rect 24946 10752 24952 10764
rect 25004 10752 25010 10804
rect 24964 10724 24992 10752
rect 24044 10696 24992 10724
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10656 21695 10659
rect 21910 10656 21916 10668
rect 21683 10628 21916 10656
rect 21683 10625 21695 10628
rect 21637 10619 21695 10625
rect 21910 10616 21916 10628
rect 21968 10616 21974 10668
rect 24044 10665 24072 10696
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10625 24087 10659
rect 24302 10656 24308 10668
rect 24263 10628 24308 10656
rect 24029 10619 24087 10625
rect 24302 10616 24308 10628
rect 24360 10616 24366 10668
rect 25406 10656 25412 10668
rect 25319 10628 25412 10656
rect 25406 10616 25412 10628
rect 25464 10656 25470 10668
rect 27706 10656 27712 10668
rect 25464 10628 27712 10656
rect 25464 10616 25470 10628
rect 27706 10616 27712 10628
rect 27764 10616 27770 10668
rect 25568 10591 25626 10597
rect 25568 10557 25580 10591
rect 25614 10588 25626 10591
rect 25614 10560 26096 10588
rect 25614 10557 25626 10560
rect 25568 10551 25626 10557
rect 21729 10523 21787 10529
rect 21729 10520 21741 10523
rect 21376 10492 21741 10520
rect 21729 10489 21741 10492
rect 21775 10520 21787 10523
rect 21818 10520 21824 10532
rect 21775 10492 21824 10520
rect 21775 10489 21787 10492
rect 21729 10483 21787 10489
rect 21818 10480 21824 10492
rect 21876 10480 21882 10532
rect 22278 10520 22284 10532
rect 22239 10492 22284 10520
rect 22278 10480 22284 10492
rect 22336 10480 22342 10532
rect 24121 10523 24179 10529
rect 24121 10489 24133 10523
rect 24167 10489 24179 10523
rect 24121 10483 24179 10489
rect 19245 10455 19303 10461
rect 19245 10452 19257 10455
rect 19024 10424 19257 10452
rect 19024 10412 19030 10424
rect 19245 10421 19257 10424
rect 19291 10421 19303 10455
rect 19245 10415 19303 10421
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 24136 10452 24164 10483
rect 26068 10464 26096 10560
rect 23532 10424 24164 10452
rect 23532 10412 23538 10424
rect 24854 10412 24860 10464
rect 24912 10452 24918 10464
rect 25639 10455 25697 10461
rect 25639 10452 25651 10455
rect 24912 10424 25651 10452
rect 24912 10412 24918 10424
rect 25639 10421 25651 10424
rect 25685 10421 25697 10455
rect 26050 10452 26056 10464
rect 26011 10424 26056 10452
rect 25639 10415 25697 10421
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1535 10251 1593 10257
rect 1535 10248 1547 10251
rect 1452 10220 1547 10248
rect 1452 10208 1458 10220
rect 1535 10217 1547 10220
rect 1581 10217 1593 10251
rect 2314 10248 2320 10260
rect 2275 10220 2320 10248
rect 1535 10211 1593 10217
rect 2314 10208 2320 10220
rect 2372 10208 2378 10260
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 3602 10248 3608 10260
rect 3559 10220 3608 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5500 10220 5733 10248
rect 5500 10208 5506 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 7837 10211 7895 10217
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 15102 10248 15108 10260
rect 12400 10220 15108 10248
rect 12400 10208 12406 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 19058 10208 19064 10260
rect 19116 10248 19122 10260
rect 19153 10251 19211 10257
rect 19153 10248 19165 10251
rect 19116 10220 19165 10248
rect 19116 10208 19122 10220
rect 19153 10217 19165 10220
rect 19199 10217 19211 10251
rect 21818 10248 21824 10260
rect 21779 10220 21824 10248
rect 19153 10211 19211 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22097 10251 22155 10257
rect 22097 10248 22109 10251
rect 21968 10220 22109 10248
rect 21968 10208 21974 10220
rect 22097 10217 22109 10220
rect 22143 10217 22155 10251
rect 22097 10211 22155 10217
rect 24581 10251 24639 10257
rect 24581 10217 24593 10251
rect 24627 10248 24639 10251
rect 24946 10248 24952 10260
rect 24627 10220 24952 10248
rect 24627 10217 24639 10220
rect 24581 10211 24639 10217
rect 24946 10208 24952 10220
rect 25004 10208 25010 10260
rect 2498 10180 2504 10192
rect 2459 10152 2504 10180
rect 2498 10140 2504 10152
rect 2556 10140 2562 10192
rect 2593 10183 2651 10189
rect 2593 10149 2605 10183
rect 2639 10180 2651 10183
rect 2682 10180 2688 10192
rect 2639 10152 2688 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2682 10140 2688 10152
rect 2740 10140 2746 10192
rect 3786 10140 3792 10192
rect 3844 10180 3850 10192
rect 4157 10183 4215 10189
rect 4157 10180 4169 10183
rect 3844 10152 4169 10180
rect 3844 10140 3850 10152
rect 4157 10149 4169 10152
rect 4203 10149 4215 10183
rect 4157 10143 4215 10149
rect 4249 10183 4307 10189
rect 4249 10149 4261 10183
rect 4295 10180 4307 10183
rect 4430 10180 4436 10192
rect 4295 10152 4436 10180
rect 4295 10149 4307 10152
rect 4249 10143 4307 10149
rect 4430 10140 4436 10152
rect 4488 10140 4494 10192
rect 6086 10180 6092 10192
rect 5920 10152 6092 10180
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2314 10112 2320 10124
rect 1510 10084 2320 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 5920 10121 5948 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 8110 10180 8116 10192
rect 8071 10152 8116 10180
rect 8110 10140 8116 10152
rect 8168 10140 8174 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8757 10183 8815 10189
rect 8260 10152 8305 10180
rect 8260 10140 8266 10152
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 8846 10180 8852 10192
rect 8803 10152 8852 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 8846 10140 8852 10152
rect 8904 10180 8910 10192
rect 10134 10180 10140 10192
rect 8904 10152 10140 10180
rect 8904 10140 8910 10152
rect 10134 10140 10140 10152
rect 10192 10140 10198 10192
rect 11330 10180 11336 10192
rect 11291 10152 11336 10180
rect 11330 10140 11336 10152
rect 11388 10140 11394 10192
rect 11514 10140 11520 10192
rect 11572 10180 11578 10192
rect 11885 10183 11943 10189
rect 11885 10180 11897 10183
rect 11572 10152 11897 10180
rect 11572 10140 11578 10152
rect 11885 10149 11897 10152
rect 11931 10180 11943 10183
rect 12526 10180 12532 10192
rect 11931 10152 12532 10180
rect 11931 10149 11943 10152
rect 11885 10143 11943 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12710 10140 12716 10192
rect 12768 10180 12774 10192
rect 13173 10183 13231 10189
rect 13173 10180 13185 10183
rect 12768 10152 13185 10180
rect 12768 10140 12774 10152
rect 13173 10149 13185 10152
rect 13219 10180 13231 10183
rect 13446 10180 13452 10192
rect 13219 10152 13452 10180
rect 13219 10149 13231 10152
rect 13173 10143 13231 10149
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 13725 10183 13783 10189
rect 13725 10149 13737 10183
rect 13771 10180 13783 10183
rect 13906 10180 13912 10192
rect 13771 10152 13912 10180
rect 13771 10149 13783 10152
rect 13725 10143 13783 10149
rect 13906 10140 13912 10152
rect 13964 10140 13970 10192
rect 13998 10140 14004 10192
rect 14056 10180 14062 10192
rect 15378 10180 15384 10192
rect 14056 10152 15384 10180
rect 14056 10140 14062 10152
rect 15378 10140 15384 10152
rect 15436 10180 15442 10192
rect 15473 10183 15531 10189
rect 15473 10180 15485 10183
rect 15436 10152 15485 10180
rect 15436 10140 15442 10152
rect 15473 10149 15485 10152
rect 15519 10149 15531 10183
rect 15473 10143 15531 10149
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 18874 10180 18880 10192
rect 17552 10152 18276 10180
rect 18835 10152 18880 10180
rect 17552 10140 17558 10152
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6181 10115 6239 10121
rect 6181 10112 6193 10115
rect 6052 10084 6193 10112
rect 6052 10072 6058 10084
rect 6181 10081 6193 10084
rect 6227 10112 6239 10115
rect 7282 10112 7288 10124
rect 6227 10084 7288 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 9582 10112 9588 10124
rect 9456 10084 9588 10112
rect 9456 10072 9462 10084
rect 9582 10072 9588 10084
rect 9640 10112 9646 10124
rect 9712 10115 9770 10121
rect 9712 10112 9724 10115
rect 9640 10084 9724 10112
rect 9640 10072 9646 10084
rect 9712 10081 9724 10084
rect 9758 10081 9770 10115
rect 17678 10112 17684 10124
rect 17639 10084 17684 10112
rect 9712 10075 9770 10081
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 17862 10112 17868 10124
rect 17775 10084 17868 10112
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 18248 10121 18276 10152
rect 18874 10140 18880 10152
rect 18932 10140 18938 10192
rect 21082 10140 21088 10192
rect 21140 10180 21146 10192
rect 21222 10183 21280 10189
rect 21222 10180 21234 10183
rect 21140 10152 21234 10180
rect 21140 10140 21146 10152
rect 21222 10149 21234 10152
rect 21268 10149 21280 10183
rect 21222 10143 21280 10149
rect 23014 10140 23020 10192
rect 23072 10180 23078 10192
rect 23569 10183 23627 10189
rect 23569 10180 23581 10183
rect 23072 10152 23581 10180
rect 23072 10140 23078 10152
rect 23569 10149 23581 10152
rect 23615 10149 23627 10183
rect 23569 10143 23627 10149
rect 23658 10140 23664 10192
rect 23716 10180 23722 10192
rect 24213 10183 24271 10189
rect 23716 10152 23761 10180
rect 23716 10140 23722 10152
rect 24213 10149 24225 10183
rect 24259 10180 24271 10183
rect 24302 10180 24308 10192
rect 24259 10152 24308 10180
rect 24259 10149 24271 10152
rect 24213 10143 24271 10149
rect 18233 10115 18291 10121
rect 18233 10081 18245 10115
rect 18279 10112 18291 10115
rect 18598 10112 18604 10124
rect 18279 10084 18604 10112
rect 18279 10081 18291 10084
rect 18233 10075 18291 10081
rect 18598 10072 18604 10084
rect 18656 10072 18662 10124
rect 18782 10112 18788 10124
rect 18743 10084 18788 10112
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 19756 10115 19814 10121
rect 19756 10081 19768 10115
rect 19802 10112 19814 10115
rect 20346 10112 20352 10124
rect 19802 10084 20352 10112
rect 19802 10081 19814 10084
rect 19756 10075 19814 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 3145 10047 3203 10053
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3418 10044 3424 10056
rect 3191 10016 3424 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3418 10004 3424 10016
rect 3476 10044 3482 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 3476 10016 4445 10044
rect 3476 10004 3482 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 9950 10044 9956 10056
rect 8904 10016 9956 10044
rect 8904 10004 8910 10016
rect 9950 10004 9956 10016
rect 10008 10044 10014 10056
rect 10137 10047 10195 10053
rect 10137 10044 10149 10047
rect 10008 10016 10149 10044
rect 10008 10004 10014 10016
rect 10137 10013 10149 10016
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10044 11299 10047
rect 12250 10044 12256 10056
rect 11287 10016 12256 10044
rect 11287 10013 11299 10016
rect 11241 10007 11299 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 12713 9979 12771 9985
rect 12713 9976 12725 9979
rect 9185 9948 12725 9976
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 3142 9868 3148 9920
rect 3200 9908 3206 9920
rect 3602 9908 3608 9920
rect 3200 9880 3608 9908
rect 3200 9868 3206 9880
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5350 9908 5356 9920
rect 5307 9880 5356 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 9185 9908 9213 9948
rect 12713 9945 12725 9948
rect 12759 9976 12771 9979
rect 13648 9976 13676 10007
rect 14642 10004 14648 10056
rect 14700 10044 14706 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14700 10016 15393 10044
rect 14700 10004 14706 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 15470 10004 15476 10056
rect 15528 10044 15534 10056
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 15528 10016 15669 10044
rect 15528 10004 15534 10016
rect 15657 10013 15669 10016
rect 15703 10013 15715 10047
rect 17880 10044 17908 10072
rect 18874 10044 18880 10056
rect 15657 10007 15715 10013
rect 17144 10016 18880 10044
rect 12759 9948 13676 9976
rect 14185 9979 14243 9985
rect 12759 9945 12771 9948
rect 12713 9939 12771 9945
rect 14185 9945 14197 9979
rect 14231 9976 14243 9979
rect 14274 9976 14280 9988
rect 14231 9948 14280 9976
rect 14231 9945 14243 9948
rect 14185 9939 14243 9945
rect 14274 9936 14280 9948
rect 14332 9976 14338 9988
rect 15488 9976 15516 10004
rect 14332 9948 15516 9976
rect 14332 9936 14338 9948
rect 16206 9936 16212 9988
rect 16264 9976 16270 9988
rect 17144 9985 17172 10016
rect 18874 10004 18880 10016
rect 18932 10004 18938 10056
rect 19150 10004 19156 10056
rect 19208 10044 19214 10056
rect 19843 10047 19901 10053
rect 19843 10044 19855 10047
rect 19208 10016 19855 10044
rect 19208 10004 19214 10016
rect 19843 10013 19855 10016
rect 19889 10013 19901 10047
rect 20898 10044 20904 10056
rect 20859 10016 20904 10044
rect 19843 10007 19901 10013
rect 20898 10004 20904 10016
rect 20956 10004 20962 10056
rect 23198 10004 23204 10056
rect 23256 10044 23262 10056
rect 24228 10044 24256 10143
rect 24302 10140 24308 10152
rect 24360 10140 24366 10192
rect 25108 10115 25166 10121
rect 25108 10081 25120 10115
rect 25154 10112 25166 10115
rect 25314 10112 25320 10124
rect 25154 10084 25320 10112
rect 25154 10081 25166 10084
rect 25108 10075 25166 10081
rect 25314 10072 25320 10084
rect 25372 10072 25378 10124
rect 23256 10016 24256 10044
rect 23256 10004 23262 10016
rect 16761 9979 16819 9985
rect 16761 9976 16773 9979
rect 16264 9948 16773 9976
rect 16264 9936 16270 9948
rect 16761 9945 16773 9948
rect 16807 9976 16819 9979
rect 17129 9979 17187 9985
rect 17129 9976 17141 9979
rect 16807 9948 17141 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 17129 9945 17141 9948
rect 17175 9945 17187 9979
rect 18892 9976 18920 10004
rect 19521 9979 19579 9985
rect 19521 9976 19533 9979
rect 18892 9948 19533 9976
rect 17129 9939 17187 9945
rect 19521 9945 19533 9948
rect 19567 9945 19579 9979
rect 19521 9939 19579 9945
rect 23106 9936 23112 9988
rect 23164 9976 23170 9988
rect 23934 9976 23940 9988
rect 23164 9948 23940 9976
rect 23164 9936 23170 9948
rect 23934 9936 23940 9948
rect 23992 9936 23998 9988
rect 7708 9880 9213 9908
rect 7708 9868 7714 9880
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 9815 9911 9873 9917
rect 9815 9908 9827 9911
rect 9456 9880 9827 9908
rect 9456 9868 9462 9880
rect 9815 9877 9827 9880
rect 9861 9877 9873 9911
rect 10870 9908 10876 9920
rect 10831 9880 10876 9908
rect 9815 9871 9873 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 16298 9908 16304 9920
rect 16259 9880 16304 9908
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 20438 9908 20444 9920
rect 20303 9880 20444 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 20438 9868 20444 9880
rect 20496 9868 20502 9920
rect 22002 9868 22008 9920
rect 22060 9908 22066 9920
rect 22557 9911 22615 9917
rect 22557 9908 22569 9911
rect 22060 9880 22569 9908
rect 22060 9868 22066 9880
rect 22557 9877 22569 9880
rect 22603 9877 22615 9911
rect 22557 9871 22615 9877
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 23566 9908 23572 9920
rect 22980 9880 23572 9908
rect 22980 9868 22986 9880
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 24670 9868 24676 9920
rect 24728 9908 24734 9920
rect 25179 9911 25237 9917
rect 25179 9908 25191 9911
rect 24728 9880 25191 9908
rect 24728 9868 24734 9880
rect 25179 9877 25191 9880
rect 25225 9877 25237 9911
rect 25179 9871 25237 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 3142 9704 3148 9716
rect 1728 9676 3148 9704
rect 1728 9664 1734 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 3844 9676 4445 9704
rect 3844 9664 3850 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 5077 9707 5135 9713
rect 5077 9673 5089 9707
rect 5123 9704 5135 9707
rect 5994 9704 6000 9716
rect 5123 9676 6000 9704
rect 5123 9673 5135 9676
rect 5077 9667 5135 9673
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 5092 9636 5120 9667
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6181 9707 6239 9713
rect 6181 9704 6193 9707
rect 6144 9676 6193 9704
rect 6144 9664 6150 9676
rect 6181 9673 6193 9676
rect 6227 9673 6239 9707
rect 6181 9667 6239 9673
rect 8110 9664 8116 9716
rect 8168 9704 8174 9716
rect 8389 9707 8447 9713
rect 8389 9704 8401 9707
rect 8168 9676 8401 9704
rect 8168 9664 8174 9676
rect 8389 9673 8401 9676
rect 8435 9673 8447 9707
rect 9030 9704 9036 9716
rect 8991 9676 9036 9704
rect 8389 9667 8447 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9582 9664 9588 9716
rect 9640 9704 9646 9716
rect 10137 9707 10195 9713
rect 10137 9704 10149 9707
rect 9640 9676 10149 9704
rect 9640 9664 9646 9676
rect 10137 9673 10149 9676
rect 10183 9673 10195 9707
rect 10137 9667 10195 9673
rect 11330 9664 11336 9716
rect 11388 9704 11394 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11388 9676 11805 9704
rect 11388 9664 11394 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 13078 9704 13084 9716
rect 13039 9676 13084 9704
rect 11793 9667 11851 9673
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13449 9707 13507 9713
rect 13449 9673 13461 9707
rect 13495 9704 13507 9707
rect 13722 9704 13728 9716
rect 13495 9676 13728 9704
rect 13495 9673 13507 9676
rect 13449 9667 13507 9673
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 14642 9704 14648 9716
rect 14603 9676 14648 9704
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 16758 9664 16764 9716
rect 16816 9704 16822 9716
rect 18509 9707 18567 9713
rect 18509 9704 18521 9707
rect 16816 9676 18521 9704
rect 16816 9664 16822 9676
rect 18509 9673 18521 9676
rect 18555 9673 18567 9707
rect 18509 9667 18567 9673
rect 20993 9707 21051 9713
rect 20993 9673 21005 9707
rect 21039 9704 21051 9707
rect 21082 9704 21088 9716
rect 21039 9676 21088 9704
rect 21039 9673 21051 9676
rect 20993 9667 21051 9673
rect 9858 9636 9864 9648
rect 2004 9608 5120 9636
rect 8220 9608 9864 9636
rect 2004 9596 2010 9608
rect 8220 9580 8248 9608
rect 9858 9596 9864 9608
rect 9916 9636 9922 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 9916 9608 10609 9636
rect 9916 9596 9922 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 10597 9599 10655 9605
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9568 3111 9571
rect 3326 9568 3332 9580
rect 3099 9540 3332 9568
rect 3099 9537 3111 9540
rect 3053 9531 3111 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 5074 9568 5080 9580
rect 3476 9540 5080 9568
rect 3476 9528 3482 9540
rect 5074 9528 5080 9540
rect 5132 9568 5138 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5132 9540 5273 9568
rect 5132 9528 5138 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 7558 9568 7564 9580
rect 5261 9531 5319 9537
rect 7116 9540 7564 9568
rect 7116 9512 7144 9540
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9568 8171 9571
rect 8202 9568 8208 9580
rect 8159 9540 8208 9568
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 9214 9568 9220 9580
rect 9175 9540 9220 9568
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 937 9503 995 9509
rect 937 9469 949 9503
rect 983 9500 995 9503
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 983 9472 1685 9500
rect 983 9469 995 9472
rect 937 9463 995 9469
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1946 9500 1952 9512
rect 1907 9472 1952 9500
rect 1673 9463 1731 9469
rect 1688 9432 1716 9463
rect 1946 9460 1952 9472
rect 2004 9460 2010 9512
rect 3878 9460 3884 9512
rect 3936 9500 3942 9512
rect 4982 9500 4988 9512
rect 3936 9472 4988 9500
rect 3936 9460 3942 9472
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7098 9500 7104 9512
rect 6687 9472 7104 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7282 9500 7288 9512
rect 7243 9472 7288 9500
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 1688 9404 1992 9432
rect 1964 9376 1992 9404
rect 2590 9392 2596 9444
rect 2648 9432 2654 9444
rect 2869 9435 2927 9441
rect 2869 9432 2881 9435
rect 2648 9404 2881 9432
rect 2648 9392 2654 9404
rect 2869 9401 2881 9404
rect 2915 9432 2927 9435
rect 3145 9435 3203 9441
rect 3145 9432 3157 9435
rect 2915 9404 3157 9432
rect 2915 9401 2927 9404
rect 2869 9395 2927 9401
rect 3145 9401 3157 9404
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 5350 9392 5356 9444
rect 5408 9432 5414 9444
rect 5902 9432 5908 9444
rect 5408 9404 5453 9432
rect 5815 9404 5908 9432
rect 5408 9392 5414 9404
rect 5902 9392 5908 9404
rect 5960 9432 5966 9444
rect 7190 9432 7196 9444
rect 5960 9404 7196 9432
rect 5960 9392 5966 9404
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 9030 9392 9036 9444
rect 9088 9432 9094 9444
rect 9309 9435 9367 9441
rect 9309 9432 9321 9435
rect 9088 9404 9321 9432
rect 9088 9392 9094 9404
rect 9309 9401 9321 9404
rect 9355 9401 9367 9435
rect 9309 9395 9367 9401
rect 9861 9435 9919 9441
rect 9861 9401 9873 9435
rect 9907 9432 9919 9435
rect 10042 9432 10048 9444
rect 9907 9404 10048 9432
rect 9907 9401 9919 9404
rect 9861 9395 9919 9401
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 10612 9432 10640 9599
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 12713 9639 12771 9645
rect 12713 9636 12725 9639
rect 11020 9608 12725 9636
rect 11020 9596 11026 9608
rect 12713 9605 12725 9608
rect 12759 9605 12771 9639
rect 12713 9599 12771 9605
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 15565 9639 15623 9645
rect 15565 9636 15577 9639
rect 13964 9608 15577 9636
rect 13964 9596 13970 9608
rect 15565 9605 15577 9608
rect 15611 9636 15623 9639
rect 15657 9639 15715 9645
rect 15657 9636 15669 9639
rect 15611 9608 15669 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 15657 9605 15669 9608
rect 15703 9605 15715 9639
rect 15657 9599 15715 9605
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17129 9639 17187 9645
rect 17129 9636 17141 9639
rect 16632 9608 17141 9636
rect 16632 9596 16638 9608
rect 17129 9605 17141 9608
rect 17175 9636 17187 9639
rect 17678 9636 17684 9648
rect 17175 9608 17684 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 10870 9568 10876 9580
rect 10831 9540 10876 9568
rect 10870 9528 10876 9540
rect 10928 9528 10934 9580
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 13630 9568 13636 9580
rect 13591 9540 13636 9568
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 14274 9568 14280 9580
rect 14235 9540 14280 9568
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 15013 9571 15071 9577
rect 15013 9537 15025 9571
rect 15059 9568 15071 9571
rect 15930 9568 15936 9580
rect 15059 9540 15936 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16390 9568 16396 9580
rect 16351 9540 16396 9568
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 17494 9568 17500 9580
rect 17455 9540 17500 9568
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 18524 9512 18552 9667
rect 21082 9664 21088 9676
rect 21140 9664 21146 9716
rect 21450 9704 21456 9716
rect 21411 9676 21456 9704
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 22649 9707 22707 9713
rect 22649 9704 22661 9707
rect 21560 9676 22661 9704
rect 20898 9596 20904 9648
rect 20956 9636 20962 9648
rect 21560 9636 21588 9676
rect 22649 9673 22661 9676
rect 22695 9673 22707 9707
rect 23106 9704 23112 9716
rect 23067 9676 23112 9704
rect 22649 9667 22707 9673
rect 23106 9664 23112 9676
rect 23164 9664 23170 9716
rect 23477 9707 23535 9713
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 23566 9704 23572 9716
rect 23523 9676 23572 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 24026 9704 24032 9716
rect 23987 9676 24032 9704
rect 24026 9664 24032 9676
rect 24084 9664 24090 9716
rect 20956 9608 21588 9636
rect 20956 9596 20962 9608
rect 21634 9596 21640 9648
rect 21692 9636 21698 9648
rect 22278 9636 22284 9648
rect 21692 9608 21772 9636
rect 22239 9608 22284 9636
rect 21692 9596 21698 9608
rect 19058 9528 19064 9580
rect 19116 9568 19122 9580
rect 21744 9577 21772 9608
rect 22278 9596 22284 9608
rect 22336 9596 22342 9648
rect 21729 9571 21787 9577
rect 19116 9540 19932 9568
rect 19116 9528 19122 9540
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 13078 9500 13084 9512
rect 12575 9472 13084 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 17402 9460 17408 9512
rect 17460 9500 17466 9512
rect 17773 9503 17831 9509
rect 17773 9500 17785 9503
rect 17460 9472 17785 9500
rect 17460 9460 17466 9472
rect 17773 9469 17785 9472
rect 17819 9469 17831 9503
rect 18506 9500 18512 9512
rect 18419 9472 18512 9500
rect 17773 9463 17831 9469
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10612 9404 10977 9432
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 13722 9432 13728 9444
rect 13683 9404 13728 9432
rect 10965 9395 11023 9401
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 16025 9435 16083 9441
rect 16025 9432 16037 9435
rect 15611 9404 16037 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16025 9401 16037 9404
rect 16071 9432 16083 9435
rect 16298 9432 16304 9444
rect 16071 9404 16304 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 16298 9392 16304 9404
rect 16356 9392 16362 9444
rect 17788 9432 17816 9463
rect 18506 9460 18512 9472
rect 18564 9500 18570 9512
rect 18693 9503 18751 9509
rect 18693 9500 18705 9503
rect 18564 9472 18705 9500
rect 18564 9460 18570 9472
rect 18693 9469 18705 9472
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 18874 9460 18880 9512
rect 18932 9500 18938 9512
rect 19904 9509 19932 9540
rect 21729 9537 21741 9571
rect 21775 9537 21787 9571
rect 21729 9531 21787 9537
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 23440 9540 24317 9568
rect 23440 9528 23446 9540
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24578 9568 24584 9580
rect 24539 9540 24584 9568
rect 24305 9531 24363 9537
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18932 9472 19165 9500
rect 18932 9460 18938 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19521 9503 19579 9509
rect 19521 9469 19533 9503
rect 19567 9469 19579 9503
rect 19521 9463 19579 9469
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 19978 9500 19984 9512
rect 19935 9472 19984 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 19334 9432 19340 9444
rect 17788 9404 19340 9432
rect 18708 9376 18736 9404
rect 19334 9392 19340 9404
rect 19392 9432 19398 9444
rect 19536 9432 19564 9463
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 19392 9404 19564 9432
rect 19392 9392 19398 9404
rect 21450 9392 21456 9444
rect 21508 9432 21514 9444
rect 21821 9435 21879 9441
rect 21821 9432 21833 9435
rect 21508 9404 21833 9432
rect 21508 9392 21514 9404
rect 21821 9401 21833 9404
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 23290 9392 23296 9444
rect 23348 9432 23354 9444
rect 24397 9435 24455 9441
rect 23348 9404 24164 9432
rect 23348 9392 23354 9404
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 1946 9324 1952 9376
rect 2004 9324 2010 9376
rect 2038 9324 2044 9376
rect 2096 9364 2102 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2096 9336 2421 9364
rect 2096 9324 2102 9336
rect 2409 9333 2421 9336
rect 2455 9364 2467 9367
rect 2682 9364 2688 9376
rect 2455 9336 2688 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 4157 9367 4215 9373
rect 4157 9333 4169 9367
rect 4203 9364 4215 9367
rect 4430 9364 4436 9376
rect 4203 9336 4436 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6696 9336 6929 9364
rect 6696 9324 6702 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 12250 9364 12256 9376
rect 12211 9336 12256 9364
rect 6917 9327 6975 9333
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 14642 9364 14648 9376
rect 13136 9336 14648 9364
rect 13136 9324 13142 9336
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 18690 9324 18696 9376
rect 18748 9324 18754 9376
rect 18966 9364 18972 9376
rect 18927 9336 18972 9364
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 20346 9324 20352 9376
rect 20404 9364 20410 9376
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 20404 9336 20453 9364
rect 20404 9324 20410 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 24136 9364 24164 9404
rect 24397 9401 24409 9435
rect 24443 9401 24455 9435
rect 24397 9395 24455 9401
rect 24412 9364 24440 9395
rect 25314 9364 25320 9376
rect 24136 9336 24440 9364
rect 25275 9336 25320 9364
rect 20441 9327 20499 9333
rect 25314 9324 25320 9336
rect 25372 9324 25378 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2498 9120 2504 9172
rect 2556 9160 2562 9172
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2556 9132 2973 9160
rect 2556 9120 2562 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 3326 9160 3332 9172
rect 3287 9132 3332 9160
rect 2961 9123 3019 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 4890 9160 4896 9172
rect 3660 9132 4896 9160
rect 3660 9120 3666 9132
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 5074 9160 5080 9172
rect 5035 9132 5080 9160
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 5408 9132 6193 9160
rect 5408 9120 5414 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 7147 9163 7205 9169
rect 7147 9129 7159 9163
rect 7193 9160 7205 9163
rect 7650 9160 7656 9172
rect 7193 9132 7656 9160
rect 7193 9129 7205 9132
rect 7147 9123 7205 9129
rect 7650 9120 7656 9132
rect 7708 9120 7714 9172
rect 7834 9160 7840 9172
rect 7795 9132 7840 9160
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 9214 9160 9220 9172
rect 9175 9132 9220 9160
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 10183 9163 10241 9169
rect 10183 9129 10195 9163
rect 10229 9160 10241 9163
rect 13078 9160 13084 9172
rect 10229 9132 13084 9160
rect 10229 9129 10241 9132
rect 10183 9123 10241 9129
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 13688 9132 14197 9160
rect 13688 9120 13694 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 14185 9123 14243 9129
rect 14568 9132 16313 9160
rect 1854 9052 1860 9104
rect 1912 9092 1918 9104
rect 2086 9095 2144 9101
rect 2086 9092 2098 9095
rect 1912 9064 2098 9092
rect 1912 9052 1918 9064
rect 2086 9061 2098 9064
rect 2132 9061 2144 9095
rect 2086 9055 2144 9061
rect 2314 9052 2320 9104
rect 2372 9092 2378 9104
rect 3697 9095 3755 9101
rect 3697 9092 3709 9095
rect 2372 9064 3709 9092
rect 2372 9052 2378 9064
rect 3697 9061 3709 9064
rect 3743 9061 3755 9095
rect 3697 9055 3755 9061
rect 5623 9095 5681 9101
rect 5623 9061 5635 9095
rect 5669 9092 5681 9095
rect 5994 9092 6000 9104
rect 5669 9064 6000 9092
rect 5669 9061 5681 9064
rect 5623 9055 5681 9061
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2866 8956 2872 8968
rect 1811 8928 2872 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3712 8956 3740 9055
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 6917 9095 6975 9101
rect 6917 9061 6929 9095
rect 6963 9092 6975 9095
rect 7282 9092 7288 9104
rect 6963 9064 7288 9092
rect 6963 9061 6975 9064
rect 6917 9055 6975 9061
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7852 9092 7880 9120
rect 8113 9095 8171 9101
rect 8113 9092 8125 9095
rect 7852 9064 8125 9092
rect 8113 9061 8125 9064
rect 8159 9061 8171 9095
rect 8113 9055 8171 9061
rect 8205 9095 8263 9101
rect 8205 9061 8217 9095
rect 8251 9092 8263 9095
rect 8294 9092 8300 9104
rect 8251 9064 8300 9092
rect 8251 9061 8263 9064
rect 8205 9055 8263 9061
rect 8294 9052 8300 9064
rect 8352 9092 8358 9104
rect 8754 9092 8760 9104
rect 8352 9064 8760 9092
rect 8352 9052 8358 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 11419 9095 11477 9101
rect 11419 9061 11431 9095
rect 11465 9092 11477 9095
rect 11514 9092 11520 9104
rect 11465 9064 11520 9092
rect 11465 9061 11477 9064
rect 11419 9055 11477 9061
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 14568 9092 14596 9132
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 16942 9120 16948 9172
rect 17000 9160 17006 9172
rect 17862 9160 17868 9172
rect 17000 9132 17868 9160
rect 17000 9120 17006 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18049 9163 18107 9169
rect 18049 9129 18061 9163
rect 18095 9160 18107 9163
rect 18417 9163 18475 9169
rect 18417 9160 18429 9163
rect 18095 9132 18429 9160
rect 18095 9129 18107 9132
rect 18049 9123 18107 9129
rect 18417 9129 18429 9132
rect 18463 9160 18475 9163
rect 18782 9160 18788 9172
rect 18463 9132 18788 9160
rect 18463 9129 18475 9132
rect 18417 9123 18475 9129
rect 11808 9064 14596 9092
rect 16316 9064 16712 9092
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 4614 9024 4620 9036
rect 4111 8996 4620 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 4614 8984 4620 8996
rect 4672 9024 4678 9036
rect 5166 9024 5172 9036
rect 4672 8996 5172 9024
rect 4672 8984 4678 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 9024 5319 9027
rect 5442 9024 5448 9036
rect 5307 8996 5448 9024
rect 5307 8993 5319 8996
rect 5261 8987 5319 8993
rect 5442 8984 5448 8996
rect 5500 8984 5506 9036
rect 7076 9027 7134 9033
rect 7076 8993 7088 9027
rect 7122 9024 7134 9027
rect 7374 9024 7380 9036
rect 7122 8996 7380 9024
rect 7122 8993 7134 8996
rect 7076 8987 7134 8993
rect 7374 8984 7380 8996
rect 7432 8984 7438 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10080 9027 10138 9033
rect 10080 9024 10092 9027
rect 10008 8996 10092 9024
rect 10008 8984 10014 8996
rect 10080 8993 10092 8996
rect 10126 8993 10138 9027
rect 11054 9024 11060 9036
rect 10967 8996 11060 9024
rect 10080 8987 10138 8993
rect 11054 8984 11060 8996
rect 11112 9024 11118 9036
rect 11808 9024 11836 9064
rect 16316 9036 16344 9064
rect 11974 9024 11980 9036
rect 11112 8996 11836 9024
rect 11887 8996 11980 9024
rect 11112 8984 11118 8996
rect 11974 8984 11980 8996
rect 12032 9024 12038 9036
rect 13446 9024 13452 9036
rect 12032 8996 13452 9024
rect 12032 8984 12038 8996
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13906 9024 13912 9036
rect 13867 8996 13912 9024
rect 13906 8984 13912 8996
rect 13964 8984 13970 9036
rect 16298 8984 16304 9036
rect 16356 8984 16362 9036
rect 16485 9027 16543 9033
rect 16485 8993 16497 9027
rect 16531 9024 16543 9027
rect 16574 9024 16580 9036
rect 16531 8996 16580 9024
rect 16531 8993 16543 8996
rect 16485 8987 16543 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 16684 9033 16712 9064
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16942 8984 16948 9036
rect 17000 9024 17006 9036
rect 17126 9024 17132 9036
rect 17000 8996 17132 9024
rect 17000 8984 17006 8996
rect 17126 8984 17132 8996
rect 17184 8984 17190 9036
rect 17218 8984 17224 9036
rect 17276 9024 17282 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17276 8996 17601 9024
rect 17276 8984 17282 8996
rect 17589 8993 17601 8996
rect 17635 9024 17647 9027
rect 18064 9024 18092 9123
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 21082 9120 21088 9172
rect 21140 9160 21146 9172
rect 21634 9160 21640 9172
rect 21140 9132 21265 9160
rect 21595 9132 21640 9160
rect 21140 9120 21146 9132
rect 18800 9092 18828 9120
rect 19518 9092 19524 9104
rect 18800 9064 19524 9092
rect 19518 9052 19524 9064
rect 19576 9092 19582 9104
rect 19981 9095 20039 9101
rect 19576 9064 19748 9092
rect 19576 9052 19582 9064
rect 18506 9024 18512 9036
rect 17635 8996 18092 9024
rect 18467 8996 18512 9024
rect 17635 8993 17647 8996
rect 17589 8987 17647 8993
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 18969 9027 19027 9033
rect 18969 9024 18981 9027
rect 18932 8996 18981 9024
rect 18932 8984 18938 8996
rect 18969 8993 18981 8996
rect 19015 8993 19027 9027
rect 19334 9024 19340 9036
rect 19295 8996 19340 9024
rect 18969 8987 19027 8993
rect 5902 8956 5908 8968
rect 3712 8928 5908 8956
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9766 8956 9772 8968
rect 8803 8928 9772 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9766 8916 9772 8928
rect 9824 8956 9830 8968
rect 10597 8959 10655 8965
rect 10597 8956 10609 8959
rect 9824 8928 10609 8956
rect 9824 8916 9830 8928
rect 10597 8925 10609 8928
rect 10643 8956 10655 8959
rect 10686 8956 10692 8968
rect 10643 8928 10692 8956
rect 10643 8925 10655 8928
rect 10597 8919 10655 8925
rect 10686 8916 10692 8928
rect 10744 8916 10750 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 11204 8928 12817 8956
rect 11204 8916 11210 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 18138 8956 18144 8968
rect 14516 8928 18144 8956
rect 14516 8916 14522 8928
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 18984 8956 19012 8987
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19720 9033 19748 9064
rect 19981 9061 19993 9095
rect 20027 9092 20039 9095
rect 20898 9092 20904 9104
rect 20027 9064 20904 9092
rect 20027 9061 20039 9064
rect 19981 9055 20039 9061
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 21237 9092 21265 9132
rect 21634 9120 21640 9132
rect 21692 9120 21698 9172
rect 22922 9160 22928 9172
rect 22883 9132 22928 9160
rect 22922 9120 22928 9132
rect 22980 9120 22986 9172
rect 25498 9120 25504 9172
rect 25556 9169 25562 9172
rect 25556 9163 25605 9169
rect 25556 9129 25559 9163
rect 25593 9129 25605 9163
rect 25556 9123 25605 9129
rect 25556 9120 25562 9123
rect 22278 9092 22284 9104
rect 21237 9064 22284 9092
rect 22278 9052 22284 9064
rect 22336 9101 22342 9104
rect 22336 9095 22384 9101
rect 22336 9061 22338 9095
rect 22372 9061 22384 9095
rect 23106 9092 23112 9104
rect 22336 9055 22384 9061
rect 22480 9064 23112 9092
rect 22336 9052 22342 9055
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 8993 19763 9027
rect 19705 8987 19763 8993
rect 20717 9027 20775 9033
rect 20717 8993 20729 9027
rect 20763 9024 20775 9027
rect 21060 9027 21118 9033
rect 21060 9024 21072 9027
rect 20763 8996 21072 9024
rect 20763 8993 20775 8996
rect 20717 8987 20775 8993
rect 21060 8993 21072 8996
rect 21106 9024 21118 9027
rect 22480 9024 22508 9064
rect 23106 9052 23112 9064
rect 23164 9052 23170 9104
rect 23934 9052 23940 9104
rect 23992 9092 23998 9104
rect 24029 9095 24087 9101
rect 24029 9092 24041 9095
rect 23992 9064 24041 9092
rect 23992 9052 23998 9064
rect 24029 9061 24041 9064
rect 24075 9061 24087 9095
rect 24029 9055 24087 9061
rect 21106 8996 22508 9024
rect 21106 8993 21118 8996
rect 21060 8987 21118 8993
rect 22554 8984 22560 9036
rect 22612 9024 22618 9036
rect 23661 9027 23719 9033
rect 23661 9024 23673 9027
rect 22612 8996 23673 9024
rect 22612 8984 22618 8996
rect 23661 8993 23673 8996
rect 23707 8993 23719 9027
rect 23661 8987 23719 8993
rect 25476 9027 25534 9033
rect 25476 8993 25488 9027
rect 25522 9024 25534 9027
rect 25774 9024 25780 9036
rect 25522 8996 25780 9024
rect 25522 8993 25534 8996
rect 25476 8987 25534 8993
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 18984 8928 20269 8956
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20257 8919 20315 8925
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 20588 8928 22017 8956
rect 20588 8916 20594 8928
rect 22005 8925 22017 8928
rect 22051 8956 22063 8959
rect 22738 8956 22744 8968
rect 22051 8928 22744 8956
rect 22051 8925 22063 8928
rect 22005 8919 22063 8925
rect 22738 8916 22744 8928
rect 22796 8916 22802 8968
rect 23676 8956 23704 8987
rect 25774 8984 25780 8996
rect 25832 8984 25838 9036
rect 23937 8959 23995 8965
rect 23937 8956 23949 8959
rect 23676 8928 23949 8956
rect 23937 8925 23949 8928
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 24026 8916 24032 8968
rect 24084 8956 24090 8968
rect 24213 8959 24271 8965
rect 24213 8956 24225 8959
rect 24084 8928 24225 8956
rect 24084 8916 24090 8928
rect 24213 8925 24225 8928
rect 24259 8956 24271 8959
rect 24578 8956 24584 8968
rect 24259 8928 24584 8956
rect 24259 8925 24271 8928
rect 24213 8919 24271 8925
rect 24578 8916 24584 8928
rect 24636 8916 24642 8968
rect 3510 8848 3516 8900
rect 3568 8888 3574 8900
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3568 8860 4261 8888
rect 3568 8848 3574 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7834 8888 7840 8900
rect 7064 8860 7840 8888
rect 7064 8848 7070 8860
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 11882 8848 11888 8900
rect 11940 8888 11946 8900
rect 12437 8891 12495 8897
rect 12437 8888 12449 8891
rect 11940 8860 12449 8888
rect 11940 8848 11946 8860
rect 12437 8857 12449 8860
rect 12483 8888 12495 8891
rect 12526 8888 12532 8900
rect 12483 8860 12532 8888
rect 12483 8857 12495 8860
rect 12437 8851 12495 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 20346 8848 20352 8900
rect 20404 8888 20410 8900
rect 20404 8860 23474 8888
rect 20404 8848 20410 8860
rect 1673 8823 1731 8829
rect 1673 8789 1685 8823
rect 1719 8820 1731 8823
rect 1946 8820 1952 8832
rect 1719 8792 1952 8820
rect 1719 8789 1731 8792
rect 1673 8783 1731 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2682 8820 2688 8832
rect 2643 8792 2688 8820
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 15749 8823 15807 8829
rect 15749 8789 15761 8823
rect 15795 8820 15807 8823
rect 15838 8820 15844 8832
rect 15795 8792 15844 8820
rect 15795 8789 15807 8792
rect 15749 8783 15807 8789
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 16117 8823 16175 8829
rect 16117 8789 16129 8823
rect 16163 8820 16175 8823
rect 16298 8820 16304 8832
rect 16163 8792 16304 8820
rect 16163 8789 16175 8792
rect 16117 8783 16175 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 21131 8823 21189 8829
rect 21131 8789 21143 8823
rect 21177 8820 21189 8823
rect 22462 8820 22468 8832
rect 21177 8792 22468 8820
rect 21177 8789 21189 8792
rect 21131 8783 21189 8789
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 23446 8820 23474 8860
rect 24762 8848 24768 8900
rect 24820 8888 24826 8900
rect 25222 8888 25228 8900
rect 24820 8860 25228 8888
rect 24820 8848 24826 8860
rect 25222 8848 25228 8860
rect 25280 8848 25286 8900
rect 25406 8820 25412 8832
rect 23446 8792 25412 8820
rect 25406 8780 25412 8792
rect 25464 8780 25470 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 4341 8619 4399 8625
rect 4341 8585 4353 8619
rect 4387 8616 4399 8619
rect 4614 8616 4620 8628
rect 4387 8588 4620 8616
rect 4387 8585 4399 8588
rect 4341 8579 4399 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 5442 8616 5448 8628
rect 4755 8588 5448 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 7374 8576 7380 8628
rect 7432 8616 7438 8628
rect 7837 8619 7895 8625
rect 7837 8616 7849 8619
rect 7432 8588 7849 8616
rect 7432 8576 7438 8588
rect 7837 8585 7849 8588
rect 7883 8585 7895 8619
rect 8294 8616 8300 8628
rect 8255 8588 8300 8616
rect 7837 8579 7895 8585
rect 8294 8576 8300 8588
rect 8352 8616 8358 8628
rect 9769 8619 9827 8625
rect 9769 8616 9781 8619
rect 8352 8588 9781 8616
rect 8352 8576 8358 8588
rect 9769 8585 9781 8588
rect 9815 8616 9827 8619
rect 9858 8616 9864 8628
rect 9815 8588 9864 8616
rect 9815 8585 9827 8588
rect 9769 8579 9827 8585
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 11609 8619 11667 8625
rect 11609 8616 11621 8619
rect 11572 8588 11621 8616
rect 11572 8576 11578 8588
rect 11609 8585 11621 8588
rect 11655 8616 11667 8619
rect 12710 8616 12716 8628
rect 11655 8588 12716 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15378 8616 15384 8628
rect 15335 8588 15384 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15378 8576 15384 8588
rect 15436 8616 15442 8628
rect 15930 8616 15936 8628
rect 15436 8588 15936 8616
rect 15436 8576 15442 8588
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 16942 8616 16948 8628
rect 16899 8588 16948 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17218 8616 17224 8628
rect 17179 8588 17224 8616
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 18230 8616 18236 8628
rect 18191 8588 18236 8616
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 22278 8576 22284 8628
rect 22336 8616 22342 8628
rect 22373 8619 22431 8625
rect 22373 8616 22385 8619
rect 22336 8588 22385 8616
rect 22336 8576 22342 8588
rect 22373 8585 22385 8588
rect 22419 8616 22431 8619
rect 22554 8616 22560 8628
rect 22419 8588 22560 8616
rect 22419 8585 22431 8588
rect 22373 8579 22431 8585
rect 22554 8576 22560 8588
rect 22612 8576 22618 8628
rect 22738 8616 22744 8628
rect 22699 8588 22744 8616
rect 22738 8576 22744 8588
rect 22796 8576 22802 8628
rect 23477 8619 23535 8625
rect 23477 8585 23489 8619
rect 23523 8616 23535 8619
rect 23750 8616 23756 8628
rect 23523 8588 23756 8616
rect 23523 8585 23535 8588
rect 23477 8579 23535 8585
rect 23750 8576 23756 8588
rect 23808 8576 23814 8628
rect 23934 8576 23940 8628
rect 23992 8616 23998 8628
rect 24762 8616 24768 8628
rect 23992 8588 24768 8616
rect 23992 8576 23998 8588
rect 24762 8576 24768 8588
rect 24820 8616 24826 8628
rect 24857 8619 24915 8625
rect 24857 8616 24869 8619
rect 24820 8588 24869 8616
rect 24820 8576 24826 8588
rect 24857 8585 24869 8588
rect 24903 8585 24915 8619
rect 24857 8579 24915 8585
rect 25593 8619 25651 8625
rect 25593 8585 25605 8619
rect 25639 8616 25651 8619
rect 26142 8616 26148 8628
rect 25639 8588 26148 8616
rect 25639 8585 25651 8588
rect 25593 8579 25651 8585
rect 26142 8576 26148 8588
rect 26200 8576 26206 8628
rect 1302 8508 1308 8560
rect 1360 8548 1366 8560
rect 4062 8548 4068 8560
rect 1360 8520 4068 8548
rect 1360 8508 1366 8520
rect 4062 8508 4068 8520
rect 4120 8548 4126 8560
rect 9950 8548 9956 8560
rect 4120 8520 9956 8548
rect 4120 8508 4126 8520
rect 9950 8508 9956 8520
rect 10008 8548 10014 8560
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 10008 8520 10057 8548
rect 10008 8508 10014 8520
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 16390 8548 16396 8560
rect 16351 8520 16396 8548
rect 10045 8511 10103 8517
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17865 8551 17923 8557
rect 17865 8548 17877 8551
rect 17184 8520 17877 8548
rect 17184 8508 17190 8520
rect 17865 8517 17877 8520
rect 17911 8548 17923 8551
rect 18506 8548 18512 8560
rect 17911 8520 18512 8548
rect 17911 8517 17923 8520
rect 17865 8511 17923 8517
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 20809 8551 20867 8557
rect 20809 8548 20821 8551
rect 19536 8520 20821 8548
rect 2314 8440 2320 8492
rect 2372 8480 2378 8492
rect 2593 8483 2651 8489
rect 2593 8480 2605 8483
rect 2372 8452 2605 8480
rect 2372 8440 2378 8452
rect 2593 8449 2605 8452
rect 2639 8449 2651 8483
rect 2593 8443 2651 8449
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5537 8483 5595 8489
rect 5537 8480 5549 8483
rect 5500 8452 5549 8480
rect 5500 8440 5506 8452
rect 5537 8449 5549 8452
rect 5583 8480 5595 8483
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5583 8452 6193 8480
rect 5583 8449 5595 8452
rect 5537 8443 5595 8449
rect 6181 8449 6193 8452
rect 6227 8480 6239 8483
rect 6917 8483 6975 8489
rect 6917 8480 6929 8483
rect 6227 8452 6929 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6917 8449 6929 8452
rect 6963 8449 6975 8483
rect 7190 8480 7196 8492
rect 7151 8452 7196 8480
rect 6917 8443 6975 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 8849 8483 8907 8489
rect 8849 8449 8861 8483
rect 8895 8480 8907 8483
rect 9214 8480 9220 8492
rect 8895 8452 9220 8480
rect 8895 8449 8907 8452
rect 8849 8443 8907 8449
rect 9214 8440 9220 8452
rect 9272 8440 9278 8492
rect 10686 8480 10692 8492
rect 10647 8452 10692 8480
rect 10686 8440 10692 8452
rect 10744 8440 10750 8492
rect 12526 8480 12532 8492
rect 12487 8452 12532 8480
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 13872 8452 14565 8480
rect 13872 8440 13878 8452
rect 14553 8449 14565 8452
rect 14599 8480 14611 8483
rect 14642 8480 14648 8492
rect 14599 8452 14648 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17828 8384 18061 8412
rect 17828 8372 17834 8384
rect 18049 8381 18061 8384
rect 18095 8412 18107 8415
rect 18509 8415 18567 8421
rect 18509 8412 18521 8415
rect 18095 8384 18521 8412
rect 18095 8381 18107 8384
rect 18049 8375 18107 8381
rect 18509 8381 18521 8384
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 18782 8372 18788 8424
rect 18840 8412 18846 8424
rect 19061 8415 19119 8421
rect 19061 8412 19073 8415
rect 18840 8384 19073 8412
rect 18840 8372 18846 8384
rect 19061 8381 19073 8384
rect 19107 8381 19119 8415
rect 19061 8375 19119 8381
rect 19242 8372 19248 8424
rect 19300 8412 19306 8424
rect 19536 8421 19564 8520
rect 20809 8517 20821 8520
rect 20855 8517 20867 8551
rect 20809 8511 20867 8517
rect 21174 8508 21180 8560
rect 21232 8548 21238 8560
rect 21542 8548 21548 8560
rect 21232 8520 21548 8548
rect 21232 8508 21238 8520
rect 21542 8508 21548 8520
rect 21600 8508 21606 8560
rect 23014 8508 23020 8560
rect 23072 8548 23078 8560
rect 23072 8520 24256 8548
rect 23072 8508 23078 8520
rect 24228 8492 24256 8520
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 21266 8440 21272 8492
rect 21324 8480 21330 8492
rect 21453 8483 21511 8489
rect 21453 8480 21465 8483
rect 21324 8452 21465 8480
rect 21324 8440 21330 8452
rect 21453 8449 21465 8452
rect 21499 8449 21511 8483
rect 21818 8480 21824 8492
rect 21779 8452 21824 8480
rect 21453 8443 21511 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 23198 8440 23204 8492
rect 23256 8480 23262 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23256 8452 23949 8480
rect 23256 8440 23262 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 24210 8480 24216 8492
rect 24123 8452 24216 8480
rect 23937 8443 23995 8449
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 19521 8415 19579 8421
rect 19521 8412 19533 8415
rect 19300 8384 19533 8412
rect 19300 8372 19306 8384
rect 19521 8381 19533 8384
rect 19567 8381 19579 8415
rect 19521 8375 19579 8381
rect 19889 8415 19947 8421
rect 19889 8381 19901 8415
rect 19935 8381 19947 8415
rect 19889 8375 19947 8381
rect 2314 8344 2320 8356
rect 2275 8316 2320 8344
rect 2314 8304 2320 8316
rect 2372 8304 2378 8356
rect 2409 8347 2467 8353
rect 2409 8313 2421 8347
rect 2455 8344 2467 8347
rect 2682 8344 2688 8356
rect 2455 8316 2688 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4338 8344 4344 8356
rect 3743 8316 4344 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 2700 8276 2728 8304
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 2700 8248 3249 8276
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3237 8239 3295 8245
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 5074 8276 5080 8288
rect 4120 8248 5080 8276
rect 4120 8236 4126 8248
rect 5074 8236 5080 8248
rect 5132 8236 5138 8288
rect 5276 8276 5304 8307
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 7009 8347 7067 8353
rect 5408 8316 5453 8344
rect 5408 8304 5414 8316
rect 7009 8313 7021 8347
rect 7055 8313 7067 8347
rect 7009 8307 7067 8313
rect 9170 8347 9228 8353
rect 9170 8313 9182 8347
rect 9216 8313 9228 8347
rect 9170 8307 9228 8313
rect 10781 8347 10839 8353
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11146 8344 11152 8356
rect 10827 8316 11152 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 5626 8276 5632 8288
rect 5276 8248 5632 8276
rect 5626 8236 5632 8248
rect 5684 8276 5690 8288
rect 6546 8276 6552 8288
rect 5684 8248 6552 8276
rect 5684 8236 5690 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 6822 8276 6828 8288
rect 6687 8248 6828 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 6822 8236 6828 8248
rect 6880 8276 6886 8288
rect 7024 8276 7052 8307
rect 8754 8276 8760 8288
rect 6880 8248 7052 8276
rect 8715 8248 8760 8276
rect 6880 8236 6886 8248
rect 8754 8236 8760 8248
rect 8812 8276 8818 8288
rect 9185 8276 9213 8307
rect 8812 8248 9213 8276
rect 10505 8279 10563 8285
rect 8812 8236 8818 8248
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10796 8276 10824 8307
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11882 8344 11888 8356
rect 11379 8316 11888 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8313 12679 8347
rect 12621 8307 12679 8313
rect 13173 8347 13231 8353
rect 13173 8313 13185 8347
rect 13219 8344 13231 8347
rect 13262 8344 13268 8356
rect 13219 8316 13268 8344
rect 13219 8313 13231 8316
rect 13173 8307 13231 8313
rect 10551 8248 10824 8276
rect 12253 8279 12311 8285
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 12434 8276 12440 8288
rect 12299 8248 12440 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 12434 8236 12440 8248
rect 12492 8276 12498 8288
rect 12636 8276 12664 8307
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 14274 8344 14280 8356
rect 14235 8316 14280 8344
rect 14274 8304 14280 8316
rect 14332 8304 14338 8356
rect 14369 8347 14427 8353
rect 14369 8313 14381 8347
rect 14415 8313 14427 8347
rect 15838 8344 15844 8356
rect 15799 8316 15844 8344
rect 14369 8307 14427 8313
rect 12492 8248 12664 8276
rect 14093 8279 14151 8285
rect 12492 8236 12498 8248
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14384 8276 14412 8307
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 15930 8304 15936 8356
rect 15988 8344 15994 8356
rect 19904 8344 19932 8375
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20036 8384 20269 8412
rect 20036 8372 20042 8384
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 25406 8412 25412 8424
rect 25367 8384 25412 8412
rect 20257 8375 20315 8381
rect 25406 8372 25412 8384
rect 25464 8412 25470 8424
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 25464 8384 25973 8412
rect 25464 8372 25470 8384
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 25961 8375 26019 8381
rect 15988 8316 16033 8344
rect 18892 8316 19932 8344
rect 21545 8347 21603 8353
rect 15988 8304 15994 8316
rect 18892 8288 18920 8316
rect 21545 8313 21557 8347
rect 21591 8313 21603 8347
rect 21545 8307 21603 8313
rect 15378 8276 15384 8288
rect 14139 8248 15384 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 15654 8276 15660 8288
rect 15615 8248 15660 8276
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 18874 8276 18880 8288
rect 18835 8248 18880 8276
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 21174 8276 21180 8288
rect 21135 8248 21180 8276
rect 21174 8236 21180 8248
rect 21232 8276 21238 8288
rect 21560 8276 21588 8307
rect 23014 8304 23020 8356
rect 23072 8344 23078 8356
rect 23750 8344 23756 8356
rect 23072 8316 23756 8344
rect 23072 8304 23078 8316
rect 23750 8304 23756 8316
rect 23808 8344 23814 8356
rect 24029 8347 24087 8353
rect 24029 8344 24041 8347
rect 23808 8316 24041 8344
rect 23808 8304 23814 8316
rect 24029 8313 24041 8316
rect 24075 8313 24087 8347
rect 24029 8307 24087 8313
rect 21232 8248 21588 8276
rect 25317 8279 25375 8285
rect 21232 8236 21238 8248
rect 25317 8245 25329 8279
rect 25363 8276 25375 8279
rect 25774 8276 25780 8288
rect 25363 8248 25780 8276
rect 25363 8245 25375 8248
rect 25317 8239 25375 8245
rect 25774 8236 25780 8248
rect 25832 8236 25838 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1728 8044 1777 8072
rect 1728 8032 1734 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2924 8044 2973 8072
rect 2924 8032 2930 8044
rect 2961 8041 2973 8044
rect 3007 8072 3019 8075
rect 6638 8072 6644 8084
rect 3007 8044 6644 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 6822 8032 6828 8084
rect 6880 8072 6886 8084
rect 6917 8075 6975 8081
rect 6917 8072 6929 8075
rect 6880 8044 6929 8072
rect 6880 8032 6886 8044
rect 6917 8041 6929 8044
rect 6963 8041 6975 8075
rect 6917 8035 6975 8041
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7064 8044 7849 8072
rect 7064 8032 7070 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 11054 8072 11060 8084
rect 11015 8044 11060 8072
rect 7837 8035 7895 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11698 8072 11704 8084
rect 11164 8044 11704 8072
rect 2133 8007 2191 8013
rect 2133 7973 2145 8007
rect 2179 8004 2191 8007
rect 2498 8004 2504 8016
rect 2179 7976 2504 8004
rect 2179 7973 2191 7976
rect 2133 7967 2191 7973
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 3142 7964 3148 8016
rect 3200 8004 3206 8016
rect 3970 8004 3976 8016
rect 3200 7976 3976 8004
rect 3200 7964 3206 7976
rect 3970 7964 3976 7976
rect 4028 8004 4034 8016
rect 4157 8007 4215 8013
rect 4157 8004 4169 8007
rect 4028 7976 4169 8004
rect 4028 7964 4034 7976
rect 4157 7973 4169 7976
rect 4203 7973 4215 8007
rect 4157 7967 4215 7973
rect 4249 8007 4307 8013
rect 4249 7973 4261 8007
rect 4295 8004 4307 8007
rect 4430 8004 4436 8016
rect 4295 7976 4436 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 4430 7964 4436 7976
rect 4488 8004 4494 8016
rect 5350 8004 5356 8016
rect 4488 7976 5356 8004
rect 4488 7964 4494 7976
rect 5350 7964 5356 7976
rect 5408 7964 5414 8016
rect 5626 8004 5632 8016
rect 5587 7976 5632 8004
rect 5626 7964 5632 7976
rect 5684 7964 5690 8016
rect 5994 7964 6000 8016
rect 6052 8004 6058 8016
rect 6359 8007 6417 8013
rect 6359 8004 6371 8007
rect 6052 7976 6371 8004
rect 6052 7964 6058 7976
rect 6359 7973 6371 7976
rect 6405 8004 6417 8007
rect 6454 8004 6460 8016
rect 6405 7976 6460 8004
rect 6405 7973 6417 7976
rect 6359 7967 6417 7973
rect 6454 7964 6460 7976
rect 6512 7964 6518 8016
rect 7282 8004 7288 8016
rect 7243 7976 7288 8004
rect 7282 7964 7288 7976
rect 7340 8004 7346 8016
rect 9858 8004 9864 8016
rect 7340 7976 8248 8004
rect 9819 7976 9864 8004
rect 7340 7964 7346 7976
rect 5074 7896 5080 7948
rect 5132 7936 5138 7948
rect 6012 7936 6040 7964
rect 5132 7908 6040 7936
rect 5132 7896 5138 7908
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7708 7908 7757 7936
rect 7708 7896 7714 7908
rect 7745 7905 7757 7908
rect 7791 7936 7803 7939
rect 7926 7936 7932 7948
rect 7791 7908 7932 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 7926 7896 7932 7908
rect 7984 7896 7990 7948
rect 8220 7945 8248 7976
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 11164 8004 11192 8044
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 14274 8072 14280 8084
rect 14235 8044 14280 8072
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 16114 8072 16120 8084
rect 16075 8044 16120 8072
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16298 8072 16304 8084
rect 16259 8044 16304 8072
rect 16298 8032 16304 8044
rect 16356 8032 16362 8084
rect 17218 8032 17224 8084
rect 17276 8072 17282 8084
rect 17957 8075 18015 8081
rect 17957 8072 17969 8075
rect 17276 8044 17969 8072
rect 17276 8032 17282 8044
rect 17957 8041 17969 8044
rect 18003 8041 18015 8075
rect 19334 8072 19340 8084
rect 17957 8035 18015 8041
rect 18064 8044 19340 8072
rect 10008 7976 11192 8004
rect 11425 8007 11483 8013
rect 10008 7964 10014 7976
rect 11425 7973 11437 8007
rect 11471 8004 11483 8007
rect 11974 8004 11980 8016
rect 11471 7976 11980 8004
rect 11471 7973 11483 7976
rect 11425 7967 11483 7973
rect 11974 7964 11980 7976
rect 12032 7964 12038 8016
rect 12894 8004 12900 8016
rect 12855 7976 12900 8004
rect 12894 7964 12900 7976
rect 12952 7964 12958 8016
rect 12986 7964 12992 8016
rect 13044 8004 13050 8016
rect 18064 8004 18092 8044
rect 19334 8032 19340 8044
rect 19392 8072 19398 8084
rect 19978 8072 19984 8084
rect 19392 8044 19984 8072
rect 19392 8032 19398 8044
rect 19978 8032 19984 8044
rect 20036 8072 20042 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 20036 8044 20269 8072
rect 20036 8032 20042 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 21266 8032 21272 8084
rect 21324 8072 21330 8084
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21324 8044 21925 8072
rect 21324 8032 21330 8044
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 23014 8072 23020 8084
rect 22975 8044 23020 8072
rect 21913 8035 21971 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 23198 8032 23204 8084
rect 23256 8072 23262 8084
rect 23661 8075 23719 8081
rect 23661 8072 23673 8075
rect 23256 8044 23673 8072
rect 23256 8032 23262 8044
rect 23661 8041 23673 8044
rect 23707 8041 23719 8075
rect 24213 8075 24271 8081
rect 24213 8072 24225 8075
rect 23661 8035 23719 8041
rect 23860 8044 24225 8072
rect 13044 7976 13089 8004
rect 17604 7976 18092 8004
rect 18141 8007 18199 8013
rect 13044 7964 13050 7976
rect 8205 7939 8263 7945
rect 8205 7905 8217 7939
rect 8251 7905 8263 7939
rect 8205 7899 8263 7905
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9214 7936 9220 7948
rect 8987 7908 9220 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15712 7908 15761 7936
rect 15712 7896 15718 7908
rect 15749 7905 15761 7908
rect 15795 7936 15807 7939
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 15795 7908 16497 7936
rect 15795 7905 15807 7908
rect 15749 7899 15807 7905
rect 16485 7905 16497 7908
rect 16531 7936 16543 7939
rect 16574 7936 16580 7948
rect 16531 7908 16580 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 16669 7899 16727 7905
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 3786 7868 3792 7880
rect 2087 7840 3792 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4338 7868 4344 7880
rect 4264 7840 4344 7868
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 2593 7803 2651 7809
rect 2593 7800 2605 7803
rect 2372 7772 2605 7800
rect 2372 7760 2378 7772
rect 2593 7769 2605 7772
rect 2639 7800 2651 7803
rect 4264 7800 4292 7840
rect 4338 7828 4344 7840
rect 4396 7868 4402 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4396 7840 4445 7868
rect 4396 7828 4402 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 5994 7868 6000 7880
rect 5955 7840 6000 7868
rect 4433 7831 4491 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7190 7868 7196 7880
rect 6972 7840 7196 7868
rect 6972 7828 6978 7840
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 9769 7871 9827 7877
rect 9769 7837 9781 7871
rect 9815 7837 9827 7871
rect 10042 7868 10048 7880
rect 10003 7840 10048 7868
rect 9769 7831 9827 7837
rect 2639 7772 4292 7800
rect 2639 7769 2651 7772
rect 2593 7763 2651 7769
rect 4890 7760 4896 7812
rect 4948 7800 4954 7812
rect 9401 7803 9459 7809
rect 9401 7800 9413 7803
rect 4948 7772 9413 7800
rect 4948 7760 4954 7772
rect 9401 7769 9413 7772
rect 9447 7800 9459 7803
rect 9784 7800 9812 7831
rect 10042 7828 10048 7840
rect 10100 7868 10106 7880
rect 11333 7871 11391 7877
rect 11333 7868 11345 7871
rect 10100 7840 11345 7868
rect 10100 7828 10106 7840
rect 11333 7837 11345 7840
rect 11379 7868 11391 7871
rect 11698 7868 11704 7880
rect 11379 7840 11704 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 13170 7868 13176 7880
rect 13131 7840 13176 7868
rect 13170 7828 13176 7840
rect 13228 7868 13234 7880
rect 14274 7868 14280 7880
rect 13228 7840 14280 7868
rect 13228 7828 13234 7840
rect 14274 7828 14280 7840
rect 14332 7828 14338 7880
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16684 7868 16712 7899
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 17000 7908 17049 7936
rect 17000 7896 17006 7908
rect 17037 7905 17049 7908
rect 17083 7905 17095 7939
rect 17037 7899 17095 7905
rect 17310 7896 17316 7948
rect 17368 7936 17374 7948
rect 17604 7945 17632 7976
rect 18141 7973 18153 8007
rect 18187 8004 18199 8007
rect 18417 8007 18475 8013
rect 18417 8004 18429 8007
rect 18187 7976 18429 8004
rect 18187 7973 18199 7976
rect 18141 7967 18199 7973
rect 18417 7973 18429 7976
rect 18463 8004 18475 8007
rect 18690 8004 18696 8016
rect 18463 7976 18696 8004
rect 18463 7973 18475 7976
rect 18417 7967 18475 7973
rect 18690 7964 18696 7976
rect 18748 7964 18754 8016
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 22459 8007 22517 8013
rect 18932 7976 19380 8004
rect 18932 7964 18938 7976
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 17368 7908 17601 7936
rect 17368 7896 17374 7908
rect 17589 7905 17601 7908
rect 17635 7905 17647 7939
rect 17589 7899 17647 7905
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 18509 7939 18567 7945
rect 18509 7936 18521 7939
rect 17920 7908 18521 7936
rect 17920 7896 17926 7908
rect 18509 7905 18521 7908
rect 18555 7936 18567 7939
rect 18782 7936 18788 7948
rect 18555 7908 18788 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 19352 7945 19380 7976
rect 22459 7973 22471 8007
rect 22505 8004 22517 8007
rect 22554 8004 22560 8016
rect 22505 7976 22560 8004
rect 22505 7973 22517 7976
rect 22459 7967 22517 7973
rect 22554 7964 22560 7976
rect 22612 8004 22618 8016
rect 23860 8004 23888 8044
rect 24213 8041 24225 8044
rect 24259 8041 24271 8075
rect 24762 8072 24768 8084
rect 24723 8044 24768 8072
rect 24213 8035 24271 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 22612 7976 23888 8004
rect 22612 7964 22618 7976
rect 18969 7939 19027 7945
rect 18969 7905 18981 7939
rect 19015 7905 19027 7939
rect 18969 7899 19027 7905
rect 19337 7939 19395 7945
rect 19337 7905 19349 7939
rect 19383 7905 19395 7939
rect 19337 7899 19395 7905
rect 16448 7840 16712 7868
rect 16448 7828 16454 7840
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18984 7868 19012 7899
rect 19518 7896 19524 7948
rect 19576 7936 19582 7948
rect 19705 7939 19763 7945
rect 19705 7936 19717 7939
rect 19576 7908 19717 7936
rect 19576 7896 19582 7908
rect 19705 7905 19717 7908
rect 19751 7905 19763 7939
rect 19705 7899 19763 7905
rect 20898 7896 20904 7948
rect 20956 7936 20962 7948
rect 21120 7939 21178 7945
rect 21120 7936 21132 7939
rect 20956 7908 21132 7936
rect 20956 7896 20962 7908
rect 21120 7905 21132 7908
rect 21166 7905 21178 7939
rect 21120 7899 21178 7905
rect 21450 7896 21456 7948
rect 21508 7936 21514 7948
rect 21508 7908 23474 7936
rect 21508 7896 21514 7908
rect 19242 7868 19248 7880
rect 17828 7840 19248 7868
rect 17828 7828 17834 7840
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19981 7871 20039 7877
rect 19981 7837 19993 7871
rect 20027 7868 20039 7871
rect 22094 7868 22100 7880
rect 20027 7840 22100 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 23446 7868 23474 7908
rect 23845 7871 23903 7877
rect 23845 7868 23857 7871
rect 23446 7840 23857 7868
rect 23845 7837 23857 7840
rect 23891 7868 23903 7871
rect 24946 7868 24952 7880
rect 23891 7840 24952 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 24946 7828 24952 7840
rect 25004 7828 25010 7880
rect 11882 7800 11888 7812
rect 9447 7772 9812 7800
rect 11795 7772 11888 7800
rect 9447 7769 9459 7772
rect 9401 7763 9459 7769
rect 11882 7760 11888 7772
rect 11940 7800 11946 7812
rect 13078 7800 13084 7812
rect 11940 7772 13084 7800
rect 11940 7760 11946 7772
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 21223 7803 21281 7809
rect 21223 7800 21235 7803
rect 15896 7772 21235 7800
rect 15896 7760 15902 7772
rect 21223 7769 21235 7772
rect 21269 7769 21281 7803
rect 21223 7763 21281 7769
rect 5166 7732 5172 7744
rect 5127 7704 5172 7732
rect 5166 7692 5172 7704
rect 5224 7732 5230 7744
rect 5350 7732 5356 7744
rect 5224 7704 5356 7732
rect 5224 7692 5230 7704
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 7098 7692 7104 7744
rect 7156 7732 7162 7744
rect 12250 7732 12256 7744
rect 7156 7704 12256 7732
rect 7156 7692 7162 7704
rect 12250 7692 12256 7704
rect 12308 7692 12314 7744
rect 12710 7732 12716 7744
rect 12671 7704 12716 7732
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15562 7732 15568 7744
rect 15151 7704 15568 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 18141 7735 18199 7741
rect 18141 7732 18153 7735
rect 15712 7704 18153 7732
rect 15712 7692 15718 7704
rect 18141 7701 18153 7704
rect 18187 7701 18199 7735
rect 20714 7732 20720 7744
rect 20675 7704 20720 7732
rect 18141 7695 18199 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21545 7735 21603 7741
rect 21545 7732 21557 7735
rect 21416 7704 21557 7732
rect 21416 7692 21422 7704
rect 21545 7701 21557 7704
rect 21591 7701 21603 7735
rect 21545 7695 21603 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2777 7531 2835 7537
rect 2777 7528 2789 7531
rect 2648 7500 2789 7528
rect 2648 7488 2654 7500
rect 2777 7497 2789 7500
rect 2823 7497 2835 7531
rect 2777 7491 2835 7497
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3786 7528 3792 7540
rect 3191 7500 3792 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 5169 7531 5227 7537
rect 5169 7528 5181 7531
rect 4028 7500 5181 7528
rect 4028 7488 4034 7500
rect 5169 7497 5181 7500
rect 5215 7497 5227 7531
rect 5169 7491 5227 7497
rect 5859 7531 5917 7537
rect 5859 7497 5871 7531
rect 5905 7528 5917 7531
rect 8846 7528 8852 7540
rect 5905 7500 8852 7528
rect 5905 7497 5917 7500
rect 5859 7491 5917 7497
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9030 7528 9036 7540
rect 8991 7500 9036 7528
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9858 7488 9864 7540
rect 9916 7528 9922 7540
rect 10137 7531 10195 7537
rect 10137 7528 10149 7531
rect 9916 7500 10149 7528
rect 9916 7488 9922 7500
rect 10137 7497 10149 7500
rect 10183 7497 10195 7531
rect 10137 7491 10195 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 11974 7528 11980 7540
rect 11931 7500 11980 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 14553 7531 14611 7537
rect 14553 7528 14565 7531
rect 13596 7500 14565 7528
rect 13596 7488 13602 7500
rect 14553 7497 14565 7500
rect 14599 7497 14611 7531
rect 14553 7491 14611 7497
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 14792 7500 14841 7528
rect 14792 7488 14798 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 16390 7528 16396 7540
rect 14829 7491 14887 7497
rect 15304 7500 16396 7528
rect 3620 7432 6960 7460
rect 3620 7404 3648 7432
rect 1670 7352 1676 7404
rect 1728 7392 1734 7404
rect 1857 7395 1915 7401
rect 1857 7392 1869 7395
rect 1728 7364 1869 7392
rect 1728 7352 1734 7364
rect 1857 7361 1869 7364
rect 1903 7361 1915 7395
rect 3602 7392 3608 7404
rect 3515 7364 3608 7392
rect 1857 7355 1915 7361
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 4522 7352 4528 7404
rect 4580 7392 4586 7404
rect 5902 7392 5908 7404
rect 4580 7364 5908 7392
rect 4580 7352 4586 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 6932 7392 6960 7432
rect 9122 7420 9128 7472
rect 9180 7460 9186 7472
rect 9766 7460 9772 7472
rect 9180 7432 9260 7460
rect 9727 7432 9772 7460
rect 9180 7420 9186 7432
rect 9232 7401 9260 7432
rect 9766 7420 9772 7432
rect 9824 7420 9830 7472
rect 11514 7420 11520 7472
rect 11572 7460 11578 7472
rect 12161 7463 12219 7469
rect 12161 7460 12173 7463
rect 11572 7432 12173 7460
rect 11572 7420 11578 7432
rect 12161 7429 12173 7432
rect 12207 7429 12219 7463
rect 12161 7423 12219 7429
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 15304 7460 15332 7500
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17405 7531 17463 7537
rect 17405 7528 17417 7531
rect 16632 7500 17417 7528
rect 16632 7488 16638 7500
rect 17405 7497 17417 7500
rect 17451 7497 17463 7531
rect 17405 7491 17463 7497
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 21140 7500 21189 7528
rect 21140 7488 21146 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 22370 7488 22376 7540
rect 22428 7528 22434 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22428 7500 23029 7528
rect 22428 7488 22434 7500
rect 23017 7497 23029 7500
rect 23063 7528 23075 7531
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 23063 7500 23213 7528
rect 23063 7497 23075 7500
rect 23017 7491 23075 7497
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 24946 7528 24952 7540
rect 24907 7500 24952 7528
rect 23201 7491 23259 7497
rect 24946 7488 24952 7500
rect 25004 7488 25010 7540
rect 14323 7432 15332 7460
rect 15565 7463 15623 7469
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 15565 7429 15577 7463
rect 15611 7460 15623 7463
rect 16942 7460 16948 7472
rect 15611 7432 16948 7460
rect 15611 7429 15623 7432
rect 15565 7423 15623 7429
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 6932 7364 7389 7392
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7361 9275 7395
rect 12176 7392 12204 7423
rect 16942 7420 16948 7432
rect 17000 7460 17006 7472
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 17000 7432 18245 7460
rect 17000 7420 17006 7432
rect 18233 7429 18245 7432
rect 18279 7460 18291 7463
rect 18874 7460 18880 7472
rect 18279 7432 18880 7460
rect 18279 7429 18291 7432
rect 18233 7423 18291 7429
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 22554 7460 22560 7472
rect 22515 7432 22560 7460
rect 22554 7420 22560 7432
rect 22612 7420 22618 7472
rect 22830 7420 22836 7472
rect 22888 7460 22894 7472
rect 22888 7432 25544 7460
rect 22888 7420 22894 7432
rect 12176 7364 12572 7392
rect 9217 7355 9275 7361
rect 4798 7284 4804 7336
rect 4856 7324 4862 7336
rect 5756 7327 5814 7333
rect 5756 7324 5768 7327
rect 4856 7296 5768 7324
rect 4856 7284 4862 7296
rect 5756 7293 5768 7296
rect 5802 7324 5814 7327
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 5802 7296 6193 7324
rect 5802 7293 5814 7296
rect 5756 7287 5814 7293
rect 6181 7293 6193 7296
rect 6227 7324 6239 7327
rect 6270 7324 6276 7336
rect 6227 7296 6276 7324
rect 6227 7293 6239 7296
rect 6181 7287 6239 7293
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 6748 7324 6776 7352
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6748 7296 6929 7324
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 6917 7287 6975 7293
rect 1765 7259 1823 7265
rect 1765 7225 1777 7259
rect 1811 7256 1823 7259
rect 1854 7256 1860 7268
rect 1811 7228 1860 7256
rect 1811 7225 1823 7228
rect 1765 7219 1823 7225
rect 1854 7216 1860 7228
rect 1912 7256 1918 7268
rect 2219 7259 2277 7265
rect 2219 7256 2231 7259
rect 1912 7228 2231 7256
rect 1912 7216 1918 7228
rect 2219 7225 2231 7228
rect 2265 7256 2277 7259
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 2265 7228 3525 7256
rect 2265 7225 2277 7228
rect 2219 7219 2277 7225
rect 3513 7225 3525 7228
rect 3559 7256 3571 7259
rect 3967 7259 4025 7265
rect 3967 7256 3979 7259
rect 3559 7228 3979 7256
rect 3559 7225 3571 7228
rect 3513 7219 3571 7225
rect 3967 7225 3979 7228
rect 4013 7256 4025 7259
rect 4062 7256 4068 7268
rect 4013 7228 4068 7256
rect 4013 7225 4025 7228
rect 3967 7219 4025 7225
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5166 7256 5172 7268
rect 4939 7228 5172 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5166 7216 5172 7228
rect 5224 7256 5230 7268
rect 6730 7256 6736 7268
rect 5224 7228 6736 7256
rect 5224 7216 5230 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 6822 7216 6828 7268
rect 6880 7256 6886 7268
rect 6932 7256 6960 7287
rect 7282 7284 7288 7296
rect 7340 7324 7346 7336
rect 8110 7324 8116 7336
rect 7340 7296 8116 7324
rect 7340 7284 7346 7296
rect 8110 7284 8116 7296
rect 8168 7324 8174 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 8168 7296 8217 7324
rect 8168 7284 8174 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 10689 7327 10747 7333
rect 10689 7293 10701 7327
rect 10735 7324 10747 7327
rect 11425 7327 11483 7333
rect 11425 7324 11437 7327
rect 10735 7296 11437 7324
rect 10735 7293 10747 7296
rect 10689 7287 10747 7293
rect 11425 7293 11437 7296
rect 11471 7324 11483 7327
rect 11471 7296 12480 7324
rect 11471 7293 11483 7296
rect 11425 7287 11483 7293
rect 8754 7256 8760 7268
rect 6880 7228 6960 7256
rect 7024 7228 8760 7256
rect 6880 7216 6886 7228
rect 2130 7148 2136 7200
rect 2188 7188 2194 7200
rect 3142 7188 3148 7200
rect 2188 7160 3148 7188
rect 2188 7148 2194 7160
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6512 7160 6653 7188
rect 6512 7148 6518 7160
rect 6641 7157 6653 7160
rect 6687 7188 6699 7191
rect 7024 7188 7052 7228
rect 8754 7216 8760 7228
rect 8812 7216 8818 7268
rect 9030 7216 9036 7268
rect 9088 7256 9094 7268
rect 9309 7259 9367 7265
rect 9309 7256 9321 7259
rect 9088 7228 9321 7256
rect 9088 7216 9094 7228
rect 9309 7225 9321 7228
rect 9355 7225 9367 7259
rect 11514 7256 11520 7268
rect 11475 7228 11520 7256
rect 9309 7219 9367 7225
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 12452 7200 12480 7296
rect 12544 7256 12572 7364
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 13817 7395 13875 7401
rect 13817 7392 13829 7395
rect 13044 7364 13829 7392
rect 13044 7352 13050 7364
rect 13817 7361 13829 7364
rect 13863 7361 13875 7395
rect 16574 7392 16580 7404
rect 13817 7355 13875 7361
rect 15948 7364 16580 7392
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7324 12679 7327
rect 12710 7324 12716 7336
rect 12667 7296 12716 7324
rect 12667 7293 12679 7296
rect 12621 7287 12679 7293
rect 12710 7284 12716 7296
rect 12768 7324 12774 7336
rect 14369 7327 14427 7333
rect 12768 7296 13814 7324
rect 12768 7284 12774 7296
rect 12942 7259 13000 7265
rect 12942 7256 12954 7259
rect 12544 7228 12954 7256
rect 12942 7225 12954 7228
rect 12988 7225 13000 7259
rect 13786 7256 13814 7296
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14734 7324 14740 7336
rect 14415 7296 14740 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 15948 7333 15976 7364
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 18598 7352 18604 7404
rect 18656 7392 18662 7404
rect 20533 7395 20591 7401
rect 18656 7364 19932 7392
rect 18656 7352 18662 7364
rect 15933 7327 15991 7333
rect 15933 7293 15945 7327
rect 15979 7293 15991 7327
rect 15933 7287 15991 7293
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7293 16175 7327
rect 16117 7287 16175 7293
rect 16132 7256 16160 7287
rect 16206 7284 16212 7336
rect 16264 7324 16270 7336
rect 16485 7327 16543 7333
rect 16485 7324 16497 7327
rect 16264 7296 16497 7324
rect 16264 7284 16270 7296
rect 16485 7293 16497 7296
rect 16531 7293 16543 7327
rect 16485 7287 16543 7293
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17037 7327 17095 7333
rect 17037 7324 17049 7327
rect 17000 7296 17049 7324
rect 17000 7284 17006 7296
rect 17037 7293 17049 7296
rect 17083 7324 17095 7327
rect 17310 7324 17316 7336
rect 17083 7296 17316 7324
rect 17083 7293 17095 7296
rect 17037 7287 17095 7293
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7324 18110 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18104 7296 18521 7324
rect 18104 7284 18110 7296
rect 18509 7293 18521 7296
rect 18555 7293 18567 7327
rect 18509 7287 18567 7293
rect 18782 7284 18788 7336
rect 18840 7324 18846 7336
rect 19058 7324 19064 7336
rect 18840 7296 19064 7324
rect 18840 7284 18846 7296
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19904 7333 19932 7364
rect 20533 7361 20545 7395
rect 20579 7392 20591 7395
rect 21450 7392 21456 7404
rect 20579 7364 21456 7392
rect 20579 7361 20591 7364
rect 20533 7355 20591 7361
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 19521 7327 19579 7333
rect 19521 7324 19533 7327
rect 19300 7296 19533 7324
rect 19300 7284 19306 7296
rect 19521 7293 19533 7296
rect 19567 7293 19579 7327
rect 19521 7287 19579 7293
rect 19889 7327 19947 7333
rect 19889 7293 19901 7327
rect 19935 7324 19947 7327
rect 19978 7324 19984 7336
rect 19935 7296 19984 7324
rect 19935 7293 19947 7296
rect 19889 7287 19947 7293
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20257 7327 20315 7333
rect 20257 7293 20269 7327
rect 20303 7293 20315 7327
rect 20257 7287 20315 7293
rect 16666 7256 16672 7268
rect 13786 7228 15608 7256
rect 16132 7228 16672 7256
rect 12942 7219 13000 7225
rect 6687 7160 7052 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 7837 7191 7895 7197
rect 7837 7188 7849 7191
rect 7708 7160 7849 7188
rect 7708 7148 7714 7160
rect 7837 7157 7849 7160
rect 7883 7157 7895 7191
rect 7837 7151 7895 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 13541 7191 13599 7197
rect 13541 7188 13553 7191
rect 12492 7160 13553 7188
rect 12492 7148 12498 7160
rect 13541 7157 13553 7160
rect 13587 7157 13599 7191
rect 15580 7188 15608 7228
rect 16666 7216 16672 7228
rect 16724 7256 16730 7268
rect 17770 7256 17776 7268
rect 16724 7228 17776 7256
rect 16724 7216 16730 7228
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 20272 7256 20300 7287
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 21361 7327 21419 7333
rect 21361 7324 21373 7327
rect 21324 7296 21373 7324
rect 21324 7284 21330 7296
rect 21361 7293 21373 7296
rect 21407 7293 21419 7327
rect 22572 7324 22600 7420
rect 23201 7395 23259 7401
rect 23201 7361 23213 7395
rect 23247 7392 23259 7395
rect 24029 7395 24087 7401
rect 24029 7392 24041 7395
rect 23247 7364 24041 7392
rect 23247 7361 23259 7364
rect 23201 7355 23259 7361
rect 24029 7361 24041 7364
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 24210 7352 24216 7404
rect 24268 7392 24274 7404
rect 24305 7395 24363 7401
rect 24305 7392 24317 7395
rect 24268 7364 24317 7392
rect 24268 7352 24274 7364
rect 24305 7361 24317 7364
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 25516 7333 25544 7432
rect 23385 7327 23443 7333
rect 23385 7324 23397 7327
rect 22572 7296 23397 7324
rect 21361 7287 21419 7293
rect 23385 7293 23397 7296
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 25501 7327 25559 7333
rect 25501 7293 25513 7327
rect 25547 7324 25559 7327
rect 26053 7327 26111 7333
rect 26053 7324 26065 7327
rect 25547 7296 26065 7324
rect 25547 7293 25559 7296
rect 25501 7287 25559 7293
rect 26053 7293 26065 7296
rect 26099 7293 26111 7327
rect 26053 7287 26111 7293
rect 19484 7228 20300 7256
rect 19484 7216 19490 7228
rect 21082 7216 21088 7268
rect 21140 7256 21146 7268
rect 21682 7259 21740 7265
rect 21682 7256 21694 7259
rect 21140 7228 21694 7256
rect 21140 7216 21146 7228
rect 21682 7225 21694 7228
rect 21728 7225 21740 7259
rect 24118 7256 24124 7268
rect 24079 7228 24124 7256
rect 21682 7219 21740 7225
rect 24118 7216 24124 7228
rect 24176 7216 24182 7268
rect 15749 7191 15807 7197
rect 15749 7188 15761 7191
rect 15580 7160 15761 7188
rect 13541 7151 13599 7157
rect 15749 7157 15761 7160
rect 15795 7157 15807 7191
rect 20898 7188 20904 7200
rect 20859 7160 20904 7188
rect 15749 7151 15807 7157
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 21358 7148 21364 7200
rect 21416 7188 21422 7200
rect 22281 7191 22339 7197
rect 22281 7188 22293 7191
rect 21416 7160 22293 7188
rect 21416 7148 21422 7160
rect 22281 7157 22293 7160
rect 22327 7157 22339 7191
rect 25682 7188 25688 7200
rect 25643 7160 25688 7188
rect 22281 7151 22339 7157
rect 25682 7148 25688 7160
rect 25740 7148 25746 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1857 6987 1915 6993
rect 1857 6984 1869 6987
rect 1728 6956 1869 6984
rect 1728 6944 1734 6956
rect 1857 6953 1869 6956
rect 1903 6984 1915 6987
rect 2590 6984 2596 6996
rect 1903 6956 2596 6984
rect 1903 6953 1915 6956
rect 1857 6947 1915 6953
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 3602 6984 3608 6996
rect 3563 6956 3608 6984
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 5994 6984 6000 6996
rect 5684 6956 6000 6984
rect 5684 6944 5690 6956
rect 5994 6944 6000 6956
rect 6052 6984 6058 6996
rect 7653 6987 7711 6993
rect 7653 6984 7665 6987
rect 6052 6956 7665 6984
rect 6052 6944 6058 6956
rect 7653 6953 7665 6956
rect 7699 6953 7711 6987
rect 9122 6984 9128 6996
rect 9083 6956 9128 6984
rect 7653 6947 7711 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 11698 6984 11704 6996
rect 11659 6956 11704 6984
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 13357 6987 13415 6993
rect 13357 6984 13369 6987
rect 12952 6956 13369 6984
rect 12952 6944 12958 6956
rect 13357 6953 13369 6956
rect 13403 6953 13415 6987
rect 13357 6947 13415 6953
rect 14369 6987 14427 6993
rect 14369 6953 14381 6987
rect 14415 6953 14427 6987
rect 14369 6947 14427 6953
rect 2038 6876 2044 6928
rect 2096 6916 2102 6928
rect 2133 6919 2191 6925
rect 2133 6916 2145 6919
rect 2096 6888 2145 6916
rect 2096 6876 2102 6888
rect 2133 6885 2145 6888
rect 2179 6916 2191 6919
rect 4249 6919 4307 6925
rect 4249 6916 4261 6919
rect 2179 6888 4261 6916
rect 2179 6885 2191 6888
rect 2133 6879 2191 6885
rect 4249 6885 4261 6888
rect 4295 6916 4307 6919
rect 4522 6916 4528 6928
rect 4295 6888 4528 6916
rect 4295 6885 4307 6888
rect 4249 6879 4307 6885
rect 4522 6876 4528 6888
rect 4580 6916 4586 6928
rect 4890 6916 4896 6928
rect 4580 6888 4896 6916
rect 4580 6876 4586 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 6175 6919 6233 6925
rect 6175 6885 6187 6919
rect 6221 6916 6233 6919
rect 6454 6916 6460 6928
rect 6221 6888 6460 6916
rect 6221 6885 6233 6888
rect 6175 6879 6233 6885
rect 6454 6876 6460 6888
rect 6512 6876 6518 6928
rect 9858 6916 9864 6928
rect 9819 6888 9864 6916
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 12434 6876 12440 6928
rect 12492 6916 12498 6928
rect 12529 6919 12587 6925
rect 12529 6916 12541 6919
rect 12492 6888 12541 6916
rect 12492 6876 12498 6888
rect 12529 6885 12541 6888
rect 12575 6885 12587 6919
rect 12529 6879 12587 6885
rect 13081 6919 13139 6925
rect 13081 6885 13093 6919
rect 13127 6916 13139 6919
rect 13170 6916 13176 6928
rect 13127 6888 13176 6916
rect 13127 6885 13139 6888
rect 13081 6879 13139 6885
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 14384 6916 14412 6947
rect 14550 6944 14556 6996
rect 14608 6984 14614 6996
rect 16393 6987 16451 6993
rect 16393 6984 16405 6987
rect 14608 6956 16405 6984
rect 14608 6944 14614 6956
rect 16393 6953 16405 6956
rect 16439 6953 16451 6987
rect 16393 6947 16451 6953
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 18782 6984 18788 6996
rect 18380 6956 18788 6984
rect 18380 6944 18386 6956
rect 18782 6944 18788 6956
rect 18840 6984 18846 6996
rect 19061 6987 19119 6993
rect 19061 6984 19073 6987
rect 18840 6956 19073 6984
rect 18840 6944 18846 6956
rect 19061 6953 19073 6956
rect 19107 6984 19119 6987
rect 19426 6984 19432 6996
rect 19107 6956 19432 6984
rect 19107 6953 19119 6956
rect 19061 6947 19119 6953
rect 19426 6944 19432 6956
rect 19484 6944 19490 6996
rect 21082 6984 21088 6996
rect 19904 6956 21088 6984
rect 15654 6916 15660 6928
rect 14384 6888 15660 6916
rect 15654 6876 15660 6888
rect 15712 6876 15718 6928
rect 16206 6876 16212 6928
rect 16264 6916 16270 6928
rect 17310 6916 17316 6928
rect 16264 6888 17316 6916
rect 16264 6876 16270 6888
rect 5534 6808 5540 6860
rect 5592 6848 5598 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5592 6820 5825 6848
rect 5592 6808 5598 6820
rect 5813 6817 5825 6820
rect 5859 6848 5871 6851
rect 7006 6848 7012 6860
rect 5859 6820 7012 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 14185 6851 14243 6857
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 14458 6848 14464 6860
rect 14231 6820 14464 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15838 6848 15844 6860
rect 15335 6820 15844 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15838 6808 15844 6820
rect 15896 6808 15902 6860
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 17144 6857 17172 6888
rect 17310 6876 17316 6888
rect 17368 6876 17374 6928
rect 18598 6876 18604 6928
rect 18656 6916 18662 6928
rect 18693 6919 18751 6925
rect 18693 6916 18705 6919
rect 18656 6888 18705 6916
rect 18656 6876 18662 6888
rect 18693 6885 18705 6888
rect 18739 6885 18751 6919
rect 18693 6879 18751 6885
rect 16761 6851 16819 6857
rect 16761 6848 16773 6851
rect 16724 6820 16773 6848
rect 16724 6808 16730 6820
rect 16761 6817 16773 6820
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 17497 6851 17555 6857
rect 17497 6848 17509 6851
rect 17276 6820 17509 6848
rect 17276 6808 17282 6820
rect 17497 6817 17509 6820
rect 17543 6817 17555 6851
rect 17497 6811 17555 6817
rect 17770 6808 17776 6860
rect 17828 6848 17834 6860
rect 19904 6857 19932 6956
rect 21082 6944 21088 6956
rect 21140 6984 21146 6996
rect 22094 6984 22100 6996
rect 21140 6956 21312 6984
rect 22055 6956 22100 6984
rect 21140 6944 21146 6956
rect 19981 6919 20039 6925
rect 19981 6885 19993 6919
rect 20027 6916 20039 6919
rect 21174 6916 21180 6928
rect 20027 6888 21180 6916
rect 20027 6885 20039 6888
rect 19981 6879 20039 6885
rect 21174 6876 21180 6888
rect 21232 6876 21238 6928
rect 21284 6925 21312 6956
rect 22094 6944 22100 6956
rect 22152 6944 22158 6996
rect 24029 6987 24087 6993
rect 24029 6953 24041 6987
rect 24075 6984 24087 6987
rect 24118 6984 24124 6996
rect 24075 6956 24124 6984
rect 24075 6953 24087 6956
rect 24029 6947 24087 6953
rect 24118 6944 24124 6956
rect 24176 6944 24182 6996
rect 25038 6984 25044 6996
rect 24320 6956 25044 6984
rect 21269 6919 21327 6925
rect 21269 6885 21281 6919
rect 21315 6916 21327 6919
rect 21358 6916 21364 6928
rect 21315 6888 21364 6916
rect 21315 6885 21327 6888
rect 21269 6879 21327 6885
rect 21358 6876 21364 6888
rect 21416 6876 21422 6928
rect 21818 6916 21824 6928
rect 21779 6888 21824 6916
rect 21818 6876 21824 6888
rect 21876 6876 21882 6928
rect 24320 6925 24348 6956
rect 25038 6944 25044 6956
rect 25096 6944 25102 6996
rect 24305 6919 24363 6925
rect 24305 6885 24317 6919
rect 24351 6885 24363 6919
rect 24305 6879 24363 6885
rect 24397 6919 24455 6925
rect 24397 6885 24409 6919
rect 24443 6916 24455 6919
rect 24670 6916 24676 6928
rect 24443 6888 24676 6916
rect 24443 6885 24455 6888
rect 24397 6879 24455 6885
rect 24670 6876 24676 6888
rect 24728 6876 24734 6928
rect 18325 6851 18383 6857
rect 18325 6848 18337 6851
rect 17828 6820 18337 6848
rect 17828 6808 17834 6820
rect 18325 6817 18337 6820
rect 18371 6817 18383 6851
rect 18325 6811 18383 6817
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6817 19947 6851
rect 22738 6848 22744 6860
rect 22699 6820 22744 6848
rect 19889 6811 19947 6817
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 2130 6780 2136 6792
rect 2087 6752 2136 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 4146 6783 4204 6789
rect 4146 6749 4158 6783
rect 4192 6780 4204 6783
rect 4614 6780 4620 6792
rect 4192 6752 4620 6780
rect 4192 6749 4204 6752
rect 4146 6743 4204 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10042 6780 10048 6792
rect 10003 6752 10048 6780
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 10744 6752 11253 6780
rect 10744 6740 10750 6752
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11330 6740 11336 6792
rect 11388 6780 11394 6792
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 11388 6752 12449 6780
rect 11388 6740 11394 6752
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6780 15807 6783
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 15795 6752 16221 6780
rect 15795 6749 15807 6752
rect 15749 6743 15807 6749
rect 16209 6749 16221 6752
rect 16255 6780 16267 6783
rect 16684 6780 16712 6808
rect 16255 6752 16712 6780
rect 21177 6783 21235 6789
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 21177 6749 21189 6783
rect 21223 6780 21235 6783
rect 21542 6780 21548 6792
rect 21223 6752 21548 6780
rect 21223 6749 21235 6752
rect 21177 6743 21235 6749
rect 21542 6740 21548 6752
rect 21600 6780 21606 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 21600 6752 22477 6780
rect 21600 6740 21606 6752
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 23382 6780 23388 6792
rect 23343 6752 23388 6780
rect 22465 6743 22523 6749
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 24762 6780 24768 6792
rect 24723 6752 24768 6780
rect 24762 6740 24768 6752
rect 24820 6740 24826 6792
rect 1210 6672 1216 6724
rect 1268 6712 1274 6724
rect 2498 6712 2504 6724
rect 1268 6684 2504 6712
rect 1268 6672 1274 6684
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2556 6684 2973 6712
rect 2556 6672 2562 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 3108 6684 4721 6712
rect 3108 6672 3114 6684
rect 4709 6681 4721 6684
rect 4755 6712 4767 6715
rect 5442 6712 5448 6724
rect 4755 6684 5448 6712
rect 4755 6681 4767 6684
rect 4709 6675 4767 6681
rect 5442 6672 5448 6684
rect 5500 6672 5506 6724
rect 6730 6712 6736 6724
rect 6691 6684 6736 6712
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 15105 6715 15163 6721
rect 15105 6681 15117 6715
rect 15151 6712 15163 6715
rect 15562 6712 15568 6724
rect 15151 6684 15568 6712
rect 15151 6681 15163 6684
rect 15105 6675 15163 6681
rect 15562 6672 15568 6684
rect 15620 6712 15626 6724
rect 16942 6712 16948 6724
rect 15620 6684 16948 6712
rect 15620 6672 15626 6684
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 845 6647 903 6653
rect 845 6613 857 6647
rect 891 6644 903 6647
rect 3970 6644 3976 6656
rect 891 6616 3976 6644
rect 891 6613 903 6616
rect 845 6607 903 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 6178 6644 6184 6656
rect 4396 6616 6184 6644
rect 4396 6604 4402 6616
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7009 6647 7067 6653
rect 7009 6644 7021 6647
rect 6880 6616 7021 6644
rect 6880 6604 6886 6616
rect 7009 6613 7021 6616
rect 7055 6613 7067 6647
rect 10778 6644 10784 6656
rect 10739 6616 10784 6644
rect 7009 6607 7067 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 16298 6644 16304 6656
rect 15519 6616 16304 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 20254 6644 20260 6656
rect 20215 6616 20260 6644
rect 20254 6604 20260 6616
rect 20312 6644 20318 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20312 6616 20637 6644
rect 20312 6604 20318 6616
rect 20625 6613 20637 6616
rect 20671 6644 20683 6647
rect 20714 6644 20720 6656
rect 20671 6616 20720 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3292 6412 3341 6440
rect 3292 6400 3298 6412
rect 3329 6409 3341 6412
rect 3375 6440 3387 6443
rect 4890 6440 4896 6452
rect 3375 6412 4016 6440
rect 4851 6412 4896 6440
rect 3375 6409 3387 6412
rect 3329 6403 3387 6409
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2498 6304 2504 6316
rect 2455 6276 2504 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 3050 6304 3056 6316
rect 3011 6276 3056 6304
rect 3050 6264 3056 6276
rect 3108 6264 3114 6316
rect 3988 6313 4016 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5534 6440 5540 6452
rect 5495 6412 5540 6440
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6086 6440 6092 6452
rect 5951 6412 6092 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6454 6440 6460 6452
rect 6319 6412 6460 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 8168 6412 8217 6440
rect 8168 6400 8174 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8205 6403 8263 6409
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6440 9827 6443
rect 9858 6440 9864 6452
rect 9815 6412 9864 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 9858 6400 9864 6412
rect 9916 6440 9922 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9916 6412 10057 6440
rect 9916 6400 9922 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10045 6403 10103 6409
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 12621 6443 12679 6449
rect 12621 6440 12633 6443
rect 11572 6412 12633 6440
rect 11572 6400 11578 6412
rect 12621 6409 12633 6412
rect 12667 6440 12679 6443
rect 12986 6440 12992 6452
rect 12667 6412 12992 6440
rect 12667 6409 12679 6412
rect 12621 6403 12679 6409
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 14093 6443 14151 6449
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 14458 6440 14464 6452
rect 14139 6412 14464 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15473 6443 15531 6449
rect 15473 6440 15485 6443
rect 15436 6412 15485 6440
rect 15436 6400 15442 6412
rect 15473 6409 15485 6412
rect 15519 6409 15531 6443
rect 15473 6403 15531 6409
rect 16574 6400 16580 6452
rect 16632 6440 16638 6452
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 16632 6412 17325 6440
rect 16632 6400 16638 6412
rect 17313 6409 17325 6412
rect 17359 6409 17371 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17313 6403 17371 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 18414 6400 18420 6452
rect 18472 6440 18478 6452
rect 18877 6443 18935 6449
rect 18877 6440 18889 6443
rect 18472 6412 18889 6440
rect 18472 6400 18478 6412
rect 18877 6409 18889 6412
rect 18923 6409 18935 6443
rect 18877 6403 18935 6409
rect 6104 6372 6132 6400
rect 11054 6372 11060 6384
rect 6104 6344 9904 6372
rect 9876 6316 9904 6344
rect 10336 6344 11060 6372
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4120 6276 4261 6304
rect 4120 6264 4126 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 9122 6304 9128 6316
rect 8895 6276 9128 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9122 6264 9128 6276
rect 9180 6304 9186 6316
rect 9490 6304 9496 6316
rect 9180 6276 9496 6304
rect 9180 6264 9186 6276
rect 9490 6264 9496 6276
rect 9548 6264 9554 6316
rect 9858 6264 9864 6316
rect 9916 6264 9922 6316
rect 5721 6239 5779 6245
rect 5721 6205 5733 6239
rect 5767 6236 5779 6239
rect 6822 6236 6828 6248
rect 5767 6208 6684 6236
rect 6783 6208 6828 6236
rect 5767 6205 5779 6208
rect 5721 6199 5779 6205
rect 2501 6171 2559 6177
rect 2501 6137 2513 6171
rect 2547 6168 2559 6171
rect 2590 6168 2596 6180
rect 2547 6140 2596 6168
rect 2547 6137 2559 6140
rect 2501 6131 2559 6137
rect 2590 6128 2596 6140
rect 2648 6128 2654 6180
rect 4065 6171 4123 6177
rect 4065 6137 4077 6171
rect 4111 6137 4123 6171
rect 4065 6131 4123 6137
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 3697 6103 3755 6109
rect 3697 6100 3709 6103
rect 3476 6072 3709 6100
rect 3476 6060 3482 6072
rect 3697 6069 3709 6072
rect 3743 6100 3755 6103
rect 4080 6100 4108 6131
rect 6656 6112 6684 6208
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7285 6239 7343 6245
rect 7285 6236 7297 6239
rect 7248 6208 7297 6236
rect 7248 6196 7254 6208
rect 7285 6205 7297 6208
rect 7331 6205 7343 6239
rect 7285 6199 7343 6205
rect 8754 6168 8760 6180
rect 8667 6140 8760 6168
rect 8754 6128 8760 6140
rect 8812 6168 8818 6180
rect 9211 6171 9269 6177
rect 9211 6168 9223 6171
rect 8812 6140 9223 6168
rect 8812 6128 8818 6140
rect 9211 6137 9223 6140
rect 9257 6168 9269 6171
rect 10336 6168 10364 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 11296 6344 11805 6372
rect 11296 6332 11302 6344
rect 11793 6341 11805 6344
rect 11839 6341 11851 6375
rect 11793 6335 11851 6341
rect 16209 6375 16267 6381
rect 16209 6341 16221 6375
rect 16255 6372 16267 6375
rect 16298 6372 16304 6384
rect 16255 6344 16304 6372
rect 16255 6341 16267 6344
rect 16209 6335 16267 6341
rect 16298 6332 16304 6344
rect 16356 6372 16362 6384
rect 18598 6372 18604 6384
rect 16356 6344 18604 6372
rect 16356 6332 16362 6344
rect 18598 6332 18604 6344
rect 18656 6332 18662 6384
rect 18892 6316 18920 6403
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 20036 6412 20821 6440
rect 20036 6400 20042 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 22738 6440 22744 6452
rect 22699 6412 22744 6440
rect 20809 6403 20867 6409
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 25038 6400 25044 6452
rect 25096 6440 25102 6452
rect 25133 6443 25191 6449
rect 25133 6440 25145 6443
rect 25096 6412 25145 6440
rect 25096 6400 25102 6412
rect 25133 6409 25145 6412
rect 25179 6409 25191 6443
rect 25133 6403 25191 6409
rect 24946 6332 24952 6384
rect 25004 6372 25010 6384
rect 25501 6375 25559 6381
rect 25501 6372 25513 6375
rect 25004 6344 25513 6372
rect 25004 6332 25010 6344
rect 25501 6341 25513 6344
rect 25547 6341 25559 6375
rect 25501 6335 25559 6341
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10778 6304 10784 6316
rect 10735 6276 10784 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10778 6264 10784 6276
rect 10836 6304 10842 6316
rect 11882 6304 11888 6316
rect 10836 6276 11888 6304
rect 10836 6264 10842 6276
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12176 6276 12909 6304
rect 11606 6196 11612 6248
rect 11664 6236 11670 6248
rect 12176 6245 12204 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 13262 6304 13268 6316
rect 13223 6276 13268 6304
rect 12897 6267 12955 6273
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 14550 6304 14556 6316
rect 14511 6276 14556 6304
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16393 6307 16451 6313
rect 16393 6304 16405 6307
rect 15804 6276 16405 6304
rect 15804 6264 15810 6276
rect 16393 6273 16405 6276
rect 16439 6273 16451 6307
rect 16758 6304 16764 6316
rect 16719 6276 16764 6304
rect 16393 6267 16451 6273
rect 16758 6264 16764 6276
rect 16816 6264 16822 6316
rect 18874 6304 18880 6316
rect 18787 6276 18880 6304
rect 18874 6264 18880 6276
rect 18932 6304 18938 6316
rect 23842 6304 23848 6316
rect 18932 6276 20300 6304
rect 23803 6276 23848 6304
rect 18932 6264 18938 6276
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11664 6208 12173 6236
rect 11664 6196 11670 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 16298 6236 16304 6248
rect 16259 6208 16304 6236
rect 12161 6199 12219 6205
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16574 6236 16580 6248
rect 16487 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6236 16638 6248
rect 17586 6236 17592 6248
rect 16632 6208 17592 6236
rect 16632 6196 16638 6208
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 17954 6196 17960 6248
rect 18012 6236 18018 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 18012 6208 18061 6236
rect 18012 6196 18018 6208
rect 18049 6205 18061 6208
rect 18095 6236 18107 6239
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 18095 6208 18521 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 19058 6236 19064 6248
rect 19019 6208 19064 6236
rect 18509 6199 18567 6205
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19242 6196 19248 6248
rect 19300 6236 19306 6248
rect 19521 6239 19579 6245
rect 19521 6236 19533 6239
rect 19300 6208 19533 6236
rect 19300 6196 19306 6208
rect 19521 6205 19533 6208
rect 19567 6205 19579 6239
rect 19978 6236 19984 6248
rect 19939 6208 19984 6236
rect 19521 6199 19579 6205
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20272 6245 20300 6276
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 24118 6264 24124 6316
rect 24176 6304 24182 6316
rect 24489 6307 24547 6313
rect 24489 6304 24501 6307
rect 24176 6276 24501 6304
rect 24176 6264 24182 6276
rect 24489 6273 24501 6276
rect 24535 6304 24547 6307
rect 24762 6304 24768 6316
rect 24535 6276 24768 6304
rect 24535 6273 24547 6276
rect 24489 6267 24547 6273
rect 24762 6264 24768 6276
rect 24820 6264 24826 6316
rect 20257 6239 20315 6245
rect 20257 6205 20269 6239
rect 20303 6205 20315 6239
rect 20257 6199 20315 6205
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6205 21511 6239
rect 21453 6199 21511 6205
rect 9257 6140 10364 6168
rect 9257 6137 9269 6140
rect 9211 6131 9269 6137
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 10836 6140 10881 6168
rect 10836 6128 10842 6140
rect 10962 6128 10968 6180
rect 11020 6168 11026 6180
rect 11333 6171 11391 6177
rect 11333 6168 11345 6171
rect 11020 6140 11345 6168
rect 11020 6128 11026 6140
rect 11333 6137 11345 6140
rect 11379 6137 11391 6171
rect 11333 6131 11391 6137
rect 12986 6128 12992 6180
rect 13044 6168 13050 6180
rect 14461 6171 14519 6177
rect 13044 6140 13089 6168
rect 13044 6128 13050 6140
rect 14461 6137 14473 6171
rect 14507 6168 14519 6171
rect 14915 6171 14973 6177
rect 14915 6168 14927 6171
rect 14507 6140 14927 6168
rect 14507 6137 14519 6140
rect 14461 6131 14519 6137
rect 14915 6137 14927 6140
rect 14961 6168 14973 6171
rect 18690 6168 18696 6180
rect 14961 6140 18696 6168
rect 14961 6137 14973 6140
rect 14915 6131 14973 6137
rect 6638 6100 6644 6112
rect 3743 6072 4108 6100
rect 6599 6072 6644 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6788 6072 6929 6100
rect 6788 6060 6794 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 7929 6103 7987 6109
rect 7929 6100 7941 6103
rect 7892 6072 7941 6100
rect 7892 6060 7898 6072
rect 7929 6069 7941 6072
rect 7975 6100 7987 6103
rect 8294 6100 8300 6112
rect 7975 6072 8300 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 10192 6072 10425 6100
rect 10192 6060 10198 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11422 6100 11428 6112
rect 11112 6072 11428 6100
rect 11112 6060 11118 6072
rect 11422 6060 11428 6072
rect 11480 6100 11486 6112
rect 14476 6100 14504 6131
rect 18690 6128 18696 6140
rect 18748 6128 18754 6180
rect 20533 6171 20591 6177
rect 20533 6137 20545 6171
rect 20579 6168 20591 6171
rect 21174 6168 21180 6180
rect 20579 6140 21180 6168
rect 20579 6137 20591 6140
rect 20533 6131 20591 6137
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 15838 6100 15844 6112
rect 11480 6072 14504 6100
rect 15799 6072 15844 6100
rect 11480 6060 11486 6072
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 18322 6100 18328 6112
rect 18279 6072 18328 6100
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 18322 6060 18328 6072
rect 18380 6100 18386 6112
rect 20070 6100 20076 6112
rect 18380 6072 20076 6100
rect 18380 6060 18386 6072
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 21269 6103 21327 6109
rect 21269 6069 21281 6103
rect 21315 6100 21327 6103
rect 21358 6100 21364 6112
rect 21315 6072 21364 6100
rect 21315 6069 21327 6072
rect 21269 6063 21327 6069
rect 21358 6060 21364 6072
rect 21416 6100 21422 6112
rect 21468 6100 21496 6199
rect 25222 6196 25228 6248
rect 25280 6236 25286 6248
rect 25317 6239 25375 6245
rect 25317 6236 25329 6239
rect 25280 6208 25329 6236
rect 25280 6196 25286 6208
rect 25317 6205 25329 6208
rect 25363 6236 25375 6239
rect 25869 6239 25927 6245
rect 25869 6236 25881 6239
rect 25363 6208 25881 6236
rect 25363 6205 25375 6208
rect 25317 6199 25375 6205
rect 25869 6205 25881 6208
rect 25915 6205 25927 6239
rect 25869 6199 25927 6205
rect 22094 6168 22100 6180
rect 22055 6140 22100 6168
rect 22094 6128 22100 6140
rect 22152 6128 22158 6180
rect 22738 6128 22744 6180
rect 22796 6168 22802 6180
rect 23477 6171 23535 6177
rect 23477 6168 23489 6171
rect 22796 6140 23489 6168
rect 22796 6128 22802 6140
rect 23477 6137 23489 6140
rect 23523 6168 23535 6171
rect 23937 6171 23995 6177
rect 23937 6168 23949 6171
rect 23523 6140 23949 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23937 6137 23949 6140
rect 23983 6168 23995 6171
rect 25038 6168 25044 6180
rect 23983 6140 25044 6168
rect 23983 6137 23995 6140
rect 23937 6131 23995 6137
rect 25038 6128 25044 6140
rect 25096 6128 25102 6180
rect 21416 6072 21496 6100
rect 21416 6060 21422 6072
rect 24670 6060 24676 6112
rect 24728 6100 24734 6112
rect 24765 6103 24823 6109
rect 24765 6100 24777 6103
rect 24728 6072 24777 6100
rect 24728 6060 24734 6072
rect 24765 6069 24777 6072
rect 24811 6069 24823 6103
rect 24765 6063 24823 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2222 5856 2228 5908
rect 2280 5896 2286 5908
rect 3421 5899 3479 5905
rect 3421 5896 3433 5899
rect 2280 5868 3433 5896
rect 2280 5856 2286 5868
rect 3421 5865 3433 5868
rect 3467 5865 3479 5899
rect 4430 5896 4436 5908
rect 4391 5868 4436 5896
rect 3421 5859 3479 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 7190 5896 7196 5908
rect 7151 5868 7196 5896
rect 7190 5856 7196 5868
rect 7248 5896 7254 5908
rect 9122 5896 9128 5908
rect 7248 5868 8984 5896
rect 9083 5868 9128 5896
rect 7248 5856 7254 5868
rect 2593 5831 2651 5837
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 2682 5828 2688 5840
rect 2639 5800 2688 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 5623 5831 5681 5837
rect 5623 5797 5635 5831
rect 5669 5828 5681 5831
rect 6454 5828 6460 5840
rect 5669 5800 6460 5828
rect 5669 5797 5681 5800
rect 5623 5791 5681 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 8199 5831 8257 5837
rect 8199 5797 8211 5831
rect 8245 5828 8257 5831
rect 8754 5828 8760 5840
rect 8245 5800 8760 5828
rect 8245 5797 8257 5800
rect 8199 5791 8257 5797
rect 8754 5788 8760 5800
rect 8812 5788 8818 5840
rect 8956 5828 8984 5868
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9493 5899 9551 5905
rect 9493 5865 9505 5899
rect 9539 5896 9551 5899
rect 9766 5896 9772 5908
rect 9539 5868 9772 5896
rect 9539 5865 9551 5868
rect 9493 5859 9551 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 10229 5899 10287 5905
rect 10229 5865 10241 5899
rect 10275 5896 10287 5899
rect 10686 5896 10692 5908
rect 10275 5868 10692 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11885 5899 11943 5905
rect 11885 5865 11897 5899
rect 11931 5896 11943 5899
rect 14550 5896 14556 5908
rect 11931 5868 12940 5896
rect 14511 5868 14556 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 10778 5828 10784 5840
rect 8956 5800 10784 5828
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 11327 5831 11385 5837
rect 11327 5797 11339 5831
rect 11373 5828 11385 5831
rect 11422 5828 11428 5840
rect 11373 5800 11428 5828
rect 11373 5797 11385 5800
rect 11327 5791 11385 5797
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 12434 5828 12440 5840
rect 12395 5800 12440 5828
rect 12434 5788 12440 5800
rect 12492 5788 12498 5840
rect 12912 5837 12940 5868
rect 14550 5856 14556 5868
rect 14608 5856 14614 5908
rect 15562 5896 15568 5908
rect 15304 5868 15568 5896
rect 12897 5831 12955 5837
rect 12897 5797 12909 5831
rect 12943 5828 12955 5831
rect 13446 5828 13452 5840
rect 12943 5800 13452 5828
rect 12943 5797 12955 5800
rect 12897 5791 12955 5797
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 1118 5720 1124 5772
rect 1176 5760 1182 5772
rect 1432 5763 1490 5769
rect 1432 5760 1444 5763
rect 1176 5732 1444 5760
rect 1176 5720 1182 5732
rect 1432 5729 1444 5732
rect 1478 5729 1490 5763
rect 4246 5760 4252 5772
rect 4159 5732 4252 5760
rect 1432 5723 1490 5729
rect 4246 5720 4252 5732
rect 4304 5760 4310 5772
rect 4304 5732 5902 5760
rect 4304 5720 4310 5732
rect 2498 5692 2504 5704
rect 2459 5664 2504 5692
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 5261 5695 5319 5701
rect 2837 5664 4154 5692
rect 1535 5627 1593 5633
rect 1535 5593 1547 5627
rect 1581 5624 1593 5627
rect 2837 5624 2865 5664
rect 3050 5624 3056 5636
rect 1581 5596 2865 5624
rect 3011 5596 3056 5624
rect 1581 5593 1593 5596
rect 1535 5587 1593 5593
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 4126 5624 4154 5664
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5534 5692 5540 5704
rect 5307 5664 5540 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5874 5692 5902 5732
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7834 5760 7840 5772
rect 7524 5732 7840 5760
rect 7524 5720 7530 5732
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9712 5763 9770 5769
rect 9712 5760 9724 5763
rect 9548 5732 9724 5760
rect 9548 5720 9554 5732
rect 9712 5729 9724 5732
rect 9758 5729 9770 5763
rect 9712 5723 9770 5729
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10928 5732 10977 5760
rect 10928 5720 10934 5732
rect 10965 5729 10977 5732
rect 11011 5760 11023 5763
rect 11514 5760 11520 5772
rect 11011 5732 11520 5760
rect 11011 5729 11023 5732
rect 10965 5723 11023 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 15304 5769 15332 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 16393 5899 16451 5905
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 16574 5896 16580 5908
rect 16439 5868 16580 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 16114 5760 16120 5772
rect 15611 5732 16120 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 16114 5720 16120 5732
rect 16172 5760 16178 5772
rect 16408 5760 16436 5859
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 17037 5899 17095 5905
rect 17037 5865 17049 5899
rect 17083 5896 17095 5899
rect 17126 5896 17132 5908
rect 17083 5868 17132 5896
rect 17083 5865 17095 5868
rect 17037 5859 17095 5865
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 17218 5856 17224 5908
rect 17276 5896 17282 5908
rect 17678 5896 17684 5908
rect 17276 5868 17684 5896
rect 17276 5856 17282 5868
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 19058 5856 19064 5908
rect 19116 5896 19122 5908
rect 19981 5899 20039 5905
rect 19981 5896 19993 5899
rect 19116 5868 19993 5896
rect 19116 5856 19122 5868
rect 19981 5865 19993 5868
rect 20027 5896 20039 5899
rect 20254 5896 20260 5908
rect 20027 5868 20260 5896
rect 20027 5865 20039 5868
rect 19981 5859 20039 5865
rect 20254 5856 20260 5868
rect 20312 5896 20318 5908
rect 20349 5899 20407 5905
rect 20349 5896 20361 5899
rect 20312 5868 20361 5896
rect 20312 5856 20318 5868
rect 20349 5865 20361 5868
rect 20395 5865 20407 5899
rect 22554 5896 22560 5908
rect 22515 5868 22560 5896
rect 20349 5859 20407 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 22830 5856 22836 5908
rect 22888 5896 22894 5908
rect 23109 5899 23167 5905
rect 23109 5896 23121 5899
rect 22888 5868 23121 5896
rect 22888 5856 22894 5868
rect 23109 5865 23121 5868
rect 23155 5865 23167 5899
rect 23842 5896 23848 5908
rect 23803 5868 23848 5896
rect 23109 5859 23167 5865
rect 16850 5760 16856 5772
rect 16172 5732 16436 5760
rect 16811 5732 16856 5760
rect 16172 5720 16178 5732
rect 16850 5720 16856 5732
rect 16908 5720 16914 5772
rect 17144 5760 17172 5856
rect 17310 5828 17316 5840
rect 17271 5800 17316 5828
rect 17310 5788 17316 5800
rect 17368 5828 17374 5840
rect 17954 5828 17960 5840
rect 17368 5800 17960 5828
rect 17368 5788 17374 5800
rect 17954 5788 17960 5800
rect 18012 5828 18018 5840
rect 18049 5831 18107 5837
rect 18049 5828 18061 5831
rect 18012 5800 18061 5828
rect 18012 5788 18018 5800
rect 18049 5797 18061 5800
rect 18095 5828 18107 5831
rect 19705 5831 19763 5837
rect 18095 5800 19104 5828
rect 18095 5797 18107 5800
rect 18049 5791 18107 5797
rect 18230 5760 18236 5772
rect 17144 5732 18236 5760
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 19076 5769 19104 5800
rect 19705 5797 19717 5831
rect 19751 5828 19763 5831
rect 21266 5828 21272 5840
rect 19751 5800 21272 5828
rect 19751 5797 19763 5800
rect 19705 5791 19763 5797
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 23124 5828 23152 5859
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 24305 5831 24363 5837
rect 24305 5828 24317 5831
rect 23124 5800 24317 5828
rect 24305 5797 24317 5800
rect 24351 5828 24363 5831
rect 25222 5828 25228 5840
rect 24351 5800 25228 5828
rect 24351 5797 24363 5800
rect 24305 5791 24363 5797
rect 25222 5788 25228 5800
rect 25280 5788 25286 5840
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5729 18751 5763
rect 18693 5723 18751 5729
rect 19061 5763 19119 5769
rect 19061 5729 19073 5763
rect 19107 5729 19119 5763
rect 19061 5723 19119 5729
rect 9306 5692 9312 5704
rect 5874 5664 9312 5692
rect 9306 5652 9312 5664
rect 9364 5652 9370 5704
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 11112 5664 12633 5692
rect 11112 5652 11118 5664
rect 12621 5661 12633 5664
rect 12667 5692 12679 5695
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12667 5664 12817 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 13081 5695 13139 5701
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13722 5692 13728 5704
rect 13127 5664 13728 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 5442 5624 5448 5636
rect 4126 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 9815 5627 9873 5633
rect 9815 5624 9827 5627
rect 8168 5596 9827 5624
rect 8168 5584 8174 5596
rect 9815 5593 9827 5596
rect 9861 5593 9873 5627
rect 9815 5587 9873 5593
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 13096 5624 13124 5655
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 15654 5692 15660 5704
rect 15427 5664 15660 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 15654 5652 15660 5664
rect 15712 5692 15718 5704
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 15712 5664 16681 5692
rect 15712 5652 15718 5664
rect 16669 5661 16681 5664
rect 16715 5692 16727 5695
rect 17402 5692 17408 5704
rect 16715 5664 17408 5692
rect 16715 5661 16727 5664
rect 16669 5655 16727 5661
rect 17402 5652 17408 5664
rect 17460 5692 17466 5704
rect 18708 5692 18736 5723
rect 19334 5720 19340 5772
rect 19392 5760 19398 5772
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 19392 5732 19441 5760
rect 19392 5720 19398 5732
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 20622 5720 20628 5772
rect 20680 5760 20686 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20680 5732 21097 5760
rect 20680 5720 20686 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 21174 5720 21180 5772
rect 21232 5760 21238 5772
rect 22186 5760 22192 5772
rect 21232 5732 22192 5760
rect 21232 5720 21238 5732
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 22646 5720 22652 5772
rect 22704 5720 22710 5772
rect 17460 5664 18736 5692
rect 22664 5692 22692 5720
rect 24210 5692 24216 5704
rect 22664 5664 23474 5692
rect 24171 5664 24216 5692
rect 17460 5652 17466 5664
rect 10100 5596 13124 5624
rect 21269 5627 21327 5633
rect 10100 5584 10106 5596
rect 21269 5593 21281 5627
rect 21315 5624 21327 5627
rect 22646 5624 22652 5636
rect 21315 5596 22652 5624
rect 21315 5593 21327 5596
rect 21269 5587 21327 5593
rect 22646 5584 22652 5596
rect 22704 5584 22710 5636
rect 23446 5624 23474 5664
rect 24210 5652 24216 5664
rect 24268 5652 24274 5704
rect 24489 5695 24547 5701
rect 24489 5661 24501 5695
rect 24535 5661 24547 5695
rect 24489 5655 24547 5661
rect 24504 5624 24532 5655
rect 24762 5624 24768 5636
rect 23446 5596 24768 5624
rect 24762 5584 24768 5596
rect 24820 5584 24826 5636
rect 2130 5556 2136 5568
rect 2091 5528 2136 5556
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 6181 5559 6239 5565
rect 6181 5556 6193 5559
rect 5408 5528 6193 5556
rect 5408 5516 5414 5528
rect 6181 5525 6193 5528
rect 6227 5525 6239 5559
rect 6822 5556 6828 5568
rect 6783 5528 6828 5556
rect 6181 5519 6239 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8260 5528 8769 5556
rect 8260 5516 8266 5528
rect 8757 5525 8769 5528
rect 8803 5556 8815 5559
rect 10134 5556 10140 5568
rect 8803 5528 10140 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 10134 5516 10140 5528
rect 10192 5556 10198 5568
rect 10318 5556 10324 5568
rect 10192 5528 10324 5556
rect 10192 5516 10198 5528
rect 10318 5516 10324 5528
rect 10376 5556 10382 5568
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 10376 5528 10517 5556
rect 10376 5516 10382 5528
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 10505 5519 10563 5525
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 12158 5556 12164 5568
rect 11112 5528 12164 5556
rect 11112 5516 11118 5528
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 12621 5559 12679 5565
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13725 5559 13783 5565
rect 13725 5556 13737 5559
rect 12667 5528 13737 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13725 5525 13737 5528
rect 13771 5525 13783 5559
rect 21818 5556 21824 5568
rect 21779 5528 21824 5556
rect 13725 5519 13783 5525
rect 21818 5516 21824 5528
rect 21876 5516 21882 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1118 5312 1124 5364
rect 1176 5352 1182 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1176 5324 1593 5352
rect 1176 5312 1182 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1854 5312 1860 5364
rect 1912 5352 1918 5364
rect 1949 5355 2007 5361
rect 1949 5352 1961 5355
rect 1912 5324 1961 5352
rect 1912 5312 1918 5324
rect 1949 5321 1961 5324
rect 1995 5321 2007 5355
rect 1949 5315 2007 5321
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4246 5352 4252 5364
rect 4111 5324 4252 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 4479 5324 4721 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4709 5321 4721 5324
rect 4755 5352 4767 5355
rect 6362 5352 6368 5364
rect 4755 5324 6368 5352
rect 4755 5321 4767 5324
rect 4709 5315 4767 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 9490 5352 9496 5364
rect 8076 5324 9496 5352
rect 8076 5312 8082 5324
rect 9490 5312 9496 5324
rect 9548 5352 9554 5364
rect 9677 5355 9735 5361
rect 9677 5352 9689 5355
rect 9548 5324 9689 5352
rect 9548 5312 9554 5324
rect 9677 5321 9689 5324
rect 9723 5321 9735 5355
rect 9677 5315 9735 5321
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 11514 5352 11520 5364
rect 9916 5324 11421 5352
rect 11475 5324 11520 5352
rect 9916 5312 9922 5324
rect 3142 5244 3148 5296
rect 3200 5284 3206 5296
rect 5626 5284 5632 5296
rect 3200 5256 5632 5284
rect 3200 5244 3206 5256
rect 5626 5244 5632 5256
rect 5684 5284 5690 5296
rect 5813 5287 5871 5293
rect 5813 5284 5825 5287
rect 5684 5256 5825 5284
rect 5684 5244 5690 5256
rect 5813 5253 5825 5256
rect 5859 5253 5871 5287
rect 5813 5247 5871 5253
rect 9766 5244 9772 5296
rect 9824 5284 9830 5296
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 9824 5256 10793 5284
rect 9824 5244 9830 5256
rect 10781 5253 10793 5256
rect 10827 5284 10839 5287
rect 10870 5284 10876 5296
rect 10827 5256 10876 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11393 5284 11421 5324
rect 11514 5312 11520 5324
rect 11572 5312 11578 5364
rect 13446 5352 13452 5364
rect 13407 5324 13452 5352
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15562 5352 15568 5364
rect 15427 5324 15568 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 17402 5352 17408 5364
rect 17363 5324 17408 5352
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 18230 5352 18236 5364
rect 18191 5324 18236 5352
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18782 5352 18788 5364
rect 18743 5324 18788 5352
rect 18782 5312 18788 5324
rect 18840 5312 18846 5364
rect 21082 5352 21088 5364
rect 21043 5324 21088 5352
rect 21082 5312 21088 5324
rect 21140 5312 21146 5364
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21729 5355 21787 5361
rect 21729 5352 21741 5355
rect 21324 5324 21741 5352
rect 21324 5312 21330 5324
rect 21729 5321 21741 5324
rect 21775 5352 21787 5355
rect 22554 5352 22560 5364
rect 21775 5324 22560 5352
rect 21775 5321 21787 5324
rect 21729 5315 21787 5321
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 11393 5256 12173 5284
rect 12161 5253 12173 5256
rect 12207 5253 12219 5287
rect 14642 5284 14648 5296
rect 14603 5256 14648 5284
rect 12161 5247 12219 5253
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 4062 5216 4068 5228
rect 3108 5188 4068 5216
rect 3108 5176 3114 5188
rect 4062 5176 4068 5188
rect 4120 5216 4126 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4120 5188 5273 5216
rect 4120 5176 4126 5188
rect 5261 5185 5273 5188
rect 5307 5216 5319 5219
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5307 5188 6193 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 6181 5185 6193 5188
rect 6227 5216 6239 5219
rect 7193 5219 7251 5225
rect 7193 5216 7205 5219
rect 6227 5188 7205 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 7193 5185 7205 5188
rect 7239 5185 7251 5219
rect 7193 5179 7251 5185
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8570 5216 8576 5228
rect 8435 5188 8576 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5216 10287 5219
rect 10686 5216 10692 5228
rect 10275 5188 10692 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11241 5219 11299 5225
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11422 5216 11428 5228
rect 11287 5188 11428 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4433 5151 4491 5157
rect 4433 5148 4445 5151
rect 4203 5120 4445 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4433 5117 4445 5120
rect 4479 5117 4491 5151
rect 12176 5148 12204 5247
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 15580 5284 15608 5312
rect 17773 5287 17831 5293
rect 17773 5284 17785 5287
rect 15580 5256 17785 5284
rect 17773 5253 17785 5256
rect 17819 5253 17831 5287
rect 17773 5247 17831 5253
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13320 5188 13814 5216
rect 13320 5176 13326 5188
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12176 5120 12449 5148
rect 4433 5111 4491 5117
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12768 5120 12909 5148
rect 12768 5108 12774 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 1854 5040 1860 5092
rect 1912 5080 1918 5092
rect 2222 5080 2228 5092
rect 1912 5052 2228 5080
rect 1912 5040 1918 5052
rect 2222 5040 2228 5052
rect 2280 5080 2286 5092
rect 2454 5083 2512 5089
rect 2454 5080 2466 5083
rect 2280 5052 2466 5080
rect 2280 5040 2286 5052
rect 2454 5049 2466 5052
rect 2500 5049 2512 5083
rect 2454 5043 2512 5049
rect 2682 5040 2688 5092
rect 2740 5080 2746 5092
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 2740 5052 3341 5080
rect 2740 5040 2746 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 4522 5080 4528 5092
rect 3329 5043 3387 5049
rect 4356 5052 4528 5080
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 4356 5021 4384 5052
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 5350 5040 5356 5092
rect 5408 5080 5414 5092
rect 5408 5052 5453 5080
rect 5408 5040 5414 5052
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6914 5080 6920 5092
rect 6052 5052 6920 5080
rect 6052 5040 6058 5052
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5049 7067 5083
rect 10318 5080 10324 5092
rect 10279 5052 10324 5080
rect 7009 5043 7067 5049
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2648 4984 3065 5012
rect 2648 4972 2654 4984
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 4981 4399 5015
rect 4341 4975 4399 4981
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 6362 5012 6368 5024
rect 5123 4984 6368 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6546 4972 6552 5024
rect 6604 5012 6610 5024
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 6604 4984 6653 5012
rect 6604 4972 6610 4984
rect 6641 4981 6653 4984
rect 6687 5012 6699 5015
rect 7024 5012 7052 5043
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 11606 5040 11612 5092
rect 11664 5080 11670 5092
rect 13786 5080 13814 5188
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 15436 5120 15669 5148
rect 15436 5108 15442 5120
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 14090 5080 14096 5092
rect 11664 5052 12480 5080
rect 13786 5052 14096 5080
rect 11664 5040 11670 5052
rect 6687 4984 7052 5012
rect 7929 5015 7987 5021
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 7975 4984 8309 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8297 4981 8309 4984
rect 8343 5012 8355 5015
rect 8754 5012 8760 5024
rect 8343 4984 8760 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9306 5012 9312 5024
rect 9267 4984 9312 5012
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 12452 5012 12480 5052
rect 14090 5040 14096 5052
rect 14148 5040 14154 5092
rect 14185 5083 14243 5089
rect 14185 5049 14197 5083
rect 14231 5049 14243 5083
rect 15565 5083 15623 5089
rect 15565 5080 15577 5083
rect 14185 5043 14243 5049
rect 14936 5052 15577 5080
rect 12529 5015 12587 5021
rect 12529 5012 12541 5015
rect 12452 4984 12541 5012
rect 12529 4981 12541 4984
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 13909 5015 13967 5021
rect 13909 4981 13921 5015
rect 13955 5012 13967 5015
rect 14200 5012 14228 5043
rect 14936 5012 14964 5052
rect 15565 5049 15577 5052
rect 15611 5049 15623 5083
rect 15565 5043 15623 5049
rect 16850 5040 16856 5092
rect 16908 5080 16914 5092
rect 16945 5083 17003 5089
rect 16945 5080 16957 5083
rect 16908 5052 16957 5080
rect 16908 5040 16914 5052
rect 16945 5049 16957 5052
rect 16991 5080 17003 5083
rect 17494 5080 17500 5092
rect 16991 5052 17500 5080
rect 16991 5049 17003 5052
rect 16945 5043 17003 5049
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 17788 5024 17816 5247
rect 18800 5216 18828 5312
rect 20441 5219 20499 5225
rect 18800 5188 20208 5216
rect 19058 5148 19064 5160
rect 19019 5120 19064 5148
rect 19058 5108 19064 5120
rect 19116 5108 19122 5160
rect 19705 5151 19763 5157
rect 19705 5117 19717 5151
rect 19751 5117 19763 5151
rect 19978 5148 19984 5160
rect 19939 5120 19984 5148
rect 19705 5111 19763 5117
rect 19426 5040 19432 5092
rect 19484 5080 19490 5092
rect 19720 5080 19748 5111
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20180 5157 20208 5188
rect 20441 5185 20453 5219
rect 20487 5216 20499 5219
rect 21818 5216 21824 5228
rect 20487 5188 21824 5216
rect 20487 5185 20499 5188
rect 20441 5179 20499 5185
rect 21818 5176 21824 5188
rect 21876 5176 21882 5228
rect 20165 5151 20223 5157
rect 20165 5117 20177 5151
rect 20211 5117 20223 5151
rect 20165 5111 20223 5117
rect 22157 5089 22185 5324
rect 22554 5312 22560 5324
rect 22612 5312 22618 5364
rect 22738 5352 22744 5364
rect 22699 5324 22744 5352
rect 22738 5312 22744 5324
rect 22796 5312 22802 5364
rect 23382 5312 23388 5364
rect 23440 5352 23446 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23440 5324 24041 5352
rect 23440 5312 23446 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24029 5315 24087 5321
rect 22572 5284 22600 5312
rect 23017 5287 23075 5293
rect 23017 5284 23029 5287
rect 22572 5256 23029 5284
rect 23017 5253 23029 5256
rect 23063 5253 23075 5287
rect 24044 5284 24072 5315
rect 24210 5312 24216 5364
rect 24268 5352 24274 5364
rect 25222 5352 25228 5364
rect 24268 5324 24624 5352
rect 25183 5324 25228 5352
rect 24268 5312 24274 5324
rect 24394 5284 24400 5296
rect 24044 5256 24400 5284
rect 23017 5247 23075 5253
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 24596 5284 24624 5324
rect 25222 5312 25228 5324
rect 25280 5312 25286 5364
rect 25593 5287 25651 5293
rect 25593 5284 25605 5287
rect 24596 5256 25605 5284
rect 25593 5253 25605 5256
rect 25639 5253 25651 5287
rect 25593 5247 25651 5253
rect 24762 5216 24768 5228
rect 24723 5188 24768 5216
rect 24762 5176 24768 5188
rect 24820 5176 24826 5228
rect 20717 5083 20775 5089
rect 20717 5080 20729 5083
rect 19484 5052 20729 5080
rect 19484 5040 19490 5052
rect 20717 5049 20729 5052
rect 20763 5049 20775 5083
rect 20717 5043 20775 5049
rect 22142 5083 22200 5089
rect 22142 5049 22154 5083
rect 22188 5049 22200 5083
rect 22142 5043 22200 5049
rect 23477 5083 23535 5089
rect 23477 5049 23489 5083
rect 23523 5080 23535 5083
rect 24305 5083 24363 5089
rect 24305 5080 24317 5083
rect 23523 5052 24317 5080
rect 23523 5049 23535 5052
rect 23477 5043 23535 5049
rect 24305 5049 24317 5052
rect 24351 5049 24363 5083
rect 24305 5043 24363 5049
rect 17770 5012 17776 5024
rect 13955 4984 14964 5012
rect 17683 4984 17776 5012
rect 13955 4981 13967 4984
rect 13909 4975 13967 4981
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 19978 5012 19984 5024
rect 17828 4984 19984 5012
rect 17828 4972 17834 4984
rect 19978 4972 19984 4984
rect 20036 4972 20042 5024
rect 24320 5012 24348 5043
rect 24394 5040 24400 5092
rect 24452 5080 24458 5092
rect 24452 5052 24497 5080
rect 24452 5040 24458 5052
rect 25130 5012 25136 5024
rect 24320 4984 25136 5012
rect 25130 4972 25136 4984
rect 25188 4972 25194 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1535 4811 1593 4817
rect 1535 4777 1547 4811
rect 1581 4808 1593 4811
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1581 4780 1961 4808
rect 1581 4777 1593 4780
rect 1535 4771 1593 4777
rect 1949 4777 1961 4780
rect 1995 4808 2007 4811
rect 2498 4808 2504 4820
rect 1995 4780 2504 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 5534 4808 5540 4820
rect 5495 4780 5540 4808
rect 5534 4768 5540 4780
rect 5592 4808 5598 4820
rect 5902 4808 5908 4820
rect 5592 4780 5908 4808
rect 5592 4768 5598 4780
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6914 4808 6920 4820
rect 6875 4780 6920 4808
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7834 4808 7840 4820
rect 7795 4780 7840 4808
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8570 4768 8576 4820
rect 8628 4808 8634 4820
rect 9033 4811 9091 4817
rect 9033 4808 9045 4811
rect 8628 4780 9045 4808
rect 8628 4768 8634 4780
rect 9033 4777 9045 4780
rect 9079 4777 9091 4811
rect 9033 4771 9091 4777
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11333 4811 11391 4817
rect 11333 4808 11345 4811
rect 11296 4780 11345 4808
rect 11296 4768 11302 4780
rect 11333 4777 11345 4780
rect 11379 4777 11391 4811
rect 12894 4808 12900 4820
rect 12855 4780 12900 4808
rect 11333 4771 11391 4777
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 14090 4808 14096 4820
rect 14051 4780 14096 4808
rect 14090 4768 14096 4780
rect 14148 4768 14154 4820
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 16393 4811 16451 4817
rect 16393 4808 16405 4811
rect 15436 4780 16405 4808
rect 15436 4768 15442 4780
rect 16393 4777 16405 4780
rect 16439 4777 16451 4811
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 16393 4771 16451 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17954 4808 17960 4820
rect 17915 4780 17960 4808
rect 17954 4768 17960 4780
rect 18012 4808 18018 4820
rect 18966 4808 18972 4820
rect 18012 4780 18972 4808
rect 18012 4768 18018 4780
rect 18966 4768 18972 4780
rect 19024 4768 19030 4820
rect 19334 4768 19340 4820
rect 19392 4808 19398 4820
rect 19889 4811 19947 4817
rect 19889 4808 19901 4811
rect 19392 4780 19901 4808
rect 19392 4768 19398 4780
rect 19889 4777 19901 4780
rect 19935 4777 19947 4811
rect 20622 4808 20628 4820
rect 20583 4780 20628 4808
rect 19889 4771 19947 4777
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 21266 4808 21272 4820
rect 21227 4780 21272 4808
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 22186 4808 22192 4820
rect 22147 4780 22192 4808
rect 22186 4768 22192 4780
rect 22244 4768 22250 4820
rect 24118 4808 24124 4820
rect 24079 4780 24124 4808
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 24670 4808 24676 4820
rect 24631 4780 24676 4808
rect 24670 4768 24676 4780
rect 24728 4768 24734 4820
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2590 4740 2596 4752
rect 2363 4712 2596 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 2590 4700 2596 4712
rect 2648 4700 2654 4752
rect 3142 4740 3148 4752
rect 3103 4712 3148 4740
rect 3142 4700 3148 4712
rect 3200 4700 3206 4752
rect 3970 4700 3976 4752
rect 4028 4740 4034 4752
rect 4146 4743 4204 4749
rect 4146 4740 4158 4743
rect 4028 4712 4158 4740
rect 4028 4700 4034 4712
rect 4146 4709 4158 4712
rect 4192 4709 4204 4743
rect 4146 4703 4204 4709
rect 4258 4743 4316 4749
rect 4258 4709 4270 4743
rect 4304 4740 4316 4743
rect 4614 4740 4620 4752
rect 4304 4712 4620 4740
rect 4304 4709 4316 4712
rect 4258 4703 4316 4709
rect 4614 4700 4620 4712
rect 4672 4700 4678 4752
rect 6083 4743 6141 4749
rect 6083 4709 6095 4743
rect 6129 4740 6141 4743
rect 6454 4740 6460 4752
rect 6129 4712 6460 4740
rect 6129 4709 6141 4712
rect 6083 4703 6141 4709
rect 6454 4700 6460 4712
rect 6512 4700 6518 4752
rect 7561 4743 7619 4749
rect 7561 4709 7573 4743
rect 7607 4740 7619 4743
rect 8110 4740 8116 4752
rect 7607 4712 8116 4740
rect 7607 4709 7619 4712
rect 7561 4703 7619 4709
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 8260 4712 8305 4740
rect 8260 4700 8266 4712
rect 9306 4700 9312 4752
rect 9364 4740 9370 4752
rect 9766 4740 9772 4752
rect 9364 4712 9772 4740
rect 9364 4700 9370 4712
rect 9766 4700 9772 4712
rect 9824 4740 9830 4752
rect 9861 4743 9919 4749
rect 9861 4740 9873 4743
rect 9824 4712 9873 4740
rect 9824 4700 9830 4712
rect 9861 4709 9873 4712
rect 9907 4709 9919 4743
rect 9861 4703 9919 4709
rect 10778 4700 10784 4752
rect 10836 4740 10842 4752
rect 12437 4743 12495 4749
rect 12437 4740 12449 4743
rect 10836 4712 12449 4740
rect 10836 4700 10842 4712
rect 11716 4684 11744 4712
rect 12437 4709 12449 4712
rect 12483 4740 12495 4743
rect 12710 4740 12716 4752
rect 12483 4712 12716 4740
rect 12483 4709 12495 4712
rect 12437 4703 12495 4709
rect 12710 4700 12716 4712
rect 12768 4740 12774 4752
rect 17034 4740 17040 4752
rect 12768 4712 13308 4740
rect 12768 4700 12774 4712
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1762 4672 1768 4684
rect 1510 4644 1768 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4641 11299 4675
rect 11698 4672 11704 4684
rect 11611 4644 11704 4672
rect 11241 4635 11299 4641
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 3142 4604 3148 4616
rect 2547 4576 3148 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 3142 4564 3148 4576
rect 3200 4604 3206 4616
rect 3421 4607 3479 4613
rect 3421 4604 3433 4607
rect 3200 4576 3433 4604
rect 3200 4564 3206 4576
rect 3421 4573 3433 4576
rect 3467 4604 3479 4607
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 3467 4576 4445 4604
rect 3467 4573 3479 4576
rect 3421 4567 3479 4573
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6638 4604 6644 4616
rect 5767 4576 6644 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 8754 4604 8760 4616
rect 8667 4576 8760 4604
rect 8754 4564 8760 4576
rect 8812 4604 8818 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8812 4576 9413 4604
rect 8812 4564 8818 4576
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9490 4564 9496 4616
rect 9548 4604 9554 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9548 4576 9781 4604
rect 9548 4564 9554 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 10042 4604 10048 4616
rect 10003 4576 10048 4604
rect 9769 4567 9827 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 11256 4536 11284 4635
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 13280 4681 13308 4712
rect 15580 4712 17040 4740
rect 15580 4684 15608 4712
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 17696 4740 17724 4768
rect 20349 4743 20407 4749
rect 17696 4712 19380 4740
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4641 13323 4675
rect 15562 4672 15568 4684
rect 15523 4644 15568 4672
rect 13265 4635 13323 4641
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 16669 4675 16727 4681
rect 16669 4672 16681 4675
rect 15712 4644 16681 4672
rect 15712 4632 15718 4644
rect 16669 4641 16681 4644
rect 16715 4641 16727 4675
rect 18230 4672 18236 4684
rect 18191 4644 18236 4672
rect 16669 4635 16727 4641
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 15746 4604 15752 4616
rect 15151 4576 15752 4604
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 16114 4604 16120 4616
rect 16075 4576 16120 4604
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 11330 4536 11336 4548
rect 4580 4508 11336 4536
rect 4580 4496 4586 4508
rect 11330 4496 11336 4508
rect 11388 4496 11394 4548
rect 14737 4539 14795 4545
rect 14737 4505 14749 4539
rect 14783 4536 14795 4539
rect 16574 4536 16580 4548
rect 14783 4508 16580 4536
rect 14783 4505 14795 4508
rect 14737 4499 14795 4505
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 16684 4536 16712 4635
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4641 18659 4675
rect 18966 4672 18972 4684
rect 18927 4644 18972 4672
rect 18601 4635 18659 4641
rect 17310 4604 17316 4616
rect 17271 4576 17316 4604
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 18616 4604 18644 4635
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19352 4681 19380 4712
rect 20349 4709 20361 4743
rect 20395 4740 20407 4743
rect 21082 4740 21088 4752
rect 20395 4712 21088 4740
rect 20395 4709 20407 4712
rect 20349 4703 20407 4709
rect 21082 4700 21088 4712
rect 21140 4700 21146 4752
rect 21910 4700 21916 4752
rect 21968 4740 21974 4752
rect 22554 4740 22560 4752
rect 21968 4712 22560 4740
rect 21968 4700 21974 4712
rect 22554 4700 22560 4712
rect 22612 4740 22618 4752
rect 22741 4743 22799 4749
rect 22741 4740 22753 4743
rect 22612 4712 22753 4740
rect 22612 4700 22618 4712
rect 22741 4709 22753 4712
rect 22787 4709 22799 4743
rect 22741 4703 22799 4709
rect 22830 4700 22836 4752
rect 22888 4740 22894 4752
rect 22888 4712 22933 4740
rect 22888 4700 22894 4712
rect 19337 4675 19395 4681
rect 19337 4641 19349 4675
rect 19383 4641 19395 4675
rect 19337 4635 19395 4641
rect 24857 4675 24915 4681
rect 24857 4641 24869 4675
rect 24903 4672 24915 4675
rect 25038 4672 25044 4684
rect 24903 4644 25044 4672
rect 24903 4641 24915 4644
rect 24857 4635 24915 4641
rect 25038 4632 25044 4644
rect 25096 4632 25102 4684
rect 17460 4576 18644 4604
rect 19613 4607 19671 4613
rect 17460 4564 17466 4576
rect 19613 4573 19625 4607
rect 19659 4604 19671 4607
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 19659 4576 20913 4604
rect 19659 4573 19671 4576
rect 19613 4567 19671 4573
rect 20901 4573 20913 4576
rect 20947 4604 20959 4607
rect 21082 4604 21088 4616
rect 20947 4576 21088 4604
rect 20947 4573 20959 4576
rect 20901 4567 20959 4573
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 22002 4564 22008 4616
rect 22060 4604 22066 4616
rect 23017 4607 23075 4613
rect 23017 4604 23029 4607
rect 22060 4576 23029 4604
rect 22060 4564 22066 4576
rect 23017 4573 23029 4576
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 21821 4539 21879 4545
rect 21821 4536 21833 4539
rect 16684 4508 21833 4536
rect 21821 4505 21833 4508
rect 21867 4505 21879 4539
rect 21821 4499 21879 4505
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 6641 4471 6699 4477
rect 6641 4468 6653 4471
rect 5408 4440 6653 4468
rect 5408 4428 5414 4440
rect 6641 4437 6653 4440
rect 6687 4437 6699 4471
rect 6641 4431 6699 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 13078 4468 13084 4480
rect 8352 4440 13084 4468
rect 8352 4428 8358 4440
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 15746 4468 15752 4480
rect 15707 4440 15752 4468
rect 15746 4428 15752 4440
rect 15804 4428 15810 4480
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 19150 4468 19156 4480
rect 16356 4440 19156 4468
rect 16356 4428 16362 4440
rect 19150 4428 19156 4440
rect 19208 4428 19214 4480
rect 21836 4468 21864 4499
rect 22462 4496 22468 4548
rect 22520 4536 22526 4548
rect 22646 4536 22652 4548
rect 22520 4508 22652 4536
rect 22520 4496 22526 4508
rect 22646 4496 22652 4508
rect 22704 4496 22710 4548
rect 22830 4468 22836 4480
rect 21836 4440 22836 4468
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 4028 4236 4445 4264
rect 4028 4224 4034 4236
rect 4433 4233 4445 4236
rect 4479 4233 4491 4267
rect 4433 4227 4491 4233
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 8202 4264 8208 4276
rect 7239 4236 8208 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 9766 4264 9772 4276
rect 9727 4236 9772 4264
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 11330 4264 11336 4276
rect 11291 4236 11336 4264
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 11698 4264 11704 4276
rect 11659 4236 11704 4264
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 13078 4224 13084 4276
rect 13136 4264 13142 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 13136 4236 13461 4264
rect 13136 4224 13142 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 16482 4264 16488 4276
rect 15804 4236 16488 4264
rect 15804 4224 15810 4236
rect 16482 4224 16488 4236
rect 16540 4264 16546 4276
rect 17126 4264 17132 4276
rect 16540 4236 17132 4264
rect 16540 4224 16546 4236
rect 17126 4224 17132 4236
rect 17184 4224 17190 4276
rect 17402 4264 17408 4276
rect 17363 4236 17408 4264
rect 17402 4224 17408 4236
rect 17460 4224 17466 4276
rect 17770 4264 17776 4276
rect 17731 4236 17776 4264
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 18230 4264 18236 4276
rect 18191 4236 18236 4264
rect 18230 4224 18236 4236
rect 18288 4224 18294 4276
rect 20162 4224 20168 4276
rect 20220 4264 20226 4276
rect 22462 4264 22468 4276
rect 20220 4236 22468 4264
rect 20220 4224 20226 4236
rect 22462 4224 22468 4236
rect 22520 4224 22526 4276
rect 22554 4224 22560 4276
rect 22612 4264 22618 4276
rect 23385 4267 23443 4273
rect 23385 4264 23397 4267
rect 22612 4236 23397 4264
rect 22612 4224 22618 4236
rect 23385 4233 23397 4236
rect 23431 4233 23443 4267
rect 25038 4264 25044 4276
rect 24999 4236 25044 4264
rect 23385 4227 23443 4233
rect 25038 4224 25044 4236
rect 25096 4224 25102 4276
rect 26142 4264 26148 4276
rect 26103 4236 26148 4264
rect 26142 4224 26148 4236
rect 26200 4224 26206 4276
rect 1762 4156 1768 4208
rect 1820 4196 1826 4208
rect 1857 4199 1915 4205
rect 1857 4196 1869 4199
rect 1820 4168 1869 4196
rect 1820 4156 1826 4168
rect 1857 4165 1869 4168
rect 1903 4165 1915 4199
rect 1857 4159 1915 4165
rect 2222 4156 2228 4208
rect 2280 4196 2286 4208
rect 2409 4199 2467 4205
rect 2409 4196 2421 4199
rect 2280 4168 2421 4196
rect 2280 4156 2286 4168
rect 2409 4165 2421 4168
rect 2455 4165 2467 4199
rect 3418 4196 3424 4208
rect 3379 4168 3424 4196
rect 2409 4159 2467 4165
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 6273 4199 6331 4205
rect 6273 4165 6285 4199
rect 6319 4196 6331 4199
rect 6454 4196 6460 4208
rect 6319 4168 6460 4196
rect 6319 4165 6331 4168
rect 6273 4159 6331 4165
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 7742 4196 7748 4208
rect 7655 4168 7748 4196
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 9490 4196 9496 4208
rect 8772 4168 9496 4196
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 5534 4128 5540 4140
rect 2372 4100 2865 4128
rect 5495 4100 5540 4128
rect 2372 4088 2378 4100
rect 1464 4063 1522 4069
rect 1464 4029 1476 4063
rect 1510 4060 1522 4063
rect 1854 4060 1860 4072
rect 1510 4032 1860 4060
rect 1510 4029 1522 4032
rect 1464 4023 1522 4029
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 1535 3927 1593 3933
rect 1535 3893 1547 3927
rect 1581 3924 1593 3927
rect 2314 3924 2320 3936
rect 1581 3896 2320 3924
rect 1581 3893 1593 3896
rect 1535 3887 1593 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2516 3924 2544 4023
rect 2837 4001 2865 4100
rect 5534 4088 5540 4100
rect 5592 4088 5598 4140
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 4430 4060 4436 4072
rect 4203 4032 4436 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 4430 4020 4436 4032
rect 4488 4020 4494 4072
rect 6638 4060 6644 4072
rect 6599 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7352 4063 7410 4069
rect 7352 4029 7364 4063
rect 7398 4060 7410 4063
rect 7760 4060 7788 4156
rect 8772 4140 8800 4168
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 14277 4199 14335 4205
rect 14277 4165 14289 4199
rect 14323 4196 14335 4199
rect 14458 4196 14464 4208
rect 14323 4168 14464 4196
rect 14323 4165 14335 4168
rect 14277 4159 14335 4165
rect 14458 4156 14464 4168
rect 14516 4156 14522 4208
rect 22830 4156 22836 4208
rect 22888 4196 22894 4208
rect 23017 4199 23075 4205
rect 23017 4196 23029 4199
rect 22888 4168 23029 4196
rect 22888 4156 22894 4168
rect 23017 4165 23029 4168
rect 23063 4165 23075 4199
rect 23017 4159 23075 4165
rect 23106 4156 23112 4208
rect 23164 4196 23170 4208
rect 23164 4168 24440 4196
rect 23164 4156 23170 4168
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9824 4100 10057 4128
rect 9824 4088 9830 4100
rect 10045 4097 10057 4100
rect 10091 4128 10103 4131
rect 10134 4128 10140 4140
rect 10091 4100 10140 4128
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10134 4088 10140 4100
rect 10192 4088 10198 4140
rect 18322 4128 18328 4140
rect 12728 4100 18328 4128
rect 7398 4032 7788 4060
rect 9401 4063 9459 4069
rect 7398 4029 7410 4032
rect 7352 4023 7410 4029
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 12250 4060 12256 4072
rect 9447 4032 10180 4060
rect 12163 4032 12256 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 2822 3995 2880 4001
rect 2822 3961 2834 3995
rect 2868 3992 2880 3995
rect 3602 3992 3608 4004
rect 2868 3964 3608 3992
rect 2868 3961 2880 3964
rect 2822 3955 2880 3961
rect 3602 3952 3608 3964
rect 3660 3952 3666 4004
rect 5258 3992 5264 4004
rect 5219 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5408 3964 5453 3992
rect 5408 3952 5414 3964
rect 7742 3952 7748 4004
rect 7800 3992 7806 4004
rect 8389 3995 8447 4001
rect 8389 3992 8401 3995
rect 7800 3964 8401 3992
rect 7800 3952 7806 3964
rect 8389 3961 8401 3964
rect 8435 3961 8447 3995
rect 8389 3955 8447 3961
rect 8481 3995 8539 4001
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 9766 3992 9772 4004
rect 8527 3964 9772 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 3786 3924 3792 3936
rect 2516 3896 3792 3924
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5368 3924 5396 3952
rect 5123 3896 5396 3924
rect 7423 3927 7481 3933
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 7423 3893 7435 3927
rect 7469 3924 7481 3927
rect 7926 3924 7932 3936
rect 7469 3896 7932 3924
rect 7469 3893 7481 3896
rect 7423 3887 7481 3893
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8496 3924 8524 3955
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 10152 3992 10180 4032
rect 12250 4020 12256 4032
rect 12308 4060 12314 4072
rect 12728 4069 12756 4100
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 19058 4128 19064 4140
rect 18984 4100 19064 4128
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 12308 4032 12725 4060
rect 12308 4020 12314 4032
rect 12713 4029 12725 4032
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 14458 4060 14464 4072
rect 14419 4032 14464 4060
rect 12897 4023 12955 4029
rect 10318 3992 10324 4004
rect 10152 3964 10324 3992
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3961 10471 3995
rect 10962 3992 10968 4004
rect 10923 3964 10968 3992
rect 10413 3955 10471 3961
rect 8251 3896 8524 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10428 3924 10456 3955
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 11698 3952 11704 4004
rect 11756 3992 11762 4004
rect 12912 3992 12940 4023
rect 14458 4020 14464 4032
rect 14516 4020 14522 4072
rect 16301 4063 16359 4069
rect 16301 4029 16313 4063
rect 16347 4060 16359 4063
rect 16574 4060 16580 4072
rect 16347 4032 16580 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16574 4020 16580 4032
rect 16632 4060 16638 4072
rect 16850 4060 16856 4072
rect 16632 4032 16856 4060
rect 16632 4020 16638 4032
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 18984 4069 19012 4100
rect 19058 4088 19064 4100
rect 19116 4088 19122 4140
rect 24118 4128 24124 4140
rect 24079 4100 24124 4128
rect 24118 4088 24124 4100
rect 24176 4088 24182 4140
rect 24412 4128 24440 4168
rect 24412 4100 24808 4128
rect 18969 4063 19027 4069
rect 18969 4029 18981 4063
rect 19015 4029 19027 4063
rect 19426 4060 19432 4072
rect 19387 4032 19432 4060
rect 18969 4023 19027 4029
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 19978 4060 19984 4072
rect 19939 4032 19984 4060
rect 19978 4020 19984 4032
rect 20036 4020 20042 4072
rect 20165 4063 20223 4069
rect 20165 4029 20177 4063
rect 20211 4029 20223 4063
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 20165 4023 20223 4029
rect 21284 4032 21833 4060
rect 20180 3992 20208 4023
rect 21284 4001 21312 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 22787 4032 23474 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 11756 3964 13814 3992
rect 11756 3952 11762 3964
rect 13786 3936 13814 3964
rect 18892 3964 20208 3992
rect 20441 3995 20499 4001
rect 18892 3936 18920 3964
rect 20441 3961 20453 3995
rect 20487 3992 20499 3995
rect 21269 3995 21327 4001
rect 21269 3992 21281 3995
rect 20487 3964 21281 3992
rect 20487 3961 20499 3964
rect 20441 3955 20499 3961
rect 21269 3961 21281 3964
rect 21315 3961 21327 3995
rect 22142 3995 22200 4001
rect 22142 3992 22154 3995
rect 21269 3955 21327 3961
rect 21652 3964 22154 3992
rect 12526 3924 12532 3936
rect 10192 3896 10456 3924
rect 12487 3896 12532 3924
rect 10192 3884 10198 3896
rect 12526 3884 12532 3896
rect 12584 3884 12590 3936
rect 13786 3896 13820 3936
rect 13814 3884 13820 3896
rect 13872 3924 13878 3936
rect 14826 3924 14832 3936
rect 13872 3896 13917 3924
rect 14787 3896 14832 3924
rect 13872 3884 13878 3896
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 15562 3924 15568 3936
rect 15523 3896 15568 3924
rect 15562 3884 15568 3896
rect 15620 3884 15626 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 18874 3924 18880 3936
rect 18835 3896 18880 3924
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20772 3896 20913 3924
rect 20772 3884 20778 3896
rect 20901 3893 20913 3896
rect 20947 3924 20959 3927
rect 21174 3924 21180 3936
rect 20947 3896 21180 3924
rect 20947 3893 20959 3896
rect 20901 3887 20959 3893
rect 21174 3884 21180 3896
rect 21232 3924 21238 3936
rect 21652 3933 21680 3964
rect 22142 3961 22154 3964
rect 22188 3961 22200 3995
rect 22142 3955 22200 3961
rect 21637 3927 21695 3933
rect 21637 3924 21649 3927
rect 21232 3896 21649 3924
rect 21232 3884 21238 3896
rect 21637 3893 21649 3896
rect 21683 3893 21695 3927
rect 23446 3924 23474 4032
rect 24780 4004 24808 4100
rect 25660 4063 25718 4069
rect 25660 4029 25672 4063
rect 25706 4060 25718 4063
rect 26142 4060 26148 4072
rect 25706 4032 26148 4060
rect 25706 4029 25718 4032
rect 25660 4023 25718 4029
rect 26142 4020 26148 4032
rect 26200 4020 26206 4072
rect 24213 3995 24271 4001
rect 24213 3961 24225 3995
rect 24259 3961 24271 3995
rect 24762 3992 24768 4004
rect 24723 3964 24768 3992
rect 24213 3955 24271 3961
rect 23750 3924 23756 3936
rect 23446 3896 23756 3924
rect 21637 3887 21695 3893
rect 23750 3884 23756 3896
rect 23808 3924 23814 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23808 3896 23857 3924
rect 23808 3884 23814 3896
rect 23845 3893 23857 3896
rect 23891 3924 23903 3927
rect 24228 3924 24256 3955
rect 24762 3952 24768 3964
rect 24820 3952 24826 4004
rect 23891 3896 24256 3924
rect 23891 3893 23903 3896
rect 23845 3887 23903 3893
rect 24670 3884 24676 3936
rect 24728 3924 24734 3936
rect 25731 3927 25789 3933
rect 25731 3924 25743 3927
rect 24728 3896 25743 3924
rect 24728 3884 24734 3896
rect 25731 3893 25743 3896
rect 25777 3893 25789 3927
rect 25731 3887 25789 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 2406 3680 2412 3732
rect 2464 3720 2470 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 2464 3692 3433 3720
rect 2464 3680 2470 3692
rect 14 3612 20 3664
rect 72 3652 78 3664
rect 1578 3652 1584 3664
rect 72 3624 1584 3652
rect 72 3612 78 3624
rect 1578 3612 1584 3624
rect 1636 3612 1642 3664
rect 2516 3661 2544 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 6546 3720 6552 3732
rect 5132 3692 6552 3720
rect 5132 3680 5138 3692
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 9122 3720 9128 3732
rect 7760 3692 8892 3720
rect 9083 3692 9128 3720
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3621 2559 3655
rect 2501 3615 2559 3621
rect 2593 3655 2651 3661
rect 2593 3621 2605 3655
rect 2639 3652 2651 3655
rect 2682 3652 2688 3664
rect 2639 3624 2688 3652
rect 2639 3621 2651 3624
rect 2593 3615 2651 3621
rect 2682 3612 2688 3624
rect 2740 3612 2746 3664
rect 3142 3652 3148 3664
rect 3103 3624 3148 3652
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 4154 3652 4160 3664
rect 3927 3624 4160 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 4154 3612 4160 3624
rect 4212 3612 4218 3664
rect 4258 3655 4316 3661
rect 4258 3621 4270 3655
rect 4304 3652 4316 3655
rect 4430 3652 4436 3664
rect 4304 3624 4436 3652
rect 4304 3621 4316 3624
rect 4258 3615 4316 3621
rect 4430 3612 4436 3624
rect 4488 3652 4494 3664
rect 5092 3652 5120 3680
rect 4488 3624 5120 3652
rect 5991 3655 6049 3661
rect 4488 3612 4494 3624
rect 5991 3621 6003 3655
rect 6037 3652 6049 3655
rect 6362 3652 6368 3664
rect 6037 3624 6368 3652
rect 6037 3621 6049 3624
rect 5991 3615 6049 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 5534 3544 5540 3596
rect 5592 3584 5598 3596
rect 5629 3587 5687 3593
rect 5629 3584 5641 3587
rect 5592 3556 5641 3584
rect 5592 3544 5598 3556
rect 5629 3553 5641 3556
rect 5675 3584 5687 3587
rect 7760 3584 7788 3692
rect 8202 3652 8208 3664
rect 8163 3624 8208 3652
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 8754 3652 8760 3664
rect 8715 3624 8760 3652
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 5675 3556 7788 3584
rect 5675 3553 5687 3556
rect 5629 3547 5687 3553
rect 1578 3476 1584 3528
rect 1636 3516 1642 3528
rect 6822 3516 6828 3528
rect 1636 3488 6828 3516
rect 1636 3476 1642 3488
rect 6822 3476 6828 3488
rect 6880 3476 6886 3528
rect 7558 3516 7564 3528
rect 7471 3488 7564 3516
rect 7558 3476 7564 3488
rect 7616 3516 7622 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7616 3488 8125 3516
rect 7616 3476 7622 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8864 3516 8892 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9306 3680 9312 3732
rect 9364 3720 9370 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9364 3692 9413 3720
rect 9364 3680 9370 3692
rect 9401 3689 9413 3692
rect 9447 3720 9459 3723
rect 9447 3692 9812 3720
rect 9447 3689 9459 3692
rect 9401 3683 9459 3689
rect 9784 3661 9812 3692
rect 10870 3680 10876 3732
rect 10928 3720 10934 3732
rect 11054 3720 11060 3732
rect 10928 3692 11060 3720
rect 10928 3680 10934 3692
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12437 3723 12495 3729
rect 12437 3720 12449 3723
rect 12400 3692 12449 3720
rect 12400 3680 12406 3692
rect 12437 3689 12449 3692
rect 12483 3689 12495 3723
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 12437 3683 12495 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 15746 3720 15752 3732
rect 13872 3692 13917 3720
rect 15707 3692 15752 3720
rect 13872 3680 13878 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 19242 3680 19248 3732
rect 19300 3720 19306 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19300 3692 19901 3720
rect 19300 3680 19306 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 19889 3683 19947 3689
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 9769 3655 9827 3661
rect 9769 3621 9781 3655
rect 9815 3621 9827 3655
rect 9769 3615 9827 3621
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 10413 3655 10471 3661
rect 9916 3624 9961 3652
rect 9916 3612 9922 3624
rect 10413 3621 10425 3655
rect 10459 3652 10471 3655
rect 10778 3652 10784 3664
rect 10459 3624 10784 3652
rect 10459 3621 10471 3624
rect 10413 3615 10471 3621
rect 10778 3612 10784 3624
rect 10836 3612 10842 3664
rect 14461 3655 14519 3661
rect 14461 3621 14473 3655
rect 14507 3652 14519 3655
rect 15654 3652 15660 3664
rect 14507 3624 15660 3652
rect 14507 3621 14519 3624
rect 14461 3615 14519 3621
rect 15654 3612 15660 3624
rect 15712 3612 15718 3664
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 21726 3652 21732 3664
rect 18196 3624 19380 3652
rect 21687 3624 21732 3652
rect 18196 3612 18202 3624
rect 10597 3587 10655 3593
rect 10597 3553 10609 3587
rect 10643 3584 10655 3587
rect 11054 3584 11060 3596
rect 10643 3556 11060 3584
rect 10643 3553 10655 3556
rect 10597 3547 10655 3553
rect 11054 3544 11060 3556
rect 11112 3584 11118 3596
rect 11241 3587 11299 3593
rect 11241 3584 11253 3587
rect 11112 3556 11253 3584
rect 11112 3544 11118 3556
rect 11241 3553 11253 3556
rect 11287 3553 11299 3587
rect 11241 3547 11299 3553
rect 11330 3544 11336 3596
rect 11388 3584 11394 3596
rect 11698 3584 11704 3596
rect 11388 3556 11704 3584
rect 11388 3544 11394 3556
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 12802 3584 12808 3596
rect 12763 3556 12808 3584
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13354 3584 13360 3596
rect 13127 3556 13360 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13354 3544 13360 3556
rect 13412 3544 13418 3596
rect 14274 3544 14280 3596
rect 14332 3584 14338 3596
rect 15289 3587 15347 3593
rect 15289 3584 15301 3587
rect 14332 3556 15301 3584
rect 14332 3544 14338 3556
rect 15289 3553 15301 3556
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 15565 3587 15623 3593
rect 15565 3553 15577 3587
rect 15611 3553 15623 3587
rect 15565 3547 15623 3553
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 8864 3488 11805 3516
rect 8113 3479 8171 3485
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 15580 3516 15608 3547
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16945 3587 17003 3593
rect 16945 3584 16957 3587
rect 16172 3556 16957 3584
rect 16172 3544 16178 3556
rect 16945 3553 16957 3556
rect 16991 3584 17003 3587
rect 17034 3584 17040 3596
rect 16991 3556 17040 3584
rect 16991 3553 17003 3556
rect 16945 3547 17003 3553
rect 17034 3544 17040 3556
rect 17092 3544 17098 3596
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 17497 3587 17555 3593
rect 17497 3584 17509 3587
rect 17184 3556 17509 3584
rect 17184 3544 17190 3556
rect 17497 3553 17509 3556
rect 17543 3584 17555 3587
rect 17678 3584 17684 3596
rect 17543 3556 17684 3584
rect 17543 3553 17555 3556
rect 17497 3547 17555 3553
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3584 17923 3587
rect 17954 3584 17960 3596
rect 17911 3556 17960 3584
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 11793 3479 11851 3485
rect 14844 3488 15608 3516
rect 16577 3519 16635 3525
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 4706 3448 4712 3460
rect 1719 3420 4153 3448
rect 4667 3420 4712 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 2406 3380 2412 3392
rect 2363 3352 2412 3380
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 2406 3340 2412 3352
rect 2464 3340 2470 3392
rect 4125 3380 4153 3420
rect 4706 3408 4712 3420
rect 4764 3448 4770 3460
rect 5169 3451 5227 3457
rect 5169 3448 5181 3451
rect 4764 3420 5181 3448
rect 4764 3408 4770 3420
rect 5169 3417 5181 3420
rect 5215 3448 5227 3451
rect 5258 3448 5264 3460
rect 5215 3420 5264 3448
rect 5215 3417 5227 3420
rect 5169 3411 5227 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 7834 3448 7840 3460
rect 7795 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 10134 3448 10140 3460
rect 7984 3420 10140 3448
rect 7984 3408 7990 3420
rect 10134 3408 10140 3420
rect 10192 3448 10198 3460
rect 10689 3451 10747 3457
rect 10689 3448 10701 3451
rect 10192 3420 10701 3448
rect 10192 3408 10198 3420
rect 10689 3417 10701 3420
rect 10735 3417 10747 3451
rect 10689 3411 10747 3417
rect 12710 3408 12716 3460
rect 12768 3448 12774 3460
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12768 3420 12909 3448
rect 12768 3408 12774 3420
rect 12897 3417 12909 3420
rect 12943 3448 12955 3451
rect 13722 3448 13728 3460
rect 12943 3420 13728 3448
rect 12943 3417 12955 3420
rect 12897 3411 12955 3417
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 14844 3392 14872 3488
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 17880 3516 17908 3547
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3584 18291 3587
rect 18782 3584 18788 3596
rect 18279 3556 18788 3584
rect 18279 3553 18291 3556
rect 18233 3547 18291 3553
rect 16623 3488 17908 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 15378 3448 15384 3460
rect 15291 3420 15384 3448
rect 15378 3408 15384 3420
rect 15436 3448 15442 3460
rect 15930 3448 15936 3460
rect 15436 3420 15936 3448
rect 15436 3408 15442 3420
rect 15930 3408 15936 3420
rect 15988 3408 15994 3460
rect 17402 3408 17408 3460
rect 17460 3448 17466 3460
rect 18248 3448 18276 3547
rect 18782 3544 18788 3556
rect 18840 3544 18846 3596
rect 19352 3593 19380 3624
rect 21726 3612 21732 3624
rect 21784 3612 21790 3664
rect 21818 3612 21824 3664
rect 21876 3652 21882 3664
rect 21876 3624 21921 3652
rect 21876 3612 21882 3624
rect 22094 3612 22100 3664
rect 22152 3652 22158 3664
rect 22830 3652 22836 3664
rect 22152 3624 22836 3652
rect 22152 3612 22158 3624
rect 22830 3612 22836 3624
rect 22888 3612 22894 3664
rect 24118 3652 24124 3664
rect 24079 3624 24124 3652
rect 24118 3612 24124 3624
rect 24176 3612 24182 3664
rect 24673 3655 24731 3661
rect 24673 3621 24685 3655
rect 24719 3652 24731 3655
rect 24762 3652 24768 3664
rect 24719 3624 24768 3652
rect 24719 3621 24731 3624
rect 24673 3615 24731 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 19337 3587 19395 3593
rect 19337 3553 19349 3587
rect 19383 3584 19395 3587
rect 21453 3587 21511 3593
rect 21453 3584 21465 3587
rect 19383 3556 21465 3584
rect 19383 3553 19395 3556
rect 19337 3547 19395 3553
rect 21453 3553 21465 3556
rect 21499 3553 21511 3587
rect 21453 3547 21511 3553
rect 22002 3516 22008 3528
rect 21963 3488 22008 3516
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 23198 3476 23204 3528
rect 23256 3516 23262 3528
rect 24029 3519 24087 3525
rect 24029 3516 24041 3519
rect 23256 3488 24041 3516
rect 23256 3476 23262 3488
rect 24029 3485 24041 3488
rect 24075 3485 24087 3519
rect 24029 3479 24087 3485
rect 18414 3448 18420 3460
rect 17460 3420 18276 3448
rect 18375 3420 18420 3448
rect 17460 3408 17466 3420
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 19521 3451 19579 3457
rect 19521 3417 19533 3451
rect 19567 3448 19579 3451
rect 20530 3448 20536 3460
rect 19567 3420 20536 3448
rect 19567 3417 19579 3420
rect 19521 3411 19579 3417
rect 20530 3408 20536 3420
rect 20588 3408 20594 3460
rect 7650 3380 7656 3392
rect 4125 3352 7656 3380
rect 7650 3340 7656 3352
rect 7708 3380 7714 3392
rect 10597 3383 10655 3389
rect 10597 3380 10609 3383
rect 7708 3352 10609 3380
rect 7708 3340 7714 3352
rect 10597 3349 10609 3352
rect 10643 3349 10655 3383
rect 14826 3380 14832 3392
rect 14787 3352 14832 3380
rect 10597 3343 10655 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 18782 3380 18788 3392
rect 18743 3352 18788 3380
rect 18782 3340 18788 3352
rect 18840 3380 18846 3392
rect 19153 3383 19211 3389
rect 19153 3380 19165 3383
rect 18840 3352 19165 3380
rect 18840 3340 18846 3352
rect 19153 3349 19165 3352
rect 19199 3380 19211 3383
rect 19426 3380 19432 3392
rect 19199 3352 19432 3380
rect 19199 3349 19211 3352
rect 19153 3343 19211 3349
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 20438 3380 20444 3392
rect 20399 3352 20444 3380
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 23750 3380 23756 3392
rect 23711 3352 23756 3380
rect 23750 3340 23756 3352
rect 23808 3340 23814 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1581 3179 1639 3185
rect 1581 3176 1593 3179
rect 1452 3148 1593 3176
rect 1452 3136 1458 3148
rect 1581 3145 1593 3148
rect 1627 3145 1639 3179
rect 1581 3139 1639 3145
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 3237 3179 3295 3185
rect 3237 3176 3249 3179
rect 2740 3148 3249 3176
rect 2740 3136 2746 3148
rect 3237 3145 3249 3148
rect 3283 3145 3295 3179
rect 3602 3176 3608 3188
rect 3563 3148 3608 3176
rect 3237 3139 3295 3145
rect 2130 3108 2136 3120
rect 2091 3080 2136 3108
rect 2130 3068 2136 3080
rect 2188 3068 2194 3120
rect 3252 3108 3280 3139
rect 3602 3136 3608 3148
rect 3660 3136 3666 3188
rect 5074 3176 5080 3188
rect 5035 3148 5080 3176
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6549 3179 6607 3185
rect 6549 3176 6561 3179
rect 6512 3148 6561 3176
rect 6512 3136 6518 3148
rect 6549 3145 6561 3148
rect 6595 3145 6607 3179
rect 6549 3139 6607 3145
rect 6963 3179 7021 3185
rect 6963 3145 6975 3179
rect 7009 3176 7021 3179
rect 7558 3176 7564 3188
rect 7009 3148 7564 3176
rect 7009 3145 7021 3148
rect 6963 3139 7021 3145
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 7837 3179 7895 3185
rect 7837 3145 7849 3179
rect 7883 3176 7895 3179
rect 8202 3176 8208 3188
rect 7883 3148 8208 3176
rect 7883 3145 7895 3148
rect 7837 3139 7895 3145
rect 8202 3136 8208 3148
rect 8260 3176 8266 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 8260 3148 9229 3176
rect 8260 3136 8266 3148
rect 9217 3145 9229 3148
rect 9263 3176 9275 3179
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 9263 3148 9505 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9493 3145 9505 3148
rect 9539 3176 9551 3179
rect 9858 3176 9864 3188
rect 9539 3148 9864 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11112 3148 11253 3176
rect 11112 3136 11118 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13412 3148 13829 3176
rect 13412 3136 13418 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 14182 3176 14188 3188
rect 14143 3148 14188 3176
rect 13817 3139 13875 3145
rect 14182 3136 14188 3148
rect 14240 3176 14246 3188
rect 21358 3176 21364 3188
rect 14240 3148 14872 3176
rect 21319 3148 21364 3176
rect 14240 3136 14246 3148
rect 4709 3111 4767 3117
rect 4709 3108 4721 3111
rect 3252 3080 4721 3108
rect 4709 3077 4721 3080
rect 4755 3077 4767 3111
rect 5534 3108 5540 3120
rect 5495 3080 5540 3108
rect 4709 3071 4767 3077
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 6273 3111 6331 3117
rect 6273 3077 6285 3111
rect 6319 3108 6331 3111
rect 6362 3108 6368 3120
rect 6319 3080 6368 3108
rect 6319 3077 6331 3080
rect 6273 3071 6331 3077
rect 6362 3068 6368 3080
rect 6420 3108 6426 3120
rect 7742 3108 7748 3120
rect 6420 3080 7748 3108
rect 6420 3068 6426 3080
rect 7742 3068 7748 3080
rect 7800 3108 7806 3120
rect 8113 3111 8171 3117
rect 8113 3108 8125 3111
rect 7800 3080 8125 3108
rect 7800 3068 7806 3080
rect 8113 3077 8125 3080
rect 8159 3077 8171 3111
rect 11790 3108 11796 3120
rect 11751 3080 11796 3108
rect 8113 3071 8171 3077
rect 2148 3040 2176 3068
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2148 3012 2329 3040
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3142 3040 3148 3052
rect 3007 3012 3148 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 6730 3040 6736 3052
rect 4126 3012 6736 3040
rect 3786 2972 3792 2984
rect 3747 2944 3792 2972
rect 3786 2932 3792 2944
rect 3844 2972 3850 2984
rect 4126 2972 4154 3012
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 3844 2944 4154 2972
rect 5721 2975 5779 2981
rect 3844 2932 3850 2944
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6454 2972 6460 2984
rect 5767 2944 6460 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6860 2975 6918 2981
rect 6860 2941 6872 2975
rect 6906 2941 6918 2975
rect 6860 2935 6918 2941
rect 2406 2904 2412 2916
rect 2319 2876 2412 2904
rect 2406 2864 2412 2876
rect 2464 2904 2470 2916
rect 2464 2876 3464 2904
rect 2464 2864 2470 2876
rect 3436 2848 3464 2876
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 4110 2907 4168 2913
rect 4110 2904 4122 2907
rect 3660 2876 4122 2904
rect 3660 2864 3666 2876
rect 4110 2873 4122 2876
rect 4156 2873 4168 2907
rect 4110 2867 4168 2873
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 6875 2904 6903 2935
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 5224 2876 7297 2904
rect 5224 2864 5230 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 8128 2904 8156 3071
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 14274 3068 14280 3120
rect 14332 3108 14338 3120
rect 14844 3117 14872 3148
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 22005 3179 22063 3185
rect 22005 3176 22017 3179
rect 21784 3148 22017 3176
rect 21784 3136 21790 3148
rect 22005 3145 22017 3148
rect 22051 3145 22063 3179
rect 22005 3139 22063 3145
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 23256 3148 23397 3176
rect 23256 3136 23262 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 14553 3111 14611 3117
rect 14553 3108 14565 3111
rect 14332 3080 14565 3108
rect 14332 3068 14338 3080
rect 14553 3077 14565 3080
rect 14599 3077 14611 3111
rect 14553 3071 14611 3077
rect 14829 3111 14887 3117
rect 14829 3077 14841 3111
rect 14875 3077 14887 3111
rect 14829 3071 14887 3077
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3040 8355 3043
rect 9122 3040 9128 3052
rect 8343 3012 9128 3040
rect 8343 3009 8355 3012
rect 8297 3003 8355 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 10134 3040 10140 3052
rect 10095 3012 10140 3040
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10778 3040 10784 3052
rect 10739 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11808 3040 11836 3068
rect 11808 3012 12940 3040
rect 12342 2932 12348 2984
rect 12400 2972 12406 2984
rect 12912 2981 12940 3012
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12400 2944 12449 2972
rect 12400 2932 12406 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2941 12955 2975
rect 14568 2972 14596 3071
rect 17034 3068 17040 3120
rect 17092 3108 17098 3120
rect 19889 3111 19947 3117
rect 19889 3108 19901 3111
rect 17092 3080 19901 3108
rect 17092 3068 17098 3080
rect 15470 3040 15476 3052
rect 15431 3012 15476 3040
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 16574 3040 16580 3052
rect 15620 3012 16580 3040
rect 15620 3000 15626 3012
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 17770 3040 17776 3052
rect 17731 3012 17776 3040
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 14737 2975 14795 2981
rect 14737 2972 14749 2975
rect 14568 2944 14749 2972
rect 12897 2935 12955 2941
rect 14737 2941 14749 2944
rect 14783 2941 14795 2975
rect 15010 2972 15016 2984
rect 14971 2944 15016 2972
rect 14737 2935 14795 2941
rect 8618 2907 8676 2913
rect 8618 2904 8630 2907
rect 8128 2876 8630 2904
rect 7285 2867 7343 2873
rect 8618 2873 8630 2876
rect 8664 2873 8676 2907
rect 8618 2867 8676 2873
rect 9766 2864 9772 2916
rect 9824 2904 9830 2916
rect 9861 2907 9919 2913
rect 9861 2904 9873 2907
rect 9824 2876 9873 2904
rect 9824 2864 9830 2876
rect 9861 2873 9873 2876
rect 9907 2904 9919 2907
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 9907 2876 10241 2904
rect 9907 2873 9919 2876
rect 9861 2867 9919 2873
rect 10229 2873 10241 2876
rect 10275 2873 10287 2907
rect 12161 2907 12219 2913
rect 12161 2904 12173 2907
rect 10229 2867 10287 2873
rect 10428 2876 12173 2904
rect 3418 2796 3424 2848
rect 3476 2836 3482 2848
rect 3970 2836 3976 2848
rect 3476 2808 3976 2836
rect 3476 2796 3482 2808
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2836 5963 2839
rect 10428 2836 10456 2876
rect 12161 2873 12173 2876
rect 12207 2904 12219 2907
rect 12802 2904 12808 2916
rect 12207 2876 12808 2904
rect 12207 2873 12219 2876
rect 12161 2867 12219 2873
rect 12802 2864 12808 2876
rect 12860 2864 12866 2916
rect 14752 2904 14780 2935
rect 15010 2932 15016 2944
rect 15068 2932 15074 2984
rect 18432 2981 18460 3080
rect 19889 3077 19901 3080
rect 19935 3077 19947 3111
rect 19889 3071 19947 3077
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 20438 3040 20444 3052
rect 19659 3012 20444 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 21729 3043 21787 3049
rect 21729 3009 21741 3043
rect 21775 3040 21787 3043
rect 21818 3040 21824 3052
rect 21775 3012 21824 3040
rect 21775 3009 21787 3012
rect 21729 3003 21787 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22612 3012 24072 3040
rect 22612 3000 22618 3012
rect 18417 2975 18475 2981
rect 18417 2941 18429 2975
rect 18463 2941 18475 2975
rect 18417 2935 18475 2941
rect 18601 2975 18659 2981
rect 18601 2941 18613 2975
rect 18647 2972 18659 2975
rect 18782 2972 18788 2984
rect 18647 2944 18788 2972
rect 18647 2941 18659 2944
rect 18601 2935 18659 2941
rect 16117 2907 16175 2913
rect 16117 2904 16129 2907
rect 14752 2876 16129 2904
rect 16117 2873 16129 2876
rect 16163 2873 16175 2907
rect 16117 2867 16175 2873
rect 16298 2864 16304 2916
rect 16356 2904 16362 2916
rect 16474 2907 16532 2913
rect 16474 2904 16486 2907
rect 16356 2876 16486 2904
rect 16356 2864 16362 2876
rect 16474 2873 16486 2876
rect 16520 2873 16532 2907
rect 16474 2867 16532 2873
rect 16577 2907 16635 2913
rect 16577 2873 16589 2907
rect 16623 2904 16635 2907
rect 16850 2904 16856 2916
rect 16623 2876 16856 2904
rect 16623 2873 16635 2876
rect 16577 2867 16635 2873
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 17126 2904 17132 2916
rect 17087 2876 17132 2904
rect 17126 2864 17132 2876
rect 17184 2864 17190 2916
rect 17678 2864 17684 2916
rect 17736 2904 17742 2916
rect 18616 2904 18644 2935
rect 18782 2932 18788 2944
rect 18840 2932 18846 2984
rect 18966 2972 18972 2984
rect 18927 2944 18972 2972
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 18874 2904 18880 2916
rect 17736 2876 18644 2904
rect 18702 2876 18880 2904
rect 17736 2864 17742 2876
rect 12526 2836 12532 2848
rect 5951 2808 10456 2836
rect 12487 2808 12532 2836
rect 5951 2805 5963 2808
rect 5905 2799 5963 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 13722 2836 13728 2848
rect 13587 2808 13728 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 15841 2839 15899 2845
rect 15841 2805 15853 2839
rect 15887 2836 15899 2839
rect 15930 2836 15936 2848
rect 15887 2808 15936 2836
rect 15887 2805 15899 2808
rect 15841 2799 15899 2805
rect 15930 2796 15936 2808
rect 15988 2796 15994 2848
rect 17402 2836 17408 2848
rect 17363 2808 17408 2836
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17770 2796 17776 2848
rect 17828 2836 17834 2848
rect 18702 2836 18730 2876
rect 18874 2864 18880 2876
rect 18932 2904 18938 2916
rect 19352 2904 19380 2935
rect 20990 2932 20996 2984
rect 21048 2972 21054 2984
rect 22189 2975 22247 2981
rect 22189 2972 22201 2975
rect 21048 2944 22201 2972
rect 21048 2932 21054 2944
rect 22189 2941 22201 2944
rect 22235 2972 22247 2975
rect 22741 2975 22799 2981
rect 22741 2972 22753 2975
rect 22235 2944 22753 2972
rect 22235 2941 22247 2944
rect 22189 2935 22247 2941
rect 22741 2941 22753 2944
rect 22787 2941 22799 2975
rect 23750 2972 23756 2984
rect 23711 2944 23756 2972
rect 22741 2935 22799 2941
rect 23750 2932 23756 2944
rect 23808 2932 23814 2984
rect 24044 2972 24072 3012
rect 24118 3000 24124 3052
rect 24176 3040 24182 3052
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 24176 3012 24409 3040
rect 24176 3000 24182 3012
rect 24397 3009 24409 3012
rect 24443 3040 24455 3043
rect 24673 3043 24731 3049
rect 24673 3040 24685 3043
rect 24443 3012 24685 3040
rect 24443 3009 24455 3012
rect 24397 3003 24455 3009
rect 24673 3009 24685 3012
rect 24719 3009 24731 3043
rect 24673 3003 24731 3009
rect 25225 2975 25283 2981
rect 25225 2972 25237 2975
rect 24044 2944 25237 2972
rect 25225 2941 25237 2944
rect 25271 2972 25283 2975
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25271 2944 25789 2972
rect 25271 2941 25283 2944
rect 25225 2935 25283 2941
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 20714 2904 20720 2916
rect 18932 2876 19380 2904
rect 20272 2876 20720 2904
rect 18932 2864 18938 2876
rect 17828 2808 18730 2836
rect 17828 2796 17834 2808
rect 18782 2796 18788 2848
rect 18840 2836 18846 2848
rect 20272 2845 20300 2876
rect 20714 2864 20720 2876
rect 20772 2913 20778 2916
rect 20772 2907 20820 2913
rect 20772 2873 20774 2907
rect 20808 2873 20820 2907
rect 20772 2867 20820 2873
rect 20772 2864 20778 2867
rect 20257 2839 20315 2845
rect 20257 2836 20269 2839
rect 18840 2808 20269 2836
rect 18840 2796 18846 2808
rect 20257 2805 20269 2808
rect 20303 2805 20315 2839
rect 20257 2799 20315 2805
rect 21726 2796 21732 2848
rect 21784 2836 21790 2848
rect 22373 2839 22431 2845
rect 22373 2836 22385 2839
rect 21784 2808 22385 2836
rect 21784 2796 21790 2808
rect 22373 2805 22385 2808
rect 22419 2805 22431 2839
rect 22373 2799 22431 2805
rect 25409 2839 25467 2845
rect 25409 2805 25421 2839
rect 25455 2836 25467 2839
rect 27522 2836 27528 2848
rect 25455 2808 27528 2836
rect 25455 2805 25467 2808
rect 25409 2799 25467 2805
rect 27522 2796 27528 2808
rect 27580 2796 27586 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 3418 2632 3424 2644
rect 2372 2604 2865 2632
rect 3379 2604 3424 2632
rect 2372 2592 2378 2604
rect 2225 2567 2283 2573
rect 2225 2533 2237 2567
rect 2271 2564 2283 2567
rect 2593 2567 2651 2573
rect 2593 2564 2605 2567
rect 2271 2536 2605 2564
rect 2271 2533 2283 2536
rect 2225 2527 2283 2533
rect 2593 2533 2605 2536
rect 2639 2564 2651 2567
rect 2682 2564 2688 2576
rect 2639 2536 2688 2564
rect 2639 2533 2651 2536
rect 2593 2527 2651 2533
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 2837 2564 2865 2604
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4154 2632 4160 2644
rect 3896 2604 4160 2632
rect 3896 2564 3924 2604
rect 4154 2592 4160 2604
rect 4212 2592 4218 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5077 2635 5135 2641
rect 5077 2632 5089 2635
rect 5040 2604 5089 2632
rect 5040 2592 5046 2604
rect 5077 2601 5089 2604
rect 5123 2601 5135 2635
rect 5077 2595 5135 2601
rect 7055 2635 7113 2641
rect 7055 2601 7067 2635
rect 7101 2632 7113 2635
rect 7834 2632 7840 2644
rect 7101 2604 7840 2632
rect 7101 2601 7113 2604
rect 7055 2595 7113 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 9217 2635 9275 2641
rect 9217 2632 9229 2635
rect 7944 2604 9229 2632
rect 2837 2536 3924 2564
rect 3970 2524 3976 2576
rect 4028 2564 4034 2576
rect 4249 2567 4307 2573
rect 4249 2564 4261 2567
rect 4028 2536 4261 2564
rect 4028 2524 4034 2536
rect 4249 2533 4261 2536
rect 4295 2533 4307 2567
rect 7742 2564 7748 2576
rect 7703 2536 7748 2564
rect 4249 2527 4307 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1946 2496 1952 2508
rect 1443 2468 1952 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5859 2468 6285 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6273 2459 6331 2465
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7282 2496 7288 2508
rect 7030 2468 7288 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2428 2559 2431
rect 3878 2428 3884 2440
rect 2547 2400 3884 2428
rect 2547 2397 2559 2400
rect 2501 2391 2559 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4154 2388 4160 2440
rect 4212 2428 4218 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 4212 2400 5457 2428
rect 4212 2388 4218 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 4706 2360 4712 2372
rect 3099 2332 4712 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 4706 2320 4712 2332
rect 4764 2320 4770 2372
rect 6288 2360 6316 2459
rect 7282 2456 7288 2468
rect 7340 2496 7346 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7340 2468 7389 2496
rect 7340 2456 7346 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 7760 2428 7788 2524
rect 7944 2505 7972 2604
rect 9217 2601 9229 2604
rect 9263 2632 9275 2635
rect 12526 2632 12532 2644
rect 9263 2604 12532 2632
rect 9263 2601 9275 2604
rect 9217 2595 9275 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 15010 2592 15016 2644
rect 15068 2632 15074 2644
rect 16117 2635 16175 2641
rect 16117 2632 16129 2635
rect 15068 2604 16129 2632
rect 15068 2592 15074 2604
rect 16117 2601 16129 2604
rect 16163 2601 16175 2635
rect 16117 2595 16175 2601
rect 16577 2635 16635 2641
rect 16577 2601 16589 2635
rect 16623 2632 16635 2635
rect 16666 2632 16672 2644
rect 16623 2604 16672 2632
rect 16623 2601 16635 2604
rect 16577 2595 16635 2601
rect 16666 2592 16672 2604
rect 16724 2632 16730 2644
rect 17678 2632 17684 2644
rect 16724 2604 16896 2632
rect 17639 2604 17684 2632
rect 16724 2592 16730 2604
rect 8250 2567 8308 2573
rect 8250 2564 8262 2567
rect 8036 2536 8262 2564
rect 7929 2499 7987 2505
rect 7929 2465 7941 2499
rect 7975 2465 7987 2499
rect 7929 2459 7987 2465
rect 8036 2428 8064 2536
rect 8250 2533 8262 2536
rect 8296 2533 8308 2567
rect 8250 2527 8308 2533
rect 9858 2524 9864 2576
rect 9916 2564 9922 2576
rect 10045 2567 10103 2573
rect 10045 2564 10057 2567
rect 9916 2536 10057 2564
rect 9916 2524 9922 2536
rect 10045 2533 10057 2536
rect 10091 2564 10103 2567
rect 10413 2567 10471 2573
rect 10413 2564 10425 2567
rect 10091 2536 10425 2564
rect 10091 2533 10103 2536
rect 10045 2527 10103 2533
rect 10413 2533 10425 2536
rect 10459 2533 10471 2567
rect 10962 2564 10968 2576
rect 10923 2536 10968 2564
rect 10413 2527 10471 2533
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 11330 2564 11336 2576
rect 11291 2536 11336 2564
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 12066 2524 12072 2576
rect 12124 2564 12130 2576
rect 12621 2567 12679 2573
rect 12621 2564 12633 2567
rect 12124 2536 12633 2564
rect 12124 2524 12130 2536
rect 12621 2533 12633 2536
rect 12667 2533 12679 2567
rect 12621 2527 12679 2533
rect 13817 2567 13875 2573
rect 13817 2533 13829 2567
rect 13863 2564 13875 2567
rect 14366 2564 14372 2576
rect 13863 2536 14372 2564
rect 13863 2533 13875 2536
rect 13817 2527 13875 2533
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 9766 2496 9772 2508
rect 8895 2468 9772 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 14292 2505 14320 2536
rect 14366 2524 14372 2536
rect 14424 2524 14430 2576
rect 15194 2564 15200 2576
rect 15155 2536 15200 2564
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 16868 2573 16896 2604
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 18141 2635 18199 2641
rect 18141 2601 18153 2635
rect 18187 2632 18199 2635
rect 18690 2632 18696 2644
rect 18187 2604 18696 2632
rect 18187 2601 18199 2604
rect 18141 2595 18199 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 18966 2592 18972 2644
rect 19024 2632 19030 2644
rect 19521 2635 19579 2641
rect 19521 2632 19533 2635
rect 19024 2604 19533 2632
rect 19024 2592 19030 2604
rect 19521 2601 19533 2604
rect 19567 2601 19579 2635
rect 19521 2595 19579 2601
rect 20622 2592 20628 2644
rect 20680 2632 20686 2644
rect 22646 2632 22652 2644
rect 20680 2604 21956 2632
rect 22607 2604 22652 2632
rect 20680 2592 20686 2604
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 20993 2567 21051 2573
rect 20993 2533 21005 2567
rect 21039 2564 21051 2567
rect 21358 2564 21364 2576
rect 21039 2536 21364 2564
rect 21039 2533 21051 2536
rect 20993 2527 21051 2533
rect 21358 2524 21364 2536
rect 21416 2524 21422 2576
rect 21928 2573 21956 2604
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 22830 2592 22836 2644
rect 22888 2632 22894 2644
rect 23753 2635 23811 2641
rect 23753 2632 23765 2635
rect 22888 2604 23765 2632
rect 22888 2592 22894 2604
rect 23753 2601 23765 2604
rect 23799 2632 23811 2635
rect 26142 2632 26148 2644
rect 23799 2604 24256 2632
rect 26103 2604 26148 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 21913 2567 21971 2573
rect 21913 2533 21925 2567
rect 21959 2564 21971 2567
rect 21959 2536 22600 2564
rect 21959 2533 21971 2536
rect 21913 2527 21971 2533
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12360 2468 12725 2496
rect 7760 2400 8064 2428
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 10318 2428 10324 2440
rect 9631 2400 10324 2428
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 11698 2360 11704 2372
rect 6288 2332 11704 2360
rect 11698 2320 11704 2332
rect 11756 2360 11762 2372
rect 12066 2360 12072 2372
rect 11756 2332 12072 2360
rect 11756 2320 11762 2332
rect 12066 2320 12072 2332
rect 12124 2360 12130 2372
rect 12360 2369 12388 2468
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 12713 2459 12771 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2465 14335 2499
rect 15212 2496 15240 2524
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15212 2468 15577 2496
rect 14277 2459 14335 2465
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18414 2496 18420 2508
rect 18371 2468 18420 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18414 2456 18420 2468
rect 18472 2496 18478 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 18472 2468 19901 2496
rect 18472 2456 18478 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20140 2499 20198 2505
rect 20140 2465 20152 2499
rect 20186 2496 20198 2499
rect 20622 2496 20628 2508
rect 20186 2468 20628 2496
rect 20186 2465 20198 2468
rect 20140 2459 20198 2465
rect 20622 2456 20628 2468
rect 20680 2456 20686 2508
rect 14182 2428 14188 2440
rect 14095 2400 14188 2428
rect 14182 2388 14188 2400
rect 14240 2428 14246 2440
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 14240 2400 16773 2428
rect 14240 2388 14246 2400
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 16761 2391 16819 2397
rect 17126 2388 17132 2400
rect 17184 2428 17190 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 17184 2400 21281 2428
rect 17184 2388 17190 2400
rect 21269 2397 21281 2400
rect 21315 2428 21327 2431
rect 22189 2431 22247 2437
rect 22189 2428 22201 2431
rect 21315 2400 22201 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 22189 2397 22201 2400
rect 22235 2397 22247 2431
rect 22572 2428 22600 2536
rect 22664 2496 22692 2592
rect 24228 2573 24256 2604
rect 26142 2592 26148 2604
rect 26200 2592 26206 2644
rect 23661 2567 23719 2573
rect 23661 2533 23673 2567
rect 23707 2564 23719 2567
rect 24121 2567 24179 2573
rect 24121 2564 24133 2567
rect 23707 2536 24133 2564
rect 23707 2533 23719 2536
rect 23661 2527 23719 2533
rect 24121 2533 24133 2536
rect 24167 2533 24179 2567
rect 24121 2527 24179 2533
rect 24213 2567 24271 2573
rect 24213 2533 24225 2567
rect 24259 2533 24271 2567
rect 24213 2527 24271 2533
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22664 2468 22845 2496
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 25660 2499 25718 2505
rect 25660 2465 25672 2499
rect 25706 2496 25718 2499
rect 26160 2496 26188 2592
rect 25706 2468 26188 2496
rect 25706 2465 25718 2468
rect 25660 2459 25718 2465
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 22572 2400 24072 2428
rect 22189 2391 22247 2397
rect 12345 2363 12403 2369
rect 12345 2360 12357 2363
rect 12124 2332 12357 2360
rect 12124 2320 12130 2332
rect 12345 2329 12357 2332
rect 12391 2329 12403 2363
rect 12345 2323 12403 2329
rect 14921 2363 14979 2369
rect 14921 2329 14933 2363
rect 14967 2360 14979 2363
rect 16298 2360 16304 2372
rect 14967 2332 16304 2360
rect 14967 2329 14979 2332
rect 14921 2323 14979 2329
rect 16298 2320 16304 2332
rect 16356 2320 16362 2372
rect 16850 2320 16856 2372
rect 16908 2360 16914 2372
rect 19245 2363 19303 2369
rect 19245 2360 19257 2363
rect 16908 2332 19257 2360
rect 16908 2320 16914 2332
rect 19245 2329 19257 2332
rect 19291 2329 19303 2363
rect 19245 2323 19303 2329
rect 23017 2363 23075 2369
rect 23017 2329 23029 2363
rect 23063 2360 23075 2363
rect 24044 2360 24072 2400
rect 24228 2400 24409 2428
rect 24228 2360 24256 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 26602 2360 26608 2372
rect 23063 2332 23980 2360
rect 24044 2332 24256 2360
rect 24596 2332 26608 2360
rect 23063 2329 23075 2332
rect 23017 2323 23075 2329
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4982 2292 4988 2304
rect 3936 2264 4988 2292
rect 3936 2252 3942 2264
rect 4982 2252 4988 2264
rect 5040 2252 5046 2304
rect 5994 2292 6000 2304
rect 5955 2264 6000 2292
rect 5994 2252 6000 2264
rect 6052 2252 6058 2304
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2292 14519 2295
rect 14734 2292 14740 2304
rect 14507 2264 14740 2292
rect 14507 2261 14519 2264
rect 14461 2255 14519 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15746 2292 15752 2304
rect 15707 2264 15752 2292
rect 15746 2252 15752 2264
rect 15804 2252 15810 2304
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 20211 2295 20269 2301
rect 20211 2292 20223 2295
rect 19392 2264 20223 2292
rect 19392 2252 19398 2264
rect 20211 2261 20223 2264
rect 20257 2261 20269 2295
rect 20622 2292 20628 2304
rect 20583 2264 20628 2292
rect 20211 2255 20269 2261
rect 20622 2252 20628 2264
rect 20680 2252 20686 2304
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 20864 2264 23397 2292
rect 20864 2252 20870 2264
rect 23385 2261 23397 2264
rect 23431 2292 23443 2295
rect 23661 2295 23719 2301
rect 23661 2292 23673 2295
rect 23431 2264 23673 2292
rect 23431 2261 23443 2264
rect 23385 2255 23443 2261
rect 23661 2261 23673 2264
rect 23707 2261 23719 2295
rect 23952 2292 23980 2332
rect 24596 2292 24624 2332
rect 26602 2320 26608 2332
rect 26660 2320 26666 2372
rect 23952 2264 24624 2292
rect 23661 2255 23719 2261
rect 24670 2252 24676 2304
rect 24728 2292 24734 2304
rect 25731 2295 25789 2301
rect 25731 2292 25743 2295
rect 24728 2264 25743 2292
rect 24728 2252 24734 2264
rect 25731 2261 25743 2264
rect 25777 2261 25789 2295
rect 25731 2255 25789 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 2590 2048 2596 2100
rect 2648 2088 2654 2100
rect 2958 2088 2964 2100
rect 2648 2060 2964 2088
rect 2648 2048 2654 2060
rect 2958 2048 2964 2060
rect 3016 2088 3022 2100
rect 7282 2088 7288 2100
rect 3016 2060 7288 2088
rect 3016 2048 3022 2060
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 19334 2088 19340 2100
rect 10744 2060 19340 2088
rect 10744 2048 10750 2060
rect 19334 2048 19340 2060
rect 19392 2048 19398 2100
rect 8478 76 8484 128
rect 8536 116 8542 128
rect 9122 116 9128 128
rect 8536 88 9128 116
rect 8536 76 8542 88
rect 9122 76 9128 88
rect 9180 76 9186 128
rect 15746 76 15752 128
rect 15804 116 15810 128
rect 19702 116 19708 128
rect 15804 88 19708 116
rect 15804 76 15810 88
rect 19702 76 19708 88
rect 19760 76 19766 128
<< via1 >>
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 1584 23851 1636 23860
rect 1584 23817 1593 23851
rect 1593 23817 1627 23851
rect 1627 23817 1636 23851
rect 1584 23808 1636 23817
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 23480 23604 23532 23656
rect 2136 23468 2188 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 24768 21675 24820 21684
rect 24768 21641 24777 21675
rect 24777 21641 24811 21675
rect 24811 21641 24820 21675
rect 24768 21632 24820 21641
rect 1124 21428 1176 21480
rect 24032 21428 24084 21480
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 1400 20383 1452 20392
rect 1400 20349 1444 20383
rect 1444 20349 1452 20383
rect 1400 20340 1452 20349
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1308 19864 1360 19916
rect 2228 19864 2280 19916
rect 1308 19660 1360 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2228 19499 2280 19508
rect 2228 19465 2237 19499
rect 2237 19465 2271 19499
rect 2271 19465 2280 19499
rect 2228 19456 2280 19465
rect 2044 19388 2096 19440
rect 1860 19295 1912 19304
rect 1860 19261 1869 19295
rect 1869 19261 1903 19295
rect 1903 19261 1912 19295
rect 1860 19252 1912 19261
rect 1952 19116 2004 19168
rect 3240 19116 3292 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 1216 18776 1268 18828
rect 2228 18776 2280 18828
rect 1768 18572 1820 18624
rect 2320 18572 2372 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1124 18300 1176 18352
rect 1400 18300 1452 18352
rect 940 18164 992 18216
rect 2228 18164 2280 18216
rect 296 18096 348 18148
rect 1216 18096 1268 18148
rect 4344 18139 4396 18148
rect 4344 18105 4353 18139
rect 4353 18105 4387 18139
rect 4387 18105 4396 18139
rect 4344 18096 4396 18105
rect 7288 18139 7340 18148
rect 7288 18105 7297 18139
rect 7297 18105 7331 18139
rect 7331 18105 7340 18139
rect 7288 18096 7340 18105
rect 1124 18028 1176 18080
rect 2780 18071 2832 18080
rect 2780 18037 2789 18071
rect 2789 18037 2823 18071
rect 2823 18037 2832 18071
rect 2780 18028 2832 18037
rect 3424 18028 3476 18080
rect 6828 18028 6880 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1584 17867 1636 17876
rect 1584 17833 1593 17867
rect 1593 17833 1627 17867
rect 1627 17833 1636 17867
rect 1584 17824 1636 17833
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 2320 17688 2372 17740
rect 3056 17688 3108 17740
rect 3976 17731 4028 17740
rect 3976 17697 3985 17731
rect 3985 17697 4019 17731
rect 4019 17697 4028 17731
rect 3976 17688 4028 17697
rect 5264 17688 5316 17740
rect 6736 17731 6788 17740
rect 6736 17697 6745 17731
rect 6745 17697 6779 17731
rect 6779 17697 6788 17731
rect 6736 17688 6788 17697
rect 13452 17731 13504 17740
rect 13452 17697 13461 17731
rect 13461 17697 13495 17731
rect 13495 17697 13504 17731
rect 13452 17688 13504 17697
rect 13912 17731 13964 17740
rect 13912 17697 13921 17731
rect 13921 17697 13955 17731
rect 13955 17697 13964 17731
rect 13912 17688 13964 17697
rect 15568 17731 15620 17740
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 24676 17688 24728 17740
rect 11612 17620 11664 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 2964 17484 3016 17536
rect 3792 17484 3844 17536
rect 5080 17484 5132 17536
rect 7196 17484 7248 17536
rect 15292 17484 15344 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 8668 17280 8720 17332
rect 10968 17280 11020 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 6368 17212 6420 17264
rect 8760 17212 8812 17264
rect 10876 17212 10928 17264
rect 112 17076 164 17128
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 4620 17144 4672 17196
rect 12992 17187 13044 17196
rect 3148 17008 3200 17060
rect 3976 17008 4028 17060
rect 3056 16940 3108 16992
rect 3700 16940 3752 16992
rect 4712 16940 4764 16992
rect 4804 16940 4856 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5356 16940 5408 16992
rect 9220 17076 9272 17128
rect 11796 17076 11848 17128
rect 11980 17076 12032 17128
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13820 17144 13872 17196
rect 15568 17187 15620 17196
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 6184 16940 6236 16992
rect 6736 16940 6788 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 9128 16940 9180 16992
rect 11060 16940 11112 16992
rect 14188 17076 14240 17128
rect 15660 17076 15712 17128
rect 15844 17008 15896 17060
rect 13912 16983 13964 16992
rect 13912 16949 13921 16983
rect 13921 16949 13955 16983
rect 13955 16949 13964 16983
rect 13912 16940 13964 16949
rect 16028 16940 16080 16992
rect 22928 16940 22980 16992
rect 24584 16983 24636 16992
rect 24584 16949 24593 16983
rect 24593 16949 24627 16983
rect 24627 16949 24636 16983
rect 24584 16940 24636 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1032 16736 1084 16788
rect 7748 16779 7800 16788
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 13728 16736 13780 16788
rect 24584 16736 24636 16788
rect 6184 16668 6236 16720
rect 1584 16600 1636 16652
rect 2596 16600 2648 16652
rect 4436 16600 4488 16652
rect 6276 16600 6328 16652
rect 7104 16600 7156 16652
rect 7840 16643 7892 16652
rect 7840 16609 7849 16643
rect 7849 16609 7883 16643
rect 7883 16609 7892 16643
rect 7840 16600 7892 16609
rect 6000 16464 6052 16516
rect 2504 16396 2556 16448
rect 3332 16396 3384 16448
rect 6092 16396 6144 16448
rect 6644 16396 6696 16448
rect 7656 16532 7708 16584
rect 8208 16532 8260 16584
rect 9772 16600 9824 16652
rect 12716 16600 12768 16652
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 13912 16600 13964 16652
rect 14280 16600 14332 16652
rect 15384 16600 15436 16652
rect 15476 16600 15528 16652
rect 16856 16643 16908 16652
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 23572 16600 23624 16652
rect 24768 16600 24820 16652
rect 10048 16532 10100 16584
rect 14556 16532 14608 16584
rect 20812 16532 20864 16584
rect 14188 16464 14240 16516
rect 16672 16464 16724 16516
rect 10876 16439 10928 16448
rect 10876 16405 10885 16439
rect 10885 16405 10919 16439
rect 10919 16405 10928 16439
rect 10876 16396 10928 16405
rect 12256 16439 12308 16448
rect 12256 16405 12265 16439
rect 12265 16405 12299 16439
rect 12299 16405 12308 16439
rect 12256 16396 12308 16405
rect 17040 16439 17092 16448
rect 17040 16405 17049 16439
rect 17049 16405 17083 16439
rect 17083 16405 17092 16439
rect 17040 16396 17092 16405
rect 18604 16396 18656 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 1492 16192 1544 16244
rect 2136 16192 2188 16244
rect 4160 16124 4212 16176
rect 11980 16192 12032 16244
rect 12072 16192 12124 16244
rect 15384 16192 15436 16244
rect 16120 16192 16172 16244
rect 16672 16235 16724 16244
rect 16672 16201 16681 16235
rect 16681 16201 16715 16235
rect 16715 16201 16724 16235
rect 16672 16192 16724 16201
rect 24768 16192 24820 16244
rect 25228 16235 25280 16244
rect 25228 16201 25237 16235
rect 25237 16201 25271 16235
rect 25271 16201 25280 16235
rect 25228 16192 25280 16201
rect 6276 16099 6328 16108
rect 6276 16065 6285 16099
rect 6285 16065 6319 16099
rect 6319 16065 6328 16099
rect 6276 16056 6328 16065
rect 1492 15920 1544 15972
rect 2688 15988 2740 16040
rect 4344 15988 4396 16040
rect 3976 15963 4028 15972
rect 3976 15929 3985 15963
rect 3985 15929 4019 15963
rect 4019 15929 4028 15963
rect 3976 15920 4028 15929
rect 7472 15988 7524 16040
rect 12716 16124 12768 16176
rect 17592 16124 17644 16176
rect 22008 16124 22060 16176
rect 23572 16124 23624 16176
rect 8208 15988 8260 16040
rect 12256 16056 12308 16108
rect 8392 15988 8444 16040
rect 9772 16031 9824 16040
rect 9772 15997 9781 16031
rect 9781 15997 9815 16031
rect 9815 15997 9824 16031
rect 9772 15988 9824 15997
rect 7840 15920 7892 15972
rect 8300 15920 8352 15972
rect 10876 15988 10928 16040
rect 11520 15963 11572 15972
rect 11520 15929 11529 15963
rect 11529 15929 11563 15963
rect 11563 15929 11572 15963
rect 11520 15920 11572 15929
rect 12624 15988 12676 16040
rect 12900 15920 12952 15972
rect 15200 16056 15252 16108
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 22744 16056 22796 16108
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 25228 15988 25280 16040
rect 18420 15920 18472 15972
rect 23112 15920 23164 15972
rect 2412 15852 2464 15904
rect 3884 15852 3936 15904
rect 4436 15895 4488 15904
rect 4436 15861 4445 15895
rect 4445 15861 4479 15895
rect 4479 15861 4488 15895
rect 4436 15852 4488 15861
rect 5540 15852 5592 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 8024 15852 8076 15904
rect 9312 15895 9364 15904
rect 9312 15861 9321 15895
rect 9321 15861 9355 15895
rect 9355 15861 9364 15895
rect 9312 15852 9364 15861
rect 10048 15852 10100 15904
rect 12440 15852 12492 15904
rect 13544 15852 13596 15904
rect 15476 15852 15528 15904
rect 16856 15852 16908 15904
rect 18144 15852 18196 15904
rect 21732 15852 21784 15904
rect 22468 15852 22520 15904
rect 24952 15852 25004 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 2044 15648 2096 15700
rect 20 15580 72 15632
rect 2688 15580 2740 15632
rect 7932 15648 7984 15700
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 2044 15555 2096 15564
rect 2044 15521 2053 15555
rect 2053 15521 2087 15555
rect 2087 15521 2096 15555
rect 2044 15512 2096 15521
rect 2872 15512 2924 15564
rect 4252 15512 4304 15564
rect 4896 15512 4948 15564
rect 6460 15512 6512 15564
rect 9772 15580 9824 15632
rect 14280 15623 14332 15632
rect 6644 15512 6696 15564
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 10968 15512 11020 15564
rect 14280 15589 14289 15623
rect 14289 15589 14323 15623
rect 14323 15589 14332 15623
rect 14280 15580 14332 15589
rect 18236 15580 18288 15632
rect 11704 15512 11756 15564
rect 12348 15512 12400 15564
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 13084 15512 13136 15564
rect 15384 15512 15436 15564
rect 17224 15555 17276 15564
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 1492 15376 1544 15428
rect 3056 15444 3108 15496
rect 7012 15487 7064 15496
rect 7012 15453 7021 15487
rect 7021 15453 7055 15487
rect 7055 15453 7064 15487
rect 7012 15444 7064 15453
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 11152 15487 11204 15496
rect 11152 15453 11161 15487
rect 11161 15453 11195 15487
rect 11195 15453 11204 15487
rect 11152 15444 11204 15453
rect 11244 15444 11296 15496
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 18420 15555 18472 15564
rect 18420 15521 18429 15555
rect 18429 15521 18463 15555
rect 18463 15521 18472 15555
rect 18420 15512 18472 15521
rect 22100 15512 22152 15564
rect 23296 15512 23348 15564
rect 17776 15444 17828 15496
rect 19340 15444 19392 15496
rect 21640 15444 21692 15496
rect 25320 15444 25372 15496
rect 4068 15376 4120 15428
rect 12256 15419 12308 15428
rect 12256 15385 12265 15419
rect 12265 15385 12299 15419
rect 12299 15385 12308 15419
rect 12256 15376 12308 15385
rect 14280 15376 14332 15428
rect 14372 15376 14424 15428
rect 15200 15376 15252 15428
rect 3056 15308 3108 15360
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 15568 15308 15620 15360
rect 18788 15308 18840 15360
rect 21180 15308 21232 15360
rect 24768 15308 24820 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2872 15104 2924 15156
rect 6460 15104 6512 15156
rect 10968 15104 11020 15156
rect 14648 15104 14700 15156
rect 7564 15036 7616 15088
rect 2872 14900 2924 14952
rect 6460 14968 6512 15020
rect 7472 14968 7524 15020
rect 5172 14900 5224 14952
rect 5632 14943 5684 14952
rect 5632 14909 5641 14943
rect 5641 14909 5675 14943
rect 5675 14909 5684 14943
rect 5632 14900 5684 14909
rect 7932 14943 7984 14952
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 4252 14764 4304 14816
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 4896 14764 4948 14773
rect 4988 14764 5040 14816
rect 6184 14832 6236 14884
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 10048 15036 10100 15088
rect 10140 15036 10192 15088
rect 8116 14832 8168 14884
rect 10048 14900 10100 14952
rect 14740 14968 14792 15020
rect 6460 14764 6512 14816
rect 7472 14764 7524 14816
rect 9036 14764 9088 14816
rect 9404 14764 9456 14816
rect 9680 14764 9732 14816
rect 10968 14900 11020 14952
rect 12440 14900 12492 14952
rect 12808 14943 12860 14952
rect 12808 14909 12817 14943
rect 12817 14909 12851 14943
rect 12851 14909 12860 14943
rect 12808 14900 12860 14909
rect 13176 14875 13228 14884
rect 13176 14841 13185 14875
rect 13185 14841 13219 14875
rect 13219 14841 13228 14875
rect 13176 14832 13228 14841
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 15752 14900 15804 14952
rect 18972 15036 19024 15088
rect 14832 14832 14884 14884
rect 13084 14764 13136 14816
rect 13912 14807 13964 14816
rect 13912 14773 13921 14807
rect 13921 14773 13955 14807
rect 13955 14773 13964 14807
rect 13912 14764 13964 14773
rect 15752 14764 15804 14816
rect 16672 14764 16724 14816
rect 18236 14900 18288 14952
rect 18328 14832 18380 14884
rect 20352 14900 20404 14952
rect 21548 14900 21600 14952
rect 24216 15104 24268 15156
rect 21456 14832 21508 14884
rect 17224 14764 17276 14816
rect 17868 14764 17920 14816
rect 18420 14764 18472 14816
rect 22100 14764 22152 14816
rect 23296 14764 23348 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 1216 14560 1268 14612
rect 1952 14560 2004 14612
rect 2596 14492 2648 14544
rect 2872 14560 2924 14612
rect 5172 14603 5224 14612
rect 5172 14569 5181 14603
rect 5181 14569 5215 14603
rect 5215 14569 5224 14603
rect 5172 14560 5224 14569
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 6644 14560 6696 14612
rect 7932 14560 7984 14612
rect 8392 14560 8444 14612
rect 10968 14560 11020 14612
rect 12256 14560 12308 14612
rect 9036 14492 9088 14544
rect 9864 14535 9916 14544
rect 9864 14501 9873 14535
rect 9873 14501 9907 14535
rect 9907 14501 9916 14535
rect 9864 14492 9916 14501
rect 11428 14535 11480 14544
rect 11428 14501 11437 14535
rect 11437 14501 11471 14535
rect 11471 14501 11480 14535
rect 11428 14492 11480 14501
rect 12348 14535 12400 14544
rect 12348 14501 12357 14535
rect 12357 14501 12391 14535
rect 12391 14501 12400 14535
rect 12348 14492 12400 14501
rect 3516 14424 3568 14476
rect 4160 14424 4212 14476
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 5632 14424 5684 14476
rect 8116 14467 8168 14476
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 5172 14356 5224 14408
rect 2872 14288 2924 14340
rect 3056 14288 3108 14340
rect 4528 14220 4580 14272
rect 4620 14220 4672 14272
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 14832 14492 14884 14544
rect 13176 14424 13228 14476
rect 13360 14424 13412 14476
rect 16120 14492 16172 14544
rect 16488 14560 16540 14612
rect 18052 14560 18104 14612
rect 24032 14560 24084 14612
rect 18328 14492 18380 14544
rect 15384 14424 15436 14476
rect 15476 14424 15528 14476
rect 17500 14424 17552 14476
rect 18880 14467 18932 14476
rect 18880 14433 18889 14467
rect 18889 14433 18923 14467
rect 18923 14433 18932 14467
rect 18880 14424 18932 14433
rect 20628 14424 20680 14476
rect 22284 14424 22336 14476
rect 23756 14424 23808 14476
rect 24676 14424 24728 14476
rect 8944 14356 8996 14408
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 10968 14356 11020 14408
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 12256 14356 12308 14408
rect 12716 14288 12768 14340
rect 7288 14220 7340 14272
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 11704 14220 11756 14272
rect 12532 14220 12584 14272
rect 14372 14220 14424 14272
rect 16396 14356 16448 14408
rect 15936 14288 15988 14340
rect 20536 14288 20588 14340
rect 16212 14220 16264 14272
rect 17316 14220 17368 14272
rect 17960 14220 18012 14272
rect 18236 14220 18288 14272
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 19432 14263 19484 14272
rect 19432 14229 19441 14263
rect 19441 14229 19475 14263
rect 19475 14229 19484 14263
rect 19432 14220 19484 14229
rect 20904 14220 20956 14272
rect 24860 14220 24912 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 1676 14016 1728 14068
rect 2136 14016 2188 14068
rect 5172 14016 5224 14068
rect 8116 14016 8168 14068
rect 9680 14016 9732 14068
rect 11428 14016 11480 14068
rect 12348 14016 12400 14068
rect 12808 14016 12860 14068
rect 13176 14016 13228 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 24676 14016 24728 14068
rect 2136 13880 2188 13932
rect 2964 13880 3016 13932
rect 4344 13880 4396 13932
rect 5632 13948 5684 14000
rect 6184 13948 6236 14000
rect 15844 13948 15896 14000
rect 16856 13948 16908 14000
rect 16948 13948 17000 14000
rect 20352 13948 20404 14000
rect 5540 13880 5592 13932
rect 7656 13880 7708 13932
rect 9956 13880 10008 13932
rect 11336 13880 11388 13932
rect 11980 13880 12032 13932
rect 12532 13923 12584 13932
rect 12532 13889 12541 13923
rect 12541 13889 12575 13923
rect 12575 13889 12584 13923
rect 12532 13880 12584 13889
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 2596 13812 2648 13864
rect 7288 13855 7340 13864
rect 2688 13744 2740 13796
rect 3148 13744 3200 13796
rect 3976 13744 4028 13796
rect 4620 13744 4672 13796
rect 5172 13787 5224 13796
rect 5172 13753 5181 13787
rect 5181 13753 5215 13787
rect 5215 13753 5224 13787
rect 5172 13744 5224 13753
rect 6644 13744 6696 13796
rect 7288 13821 7297 13855
rect 7297 13821 7331 13855
rect 7331 13821 7340 13855
rect 7288 13812 7340 13821
rect 7932 13812 7984 13864
rect 8760 13855 8812 13864
rect 8760 13821 8762 13855
rect 8762 13821 8812 13855
rect 8760 13812 8812 13821
rect 8852 13812 8904 13864
rect 13360 13812 13412 13864
rect 14464 13812 14516 13864
rect 15752 13812 15804 13864
rect 17316 13880 17368 13932
rect 23940 13948 23992 14000
rect 16488 13812 16540 13864
rect 16764 13812 16816 13864
rect 17776 13812 17828 13864
rect 19432 13855 19484 13864
rect 19432 13821 19441 13855
rect 19441 13821 19475 13855
rect 19475 13821 19484 13855
rect 19432 13812 19484 13821
rect 20444 13812 20496 13864
rect 204 13676 256 13728
rect 3240 13676 3292 13728
rect 4160 13719 4212 13728
rect 4160 13685 4169 13719
rect 4169 13685 4203 13719
rect 4203 13685 4212 13719
rect 6920 13719 6972 13728
rect 4160 13676 4212 13685
rect 6920 13685 6929 13719
rect 6929 13685 6963 13719
rect 6963 13685 6972 13719
rect 6920 13676 6972 13685
rect 7656 13676 7708 13728
rect 7840 13676 7892 13728
rect 8300 13676 8352 13728
rect 9036 13676 9088 13728
rect 10692 13744 10744 13796
rect 9496 13676 9548 13728
rect 10784 13676 10836 13728
rect 12440 13676 12492 13728
rect 12716 13676 12768 13728
rect 13268 13676 13320 13728
rect 14004 13676 14056 13728
rect 15476 13744 15528 13796
rect 20628 13744 20680 13796
rect 15936 13719 15988 13728
rect 15936 13685 15945 13719
rect 15945 13685 15979 13719
rect 15979 13685 15988 13719
rect 15936 13676 15988 13685
rect 16580 13719 16632 13728
rect 16580 13685 16589 13719
rect 16589 13685 16623 13719
rect 16623 13685 16632 13719
rect 16580 13676 16632 13685
rect 16856 13676 16908 13728
rect 17040 13676 17092 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 19984 13676 20036 13728
rect 22284 13676 22336 13728
rect 22560 13676 22612 13728
rect 23020 13719 23072 13728
rect 23020 13685 23029 13719
rect 23029 13685 23063 13719
rect 23063 13685 23072 13719
rect 23020 13676 23072 13685
rect 23756 13676 23808 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1308 13472 1360 13524
rect 2044 13515 2096 13524
rect 2044 13481 2053 13515
rect 2053 13481 2087 13515
rect 2087 13481 2096 13515
rect 2044 13472 2096 13481
rect 2504 13472 2556 13524
rect 3148 13515 3200 13524
rect 3148 13481 3157 13515
rect 3157 13481 3191 13515
rect 3191 13481 3200 13515
rect 3148 13472 3200 13481
rect 3516 13515 3568 13524
rect 3516 13481 3525 13515
rect 3525 13481 3559 13515
rect 3559 13481 3568 13515
rect 3516 13472 3568 13481
rect 5172 13472 5224 13524
rect 9864 13515 9916 13524
rect 9864 13481 9873 13515
rect 9873 13481 9907 13515
rect 9907 13481 9916 13515
rect 9864 13472 9916 13481
rect 3240 13404 3292 13456
rect 2504 13336 2556 13388
rect 3884 13336 3936 13388
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 5172 13336 5224 13388
rect 8852 13404 8904 13456
rect 9588 13404 9640 13456
rect 9772 13404 9824 13456
rect 11244 13472 11296 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 14004 13515 14056 13524
rect 14004 13481 14013 13515
rect 14013 13481 14047 13515
rect 14047 13481 14056 13515
rect 14004 13472 14056 13481
rect 14372 13472 14424 13524
rect 14648 13472 14700 13524
rect 16212 13472 16264 13524
rect 17040 13472 17092 13524
rect 17316 13472 17368 13524
rect 17500 13472 17552 13524
rect 18512 13472 18564 13524
rect 10692 13404 10744 13456
rect 12164 13404 12216 13456
rect 16396 13404 16448 13456
rect 18052 13404 18104 13456
rect 18880 13404 18932 13456
rect 24124 13472 24176 13524
rect 20076 13404 20128 13456
rect 27620 13404 27672 13456
rect 3148 13268 3200 13320
rect 3516 13268 3568 13320
rect 4252 13268 4304 13320
rect 7104 13336 7156 13388
rect 7932 13336 7984 13388
rect 9312 13336 9364 13388
rect 12072 13336 12124 13388
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 14096 13336 14148 13388
rect 14832 13336 14884 13388
rect 16672 13336 16724 13388
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10508 13268 10560 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11244 13268 11296 13320
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 3700 13200 3752 13252
rect 3884 13200 3936 13252
rect 13268 13200 13320 13252
rect 14280 13200 14332 13252
rect 14924 13200 14976 13252
rect 15844 13200 15896 13252
rect 2688 13132 2740 13184
rect 8116 13132 8168 13184
rect 10784 13132 10836 13184
rect 11336 13132 11388 13184
rect 13912 13132 13964 13184
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 17040 13379 17092 13388
rect 17040 13345 17049 13379
rect 17049 13345 17083 13379
rect 17083 13345 17092 13379
rect 17316 13379 17368 13388
rect 17040 13336 17092 13345
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 20720 13336 20772 13388
rect 22652 13336 22704 13388
rect 23940 13336 23992 13388
rect 24216 13336 24268 13388
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 19984 13268 20036 13320
rect 22192 13268 22244 13320
rect 22744 13268 22796 13320
rect 17040 13200 17092 13252
rect 19248 13243 19300 13252
rect 19248 13209 19257 13243
rect 19257 13209 19291 13243
rect 19291 13209 19300 13243
rect 19248 13200 19300 13209
rect 21824 13200 21876 13252
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 22836 13132 22888 13184
rect 23848 13132 23900 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2044 12928 2096 12980
rect 2228 12928 2280 12980
rect 3240 12928 3292 12980
rect 2596 12860 2648 12912
rect 4160 12928 4212 12980
rect 4988 12928 5040 12980
rect 5172 12928 5224 12980
rect 6000 12928 6052 12980
rect 7104 12971 7156 12980
rect 7104 12937 7113 12971
rect 7113 12937 7147 12971
rect 7147 12937 7156 12971
rect 7104 12928 7156 12937
rect 7196 12928 7248 12980
rect 8852 12928 8904 12980
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 10508 12928 10560 12937
rect 14832 12928 14884 12980
rect 17132 12928 17184 12980
rect 18604 12928 18656 12980
rect 5356 12860 5408 12912
rect 8300 12860 8352 12912
rect 1308 12792 1360 12844
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 5540 12835 5592 12844
rect 5540 12801 5549 12835
rect 5549 12801 5583 12835
rect 5583 12801 5592 12835
rect 5540 12792 5592 12801
rect 7012 12792 7064 12844
rect 8852 12792 8904 12844
rect 2136 12656 2188 12708
rect 2872 12588 2924 12640
rect 3240 12588 3292 12640
rect 4160 12656 4212 12708
rect 5172 12588 5224 12640
rect 5356 12699 5408 12708
rect 5356 12665 5365 12699
rect 5365 12665 5399 12699
rect 5399 12665 5408 12699
rect 5356 12656 5408 12665
rect 7104 12656 7156 12708
rect 6644 12588 6696 12640
rect 7012 12588 7064 12640
rect 7564 12588 7616 12640
rect 10692 12860 10744 12912
rect 12164 12860 12216 12912
rect 14004 12860 14056 12912
rect 16396 12860 16448 12912
rect 16672 12860 16724 12912
rect 16856 12860 16908 12912
rect 18236 12860 18288 12912
rect 19248 12903 19300 12912
rect 19248 12869 19257 12903
rect 19257 12869 19291 12903
rect 19291 12869 19300 12903
rect 19248 12860 19300 12869
rect 19984 12928 20036 12980
rect 20168 12928 20220 12980
rect 22836 12928 22888 12980
rect 23020 12928 23072 12980
rect 24216 12928 24268 12980
rect 10968 12835 11020 12844
rect 10968 12801 10977 12835
rect 10977 12801 11011 12835
rect 11011 12801 11020 12835
rect 10968 12792 11020 12801
rect 18512 12792 18564 12844
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 23664 12860 23716 12912
rect 12808 12724 12860 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14832 12724 14884 12776
rect 15476 12724 15528 12776
rect 10692 12699 10744 12708
rect 10692 12665 10701 12699
rect 10701 12665 10735 12699
rect 10735 12665 10744 12699
rect 10692 12656 10744 12665
rect 10784 12699 10836 12708
rect 10784 12665 10793 12699
rect 10793 12665 10827 12699
rect 10827 12665 10836 12699
rect 10784 12656 10836 12665
rect 14004 12656 14056 12708
rect 15384 12656 15436 12708
rect 15752 12699 15804 12708
rect 15752 12665 15761 12699
rect 15761 12665 15795 12699
rect 15795 12665 15804 12699
rect 15752 12656 15804 12665
rect 16856 12656 16908 12708
rect 17316 12656 17368 12708
rect 17960 12656 18012 12708
rect 18696 12699 18748 12708
rect 18696 12665 18705 12699
rect 18705 12665 18739 12699
rect 18739 12665 18748 12699
rect 18696 12656 18748 12665
rect 8484 12588 8536 12640
rect 9312 12588 9364 12640
rect 12072 12588 12124 12640
rect 12624 12588 12676 12640
rect 13176 12588 13228 12640
rect 13268 12588 13320 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 17040 12588 17092 12597
rect 18604 12588 18656 12640
rect 19156 12588 19208 12640
rect 19524 12588 19576 12640
rect 20444 12656 20496 12708
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 22652 12588 22704 12640
rect 23940 12631 23992 12640
rect 23940 12597 23949 12631
rect 23949 12597 23983 12631
rect 23983 12597 23992 12631
rect 23940 12588 23992 12597
rect 24216 12588 24268 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1860 12384 1912 12436
rect 1952 12384 2004 12436
rect 2320 12384 2372 12436
rect 3516 12384 3568 12436
rect 3700 12427 3752 12436
rect 3700 12393 3709 12427
rect 3709 12393 3743 12427
rect 3743 12393 3752 12427
rect 3700 12384 3752 12393
rect 7932 12427 7984 12436
rect 7932 12393 7941 12427
rect 7941 12393 7975 12427
rect 7975 12393 7984 12427
rect 7932 12384 7984 12393
rect 8852 12384 8904 12436
rect 9312 12384 9364 12436
rect 2136 12316 2188 12368
rect 6000 12316 6052 12368
rect 7564 12316 7616 12368
rect 8208 12359 8260 12368
rect 8208 12325 8217 12359
rect 8217 12325 8251 12359
rect 8251 12325 8260 12359
rect 8208 12316 8260 12325
rect 10140 12316 10192 12368
rect 10968 12384 11020 12436
rect 11428 12316 11480 12368
rect 14004 12316 14056 12368
rect 3700 12248 3752 12300
rect 4988 12248 5040 12300
rect 5356 12248 5408 12300
rect 8852 12248 8904 12300
rect 9588 12248 9640 12300
rect 11888 12248 11940 12300
rect 13544 12248 13596 12300
rect 17868 12384 17920 12436
rect 18880 12384 18932 12436
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 14464 12316 14516 12368
rect 15384 12316 15436 12368
rect 16396 12316 16448 12368
rect 17960 12316 18012 12368
rect 18696 12248 18748 12300
rect 19892 12291 19944 12300
rect 19892 12257 19910 12291
rect 19910 12257 19944 12291
rect 19892 12248 19944 12257
rect 20076 12248 20128 12300
rect 21088 12248 21140 12300
rect 23572 12291 23624 12300
rect 23572 12257 23581 12291
rect 23581 12257 23615 12291
rect 23615 12257 23624 12291
rect 23572 12248 23624 12257
rect 25136 12248 25188 12300
rect 2320 12223 2372 12232
rect 2320 12189 2329 12223
rect 2329 12189 2363 12223
rect 2363 12189 2372 12223
rect 2320 12180 2372 12189
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 6920 12180 6972 12232
rect 10692 12180 10744 12232
rect 13728 12180 13780 12232
rect 15476 12180 15528 12232
rect 4252 12155 4304 12164
rect 4252 12121 4261 12155
rect 4261 12121 4295 12155
rect 4295 12121 4304 12155
rect 4252 12112 4304 12121
rect 6552 12112 6604 12164
rect 6736 12112 6788 12164
rect 9680 12112 9732 12164
rect 9956 12112 10008 12164
rect 12440 12112 12492 12164
rect 13084 12112 13136 12164
rect 16580 12180 16632 12232
rect 17224 12180 17276 12232
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 23480 12180 23532 12189
rect 8392 12044 8444 12096
rect 12348 12044 12400 12096
rect 12624 12044 12676 12096
rect 13912 12087 13964 12096
rect 13912 12053 13921 12087
rect 13921 12053 13955 12087
rect 13955 12053 13964 12087
rect 13912 12044 13964 12053
rect 15292 12044 15344 12096
rect 15752 12044 15804 12096
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 20904 12044 20956 12096
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 25044 12044 25096 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2136 11840 2188 11892
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2964 11568 3016 11620
rect 5540 11840 5592 11892
rect 6000 11840 6052 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 8208 11840 8260 11892
rect 10140 11840 10192 11892
rect 11428 11883 11480 11892
rect 11428 11849 11437 11883
rect 11437 11849 11471 11883
rect 11471 11849 11480 11883
rect 11428 11840 11480 11849
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 14004 11840 14056 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 4160 11772 4212 11824
rect 6368 11772 6420 11824
rect 6828 11772 6880 11824
rect 3792 11747 3844 11756
rect 3792 11713 3801 11747
rect 3801 11713 3835 11747
rect 3835 11713 3844 11747
rect 3792 11704 3844 11713
rect 3976 11704 4028 11756
rect 4252 11704 4304 11756
rect 4436 11704 4488 11756
rect 9312 11772 9364 11824
rect 7104 11704 7156 11756
rect 9036 11704 9088 11756
rect 10140 11704 10192 11756
rect 10692 11704 10744 11756
rect 11704 11772 11756 11824
rect 13544 11772 13596 11824
rect 17960 11840 18012 11892
rect 19156 11883 19208 11892
rect 19156 11849 19165 11883
rect 19165 11849 19199 11883
rect 19199 11849 19208 11883
rect 19156 11840 19208 11849
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 20168 11840 20220 11892
rect 21088 11883 21140 11892
rect 21088 11849 21097 11883
rect 21097 11849 21131 11883
rect 21131 11849 21140 11883
rect 21088 11840 21140 11849
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 23572 11840 23624 11892
rect 25412 11883 25464 11892
rect 25412 11849 25421 11883
rect 25421 11849 25455 11883
rect 25455 11849 25464 11883
rect 25412 11840 25464 11849
rect 15568 11772 15620 11824
rect 17408 11772 17460 11824
rect 19892 11815 19944 11824
rect 19892 11781 19901 11815
rect 19901 11781 19935 11815
rect 19935 11781 19944 11815
rect 19892 11772 19944 11781
rect 20628 11815 20680 11824
rect 20628 11781 20637 11815
rect 20637 11781 20671 11815
rect 20671 11781 20680 11815
rect 20628 11772 20680 11781
rect 21548 11772 21600 11824
rect 12256 11704 12308 11756
rect 12808 11704 12860 11756
rect 13268 11704 13320 11756
rect 15292 11704 15344 11756
rect 16028 11704 16080 11756
rect 16396 11747 16448 11756
rect 16396 11713 16405 11747
rect 16405 11713 16439 11747
rect 16439 11713 16448 11747
rect 16396 11704 16448 11713
rect 19340 11704 19392 11756
rect 20260 11704 20312 11756
rect 21916 11747 21968 11756
rect 21916 11713 21925 11747
rect 21925 11713 21959 11747
rect 21959 11713 21968 11747
rect 21916 11704 21968 11713
rect 6276 11636 6328 11688
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 6368 11568 6420 11620
rect 1216 11500 1268 11552
rect 4988 11500 5040 11552
rect 6460 11500 6512 11552
rect 9036 11500 9088 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 10048 11500 10100 11552
rect 10784 11500 10836 11552
rect 11796 11500 11848 11552
rect 12624 11636 12676 11688
rect 15752 11636 15804 11688
rect 18880 11636 18932 11688
rect 23756 11679 23808 11688
rect 23756 11645 23765 11679
rect 23765 11645 23799 11679
rect 23799 11645 23808 11679
rect 23756 11636 23808 11645
rect 25228 11679 25280 11688
rect 25228 11645 25237 11679
rect 25237 11645 25271 11679
rect 25271 11645 25280 11679
rect 25228 11636 25280 11645
rect 14372 11611 14424 11620
rect 14372 11577 14381 11611
rect 14381 11577 14415 11611
rect 14415 11577 14424 11611
rect 14372 11568 14424 11577
rect 12256 11500 12308 11552
rect 14004 11500 14056 11552
rect 16212 11568 16264 11620
rect 17960 11568 18012 11620
rect 19524 11568 19576 11620
rect 20168 11611 20220 11620
rect 20168 11577 20177 11611
rect 20177 11577 20211 11611
rect 20211 11577 20220 11611
rect 20168 11568 20220 11577
rect 25136 11611 25188 11620
rect 17224 11500 17276 11552
rect 21364 11500 21416 11552
rect 25136 11577 25145 11611
rect 25145 11577 25179 11611
rect 25179 11577 25188 11611
rect 25136 11568 25188 11577
rect 27620 11568 27672 11620
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 5080 11296 5132 11348
rect 6368 11339 6420 11348
rect 6368 11305 6377 11339
rect 6377 11305 6411 11339
rect 6411 11305 6420 11339
rect 6368 11296 6420 11305
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7564 11296 7616 11348
rect 10140 11296 10192 11348
rect 11520 11296 11572 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 14372 11339 14424 11348
rect 1768 11228 1820 11280
rect 3976 11228 4028 11280
rect 4160 11228 4212 11280
rect 6000 11228 6052 11280
rect 8300 11228 8352 11280
rect 10048 11228 10100 11280
rect 4620 11160 4672 11212
rect 5448 11203 5500 11212
rect 5448 11169 5457 11203
rect 5457 11169 5491 11203
rect 5491 11169 5500 11203
rect 5448 11160 5500 11169
rect 7748 11160 7800 11212
rect 11980 11160 12032 11212
rect 14372 11305 14381 11339
rect 14381 11305 14415 11339
rect 14415 11305 14424 11339
rect 14372 11296 14424 11305
rect 15476 11296 15528 11348
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 20260 11339 20312 11348
rect 20260 11305 20269 11339
rect 20269 11305 20303 11339
rect 20303 11305 20312 11339
rect 20260 11296 20312 11305
rect 21548 11296 21600 11348
rect 13912 11228 13964 11280
rect 17500 11228 17552 11280
rect 2320 11092 2372 11144
rect 3424 11092 3476 11144
rect 6460 11092 6512 11144
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10692 11092 10744 11144
rect 13636 11092 13688 11144
rect 15568 11135 15620 11144
rect 388 11024 440 11076
rect 6368 11024 6420 11076
rect 9772 11024 9824 11076
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 17592 11160 17644 11212
rect 17868 11203 17920 11212
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 20720 11228 20772 11280
rect 21916 11228 21968 11280
rect 18972 11160 19024 11212
rect 20444 11160 20496 11212
rect 22008 11160 22060 11212
rect 23112 11160 23164 11212
rect 25412 11160 25464 11212
rect 18144 11092 18196 11144
rect 20904 11092 20956 11144
rect 22468 11092 22520 11144
rect 23296 11092 23348 11144
rect 24032 11092 24084 11144
rect 1768 10956 1820 11008
rect 6092 10956 6144 11008
rect 6920 10956 6972 11008
rect 10048 10956 10100 11008
rect 12808 10956 12860 11008
rect 13728 10956 13780 11008
rect 14096 10956 14148 11008
rect 15844 11024 15896 11076
rect 17960 10956 18012 11008
rect 18880 10999 18932 11008
rect 18880 10965 18889 10999
rect 18889 10965 18923 10999
rect 18923 10965 18932 10999
rect 18880 10956 18932 10965
rect 19340 10999 19392 11008
rect 19340 10965 19349 10999
rect 19349 10965 19383 10999
rect 19383 10965 19392 10999
rect 19340 10956 19392 10965
rect 20168 10956 20220 11008
rect 20260 10956 20312 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 5448 10752 5500 10804
rect 8300 10752 8352 10804
rect 10508 10752 10560 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 15292 10752 15344 10804
rect 15936 10752 15988 10804
rect 17500 10795 17552 10804
rect 17500 10761 17509 10795
rect 17509 10761 17543 10795
rect 17543 10761 17552 10795
rect 17500 10752 17552 10761
rect 17684 10752 17736 10804
rect 18144 10752 18196 10804
rect 19524 10752 19576 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 21088 10752 21140 10804
rect 4804 10684 4856 10736
rect 1860 10616 1912 10668
rect 2596 10616 2648 10668
rect 3608 10616 3660 10668
rect 5080 10616 5132 10668
rect 5172 10616 5224 10668
rect 13636 10684 13688 10736
rect 14648 10684 14700 10736
rect 15752 10684 15804 10736
rect 16028 10727 16080 10736
rect 16028 10693 16037 10727
rect 16037 10693 16071 10727
rect 16071 10693 16080 10727
rect 16028 10684 16080 10693
rect 16396 10684 16448 10736
rect 8024 10616 8076 10668
rect 10140 10616 10192 10668
rect 11980 10616 12032 10668
rect 12992 10616 13044 10668
rect 15568 10616 15620 10668
rect 19340 10616 19392 10668
rect 1768 10523 1820 10532
rect 1768 10489 1777 10523
rect 1777 10489 1811 10523
rect 1811 10489 1820 10523
rect 1768 10480 1820 10489
rect 2964 10480 3016 10532
rect 4160 10480 4212 10532
rect 4620 10412 4672 10464
rect 6184 10548 6236 10600
rect 6000 10523 6052 10532
rect 6000 10489 6009 10523
rect 6009 10489 6043 10523
rect 6043 10489 6052 10523
rect 6000 10480 6052 10489
rect 8300 10480 8352 10532
rect 9956 10523 10008 10532
rect 9956 10489 9965 10523
rect 9965 10489 9999 10523
rect 9999 10489 10008 10523
rect 9956 10480 10008 10489
rect 10048 10523 10100 10532
rect 10048 10489 10057 10523
rect 10057 10489 10091 10523
rect 10091 10489 10100 10523
rect 10048 10480 10100 10489
rect 8208 10412 8260 10464
rect 11336 10480 11388 10532
rect 15108 10480 15160 10532
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 14096 10412 14148 10464
rect 19064 10480 19116 10532
rect 18972 10412 19024 10464
rect 19524 10480 19576 10532
rect 21088 10480 21140 10532
rect 22468 10752 22520 10804
rect 23112 10795 23164 10804
rect 23112 10761 23121 10795
rect 23121 10761 23155 10795
rect 23155 10761 23164 10795
rect 23112 10752 23164 10761
rect 23480 10795 23532 10804
rect 23480 10761 23489 10795
rect 23489 10761 23523 10795
rect 23523 10761 23532 10795
rect 24952 10795 25004 10804
rect 23480 10752 23532 10761
rect 24952 10761 24961 10795
rect 24961 10761 24995 10795
rect 24995 10761 25004 10795
rect 24952 10752 25004 10761
rect 21916 10616 21968 10668
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 27712 10616 27764 10668
rect 21824 10480 21876 10532
rect 22284 10523 22336 10532
rect 22284 10489 22293 10523
rect 22293 10489 22327 10523
rect 22327 10489 22336 10523
rect 22284 10480 22336 10489
rect 23480 10412 23532 10464
rect 24860 10412 24912 10464
rect 26056 10455 26108 10464
rect 26056 10421 26065 10455
rect 26065 10421 26099 10455
rect 26099 10421 26108 10455
rect 26056 10412 26108 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1400 10208 1452 10260
rect 2320 10251 2372 10260
rect 2320 10217 2329 10251
rect 2329 10217 2363 10251
rect 2363 10217 2372 10251
rect 2320 10208 2372 10217
rect 3608 10208 3660 10260
rect 5448 10208 5500 10260
rect 7748 10208 7800 10260
rect 12348 10208 12400 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 19064 10208 19116 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 21916 10208 21968 10260
rect 24952 10208 25004 10260
rect 2504 10183 2556 10192
rect 2504 10149 2513 10183
rect 2513 10149 2547 10183
rect 2547 10149 2556 10183
rect 2504 10140 2556 10149
rect 2688 10140 2740 10192
rect 3792 10140 3844 10192
rect 4436 10140 4488 10192
rect 2320 10072 2372 10124
rect 6092 10140 6144 10192
rect 8116 10183 8168 10192
rect 8116 10149 8125 10183
rect 8125 10149 8159 10183
rect 8159 10149 8168 10183
rect 8116 10140 8168 10149
rect 8208 10183 8260 10192
rect 8208 10149 8217 10183
rect 8217 10149 8251 10183
rect 8251 10149 8260 10183
rect 8208 10140 8260 10149
rect 8852 10140 8904 10192
rect 10140 10140 10192 10192
rect 11336 10183 11388 10192
rect 11336 10149 11345 10183
rect 11345 10149 11379 10183
rect 11379 10149 11388 10183
rect 11336 10140 11388 10149
rect 11520 10140 11572 10192
rect 12532 10140 12584 10192
rect 12716 10140 12768 10192
rect 13452 10140 13504 10192
rect 13912 10140 13964 10192
rect 14004 10140 14056 10192
rect 15384 10140 15436 10192
rect 17500 10140 17552 10192
rect 18880 10183 18932 10192
rect 6000 10072 6052 10124
rect 7288 10072 7340 10124
rect 9404 10072 9456 10124
rect 9588 10072 9640 10124
rect 17684 10115 17736 10124
rect 17684 10081 17693 10115
rect 17693 10081 17727 10115
rect 17727 10081 17736 10115
rect 17684 10072 17736 10081
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 18880 10149 18889 10183
rect 18889 10149 18923 10183
rect 18923 10149 18932 10183
rect 18880 10140 18932 10149
rect 21088 10140 21140 10192
rect 23020 10140 23072 10192
rect 23664 10183 23716 10192
rect 23664 10149 23673 10183
rect 23673 10149 23707 10183
rect 23707 10149 23716 10183
rect 23664 10140 23716 10149
rect 18604 10072 18656 10124
rect 18788 10115 18840 10124
rect 18788 10081 18797 10115
rect 18797 10081 18831 10115
rect 18831 10081 18840 10115
rect 18788 10072 18840 10081
rect 20352 10072 20404 10124
rect 3424 10004 3476 10056
rect 8852 10004 8904 10056
rect 9956 10004 10008 10056
rect 12256 10004 12308 10056
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 3148 9868 3200 9920
rect 3608 9868 3660 9920
rect 5356 9868 5408 9920
rect 7656 9868 7708 9920
rect 14648 10004 14700 10056
rect 15476 10004 15528 10056
rect 14280 9936 14332 9988
rect 16212 9936 16264 9988
rect 18880 10004 18932 10056
rect 19156 10004 19208 10056
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 23204 10004 23256 10056
rect 24308 10140 24360 10192
rect 25320 10072 25372 10124
rect 23112 9936 23164 9988
rect 23940 9936 23992 9988
rect 9404 9868 9456 9920
rect 10876 9911 10928 9920
rect 10876 9877 10885 9911
rect 10885 9877 10919 9911
rect 10919 9877 10928 9911
rect 10876 9868 10928 9877
rect 16304 9911 16356 9920
rect 16304 9877 16313 9911
rect 16313 9877 16347 9911
rect 16347 9877 16356 9911
rect 16304 9868 16356 9877
rect 20444 9868 20496 9920
rect 22008 9868 22060 9920
rect 22928 9868 22980 9920
rect 23572 9868 23624 9920
rect 24676 9868 24728 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1676 9664 1728 9716
rect 3148 9664 3200 9716
rect 3792 9664 3844 9716
rect 1952 9596 2004 9648
rect 6000 9664 6052 9716
rect 6092 9664 6144 9716
rect 8116 9664 8168 9716
rect 9036 9707 9088 9716
rect 9036 9673 9045 9707
rect 9045 9673 9079 9707
rect 9079 9673 9088 9707
rect 9036 9664 9088 9673
rect 9588 9664 9640 9716
rect 11336 9664 11388 9716
rect 13084 9707 13136 9716
rect 13084 9673 13093 9707
rect 13093 9673 13127 9707
rect 13127 9673 13136 9707
rect 13084 9664 13136 9673
rect 13728 9664 13780 9716
rect 14648 9707 14700 9716
rect 14648 9673 14657 9707
rect 14657 9673 14691 9707
rect 14691 9673 14700 9707
rect 14648 9664 14700 9673
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 16764 9664 16816 9716
rect 9864 9596 9916 9648
rect 3332 9528 3384 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 5080 9528 5132 9580
rect 7564 9528 7616 9580
rect 8208 9528 8260 9580
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 1952 9503 2004 9512
rect 1952 9469 1961 9503
rect 1961 9469 1995 9503
rect 1995 9469 2004 9503
rect 1952 9460 2004 9469
rect 3884 9460 3936 9512
rect 4988 9460 5040 9512
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 2596 9392 2648 9444
rect 5356 9435 5408 9444
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5908 9435 5960 9444
rect 5356 9392 5408 9401
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 7196 9392 7248 9444
rect 9036 9392 9088 9444
rect 10048 9392 10100 9444
rect 10968 9596 11020 9648
rect 13912 9596 13964 9648
rect 16580 9596 16632 9648
rect 17684 9596 17736 9648
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 13636 9571 13688 9580
rect 13636 9537 13645 9571
rect 13645 9537 13679 9571
rect 13679 9537 13688 9571
rect 13636 9528 13688 9537
rect 14280 9571 14332 9580
rect 14280 9537 14289 9571
rect 14289 9537 14323 9571
rect 14323 9537 14332 9571
rect 14280 9528 14332 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 21088 9664 21140 9716
rect 21456 9707 21508 9716
rect 21456 9673 21465 9707
rect 21465 9673 21499 9707
rect 21499 9673 21508 9707
rect 21456 9664 21508 9673
rect 20904 9596 20956 9648
rect 23112 9707 23164 9716
rect 23112 9673 23121 9707
rect 23121 9673 23155 9707
rect 23155 9673 23164 9707
rect 23112 9664 23164 9673
rect 23572 9664 23624 9716
rect 24032 9707 24084 9716
rect 24032 9673 24041 9707
rect 24041 9673 24075 9707
rect 24075 9673 24084 9707
rect 24032 9664 24084 9673
rect 21640 9596 21692 9648
rect 22284 9639 22336 9648
rect 19064 9528 19116 9580
rect 22284 9605 22293 9639
rect 22293 9605 22327 9639
rect 22327 9605 22336 9639
rect 22284 9596 22336 9605
rect 13084 9460 13136 9512
rect 17408 9460 17460 9512
rect 13728 9435 13780 9444
rect 13728 9401 13737 9435
rect 13737 9401 13771 9435
rect 13771 9401 13780 9435
rect 13728 9392 13780 9401
rect 16304 9392 16356 9444
rect 18512 9460 18564 9512
rect 18880 9460 18932 9512
rect 23388 9528 23440 9580
rect 24584 9571 24636 9580
rect 24584 9537 24593 9571
rect 24593 9537 24627 9571
rect 24627 9537 24636 9571
rect 24584 9528 24636 9537
rect 19340 9392 19392 9444
rect 19984 9460 20036 9512
rect 21456 9392 21508 9444
rect 23296 9392 23348 9444
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 1952 9324 2004 9376
rect 2044 9324 2096 9376
rect 2688 9324 2740 9376
rect 4436 9324 4488 9376
rect 6644 9324 6696 9376
rect 12256 9367 12308 9376
rect 12256 9333 12265 9367
rect 12265 9333 12299 9367
rect 12299 9333 12308 9367
rect 12256 9324 12308 9333
rect 13084 9324 13136 9376
rect 14648 9324 14700 9376
rect 18696 9324 18748 9376
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 20352 9324 20404 9376
rect 25320 9367 25372 9376
rect 25320 9333 25329 9367
rect 25329 9333 25363 9367
rect 25363 9333 25372 9367
rect 25320 9324 25372 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2504 9120 2556 9172
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 3608 9120 3660 9172
rect 4896 9120 4948 9172
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5356 9120 5408 9172
rect 7656 9120 7708 9172
rect 7840 9163 7892 9172
rect 7840 9129 7849 9163
rect 7849 9129 7883 9163
rect 7883 9129 7892 9163
rect 7840 9120 7892 9129
rect 9220 9163 9272 9172
rect 9220 9129 9229 9163
rect 9229 9129 9263 9163
rect 9263 9129 9272 9163
rect 9220 9120 9272 9129
rect 13084 9120 13136 9172
rect 13636 9120 13688 9172
rect 1860 9052 1912 9104
rect 2320 9052 2372 9104
rect 2872 8916 2924 8968
rect 6000 9052 6052 9104
rect 7288 9052 7340 9104
rect 8300 9052 8352 9104
rect 8760 9052 8812 9104
rect 11520 9052 11572 9104
rect 16948 9120 17000 9172
rect 17868 9120 17920 9172
rect 4620 8984 4672 9036
rect 5172 8984 5224 9036
rect 5448 8984 5500 9036
rect 7380 8984 7432 9036
rect 9956 8984 10008 9036
rect 11060 9027 11112 9036
rect 11060 8993 11069 9027
rect 11069 8993 11103 9027
rect 11103 8993 11112 9027
rect 11980 9027 12032 9036
rect 11060 8984 11112 8993
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 13452 9027 13504 9036
rect 11980 8984 12032 8993
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 13912 9027 13964 9036
rect 13912 8993 13921 9027
rect 13921 8993 13955 9027
rect 13955 8993 13964 9027
rect 13912 8984 13964 8993
rect 16304 8984 16356 9036
rect 16580 8984 16632 9036
rect 16948 8984 17000 9036
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 17224 8984 17276 9036
rect 18788 9120 18840 9172
rect 21088 9120 21140 9172
rect 21640 9163 21692 9172
rect 19524 9052 19576 9104
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 18880 8984 18932 9036
rect 19340 9027 19392 9036
rect 5908 8916 5960 8968
rect 9772 8916 9824 8968
rect 10692 8916 10744 8968
rect 11152 8916 11204 8968
rect 14464 8916 14516 8968
rect 18144 8916 18196 8968
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 20904 9052 20956 9104
rect 21640 9129 21649 9163
rect 21649 9129 21683 9163
rect 21683 9129 21692 9163
rect 21640 9120 21692 9129
rect 22928 9163 22980 9172
rect 22928 9129 22937 9163
rect 22937 9129 22971 9163
rect 22971 9129 22980 9163
rect 22928 9120 22980 9129
rect 25504 9120 25556 9172
rect 22284 9052 22336 9104
rect 23112 9052 23164 9104
rect 23940 9052 23992 9104
rect 22560 8984 22612 9036
rect 20536 8916 20588 8968
rect 22744 8916 22796 8968
rect 25780 8984 25832 9036
rect 24032 8916 24084 8968
rect 24584 8916 24636 8968
rect 3516 8848 3568 8900
rect 7012 8848 7064 8900
rect 7840 8848 7892 8900
rect 11888 8848 11940 8900
rect 12532 8848 12584 8900
rect 20352 8848 20404 8900
rect 1952 8780 2004 8832
rect 2688 8823 2740 8832
rect 2688 8789 2697 8823
rect 2697 8789 2731 8823
rect 2731 8789 2740 8823
rect 2688 8780 2740 8789
rect 15844 8780 15896 8832
rect 16304 8780 16356 8832
rect 22468 8780 22520 8832
rect 24768 8848 24820 8900
rect 25228 8848 25280 8900
rect 25412 8780 25464 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 4620 8576 4672 8628
rect 5448 8576 5500 8628
rect 7380 8576 7432 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 9864 8576 9916 8628
rect 11520 8576 11572 8628
rect 12716 8576 12768 8628
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 15384 8576 15436 8628
rect 15936 8576 15988 8628
rect 16948 8576 17000 8628
rect 17224 8619 17276 8628
rect 17224 8585 17233 8619
rect 17233 8585 17267 8619
rect 17267 8585 17276 8619
rect 17224 8576 17276 8585
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 22284 8576 22336 8628
rect 22560 8576 22612 8628
rect 22744 8619 22796 8628
rect 22744 8585 22753 8619
rect 22753 8585 22787 8619
rect 22787 8585 22796 8619
rect 22744 8576 22796 8585
rect 23756 8576 23808 8628
rect 23940 8576 23992 8628
rect 24768 8576 24820 8628
rect 26148 8576 26200 8628
rect 1308 8508 1360 8560
rect 4068 8508 4120 8560
rect 9956 8508 10008 8560
rect 16396 8551 16448 8560
rect 16396 8517 16405 8551
rect 16405 8517 16439 8551
rect 16439 8517 16448 8551
rect 16396 8508 16448 8517
rect 17132 8508 17184 8560
rect 18512 8508 18564 8560
rect 2320 8440 2372 8492
rect 5448 8440 5500 8492
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 9220 8440 9272 8492
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13820 8440 13872 8492
rect 14648 8440 14700 8492
rect 17776 8372 17828 8424
rect 18788 8372 18840 8424
rect 19248 8372 19300 8424
rect 21180 8508 21232 8560
rect 21548 8508 21600 8560
rect 23020 8508 23072 8560
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 21272 8440 21324 8492
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 23204 8440 23256 8492
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 2320 8347 2372 8356
rect 2320 8313 2329 8347
rect 2329 8313 2363 8347
rect 2363 8313 2372 8347
rect 2320 8304 2372 8313
rect 2688 8304 2740 8356
rect 4344 8304 4396 8356
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 4068 8236 4120 8288
rect 5080 8279 5132 8288
rect 5080 8245 5089 8279
rect 5089 8245 5123 8279
rect 5123 8245 5132 8279
rect 5080 8236 5132 8245
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 5632 8236 5684 8288
rect 6552 8236 6604 8288
rect 6828 8236 6880 8288
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 11152 8304 11204 8356
rect 11888 8304 11940 8356
rect 12440 8236 12492 8288
rect 13268 8304 13320 8356
rect 14280 8347 14332 8356
rect 14280 8313 14289 8347
rect 14289 8313 14323 8347
rect 14323 8313 14332 8347
rect 14280 8304 14332 8313
rect 15844 8347 15896 8356
rect 15844 8313 15853 8347
rect 15853 8313 15887 8347
rect 15887 8313 15896 8347
rect 15844 8304 15896 8313
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 19984 8372 20036 8424
rect 25412 8415 25464 8424
rect 25412 8381 25421 8415
rect 25421 8381 25455 8415
rect 25455 8381 25464 8415
rect 25412 8372 25464 8381
rect 15936 8304 15988 8313
rect 15384 8236 15436 8288
rect 15660 8279 15712 8288
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 18880 8279 18932 8288
rect 18880 8245 18889 8279
rect 18889 8245 18923 8279
rect 18923 8245 18932 8279
rect 18880 8236 18932 8245
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 23020 8304 23072 8356
rect 23756 8304 23808 8356
rect 21180 8236 21232 8245
rect 25780 8236 25832 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1676 8032 1728 8084
rect 2872 8032 2924 8084
rect 6644 8032 6696 8084
rect 6828 8032 6880 8084
rect 7012 8032 7064 8084
rect 11060 8075 11112 8084
rect 11060 8041 11069 8075
rect 11069 8041 11103 8075
rect 11103 8041 11112 8075
rect 11060 8032 11112 8041
rect 2504 7964 2556 8016
rect 3148 7964 3200 8016
rect 3976 7964 4028 8016
rect 4436 7964 4488 8016
rect 5356 7964 5408 8016
rect 5632 8007 5684 8016
rect 5632 7973 5641 8007
rect 5641 7973 5675 8007
rect 5675 7973 5684 8007
rect 5632 7964 5684 7973
rect 6000 7964 6052 8016
rect 6460 7964 6512 8016
rect 7288 8007 7340 8016
rect 7288 7973 7297 8007
rect 7297 7973 7331 8007
rect 7331 7973 7340 8007
rect 9864 8007 9916 8016
rect 7288 7964 7340 7973
rect 5080 7896 5132 7948
rect 7656 7896 7708 7948
rect 7932 7896 7984 7948
rect 9864 7973 9873 8007
rect 9873 7973 9907 8007
rect 9907 7973 9916 8007
rect 9864 7964 9916 7973
rect 9956 7964 10008 8016
rect 11704 8032 11756 8084
rect 14280 8075 14332 8084
rect 14280 8041 14289 8075
rect 14289 8041 14323 8075
rect 14323 8041 14332 8075
rect 14280 8032 14332 8041
rect 16120 8075 16172 8084
rect 16120 8041 16129 8075
rect 16129 8041 16163 8075
rect 16163 8041 16172 8075
rect 16120 8032 16172 8041
rect 16304 8075 16356 8084
rect 16304 8041 16313 8075
rect 16313 8041 16347 8075
rect 16347 8041 16356 8075
rect 16304 8032 16356 8041
rect 17224 8032 17276 8084
rect 11980 7964 12032 8016
rect 12900 8007 12952 8016
rect 12900 7973 12909 8007
rect 12909 7973 12943 8007
rect 12943 7973 12952 8007
rect 12900 7964 12952 7973
rect 12992 8007 13044 8016
rect 12992 7973 13001 8007
rect 13001 7973 13035 8007
rect 13035 7973 13044 8007
rect 19340 8032 19392 8084
rect 19984 8032 20036 8084
rect 21272 8032 21324 8084
rect 23020 8075 23072 8084
rect 23020 8041 23029 8075
rect 23029 8041 23063 8075
rect 23063 8041 23072 8075
rect 23020 8032 23072 8041
rect 23204 8032 23256 8084
rect 12992 7964 13044 7973
rect 9220 7896 9272 7948
rect 15660 7896 15712 7948
rect 16580 7896 16632 7948
rect 3792 7828 3844 7880
rect 2320 7760 2372 7812
rect 4344 7828 4396 7880
rect 6000 7871 6052 7880
rect 6000 7837 6009 7871
rect 6009 7837 6043 7871
rect 6043 7837 6052 7871
rect 6000 7828 6052 7837
rect 6920 7828 6972 7880
rect 7196 7828 7248 7880
rect 10048 7871 10100 7880
rect 4896 7760 4948 7812
rect 10048 7837 10057 7871
rect 10057 7837 10091 7871
rect 10091 7837 10100 7871
rect 10048 7828 10100 7837
rect 11704 7828 11756 7880
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 14280 7828 14332 7880
rect 16396 7828 16448 7880
rect 16948 7896 17000 7948
rect 17316 7896 17368 7948
rect 18696 7964 18748 8016
rect 18880 7964 18932 8016
rect 17868 7896 17920 7948
rect 18788 7896 18840 7948
rect 22560 7964 22612 8016
rect 24768 8075 24820 8084
rect 24768 8041 24777 8075
rect 24777 8041 24811 8075
rect 24811 8041 24820 8075
rect 24768 8032 24820 8041
rect 17776 7828 17828 7880
rect 19524 7896 19576 7948
rect 20904 7896 20956 7948
rect 21456 7896 21508 7948
rect 19248 7828 19300 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 24952 7828 25004 7880
rect 11888 7803 11940 7812
rect 11888 7769 11897 7803
rect 11897 7769 11931 7803
rect 11931 7769 11940 7803
rect 11888 7760 11940 7769
rect 13084 7760 13136 7812
rect 15844 7760 15896 7812
rect 5172 7735 5224 7744
rect 5172 7701 5181 7735
rect 5181 7701 5215 7735
rect 5215 7701 5224 7735
rect 5172 7692 5224 7701
rect 5356 7692 5408 7744
rect 7104 7692 7156 7744
rect 12256 7692 12308 7744
rect 12716 7735 12768 7744
rect 12716 7701 12725 7735
rect 12725 7701 12759 7735
rect 12759 7701 12768 7735
rect 12716 7692 12768 7701
rect 15568 7692 15620 7744
rect 15660 7692 15712 7744
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 21364 7692 21416 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2596 7488 2648 7540
rect 3792 7488 3844 7540
rect 3976 7488 4028 7540
rect 8852 7488 8904 7540
rect 9036 7531 9088 7540
rect 9036 7497 9045 7531
rect 9045 7497 9079 7531
rect 9079 7497 9088 7531
rect 9036 7488 9088 7497
rect 9864 7488 9916 7540
rect 11980 7488 12032 7540
rect 13544 7488 13596 7540
rect 14740 7488 14792 7540
rect 1676 7352 1728 7404
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 4528 7352 4580 7404
rect 5908 7352 5960 7404
rect 6736 7352 6788 7404
rect 9128 7420 9180 7472
rect 9772 7463 9824 7472
rect 9772 7429 9781 7463
rect 9781 7429 9815 7463
rect 9815 7429 9824 7463
rect 9772 7420 9824 7429
rect 11520 7420 11572 7472
rect 16396 7488 16448 7540
rect 16580 7488 16632 7540
rect 21088 7488 21140 7540
rect 22376 7488 22428 7540
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 16948 7420 17000 7472
rect 18880 7463 18932 7472
rect 18880 7429 18889 7463
rect 18889 7429 18923 7463
rect 18923 7429 18932 7463
rect 18880 7420 18932 7429
rect 22560 7463 22612 7472
rect 22560 7429 22569 7463
rect 22569 7429 22603 7463
rect 22603 7429 22612 7463
rect 22560 7420 22612 7429
rect 22836 7420 22888 7472
rect 4804 7284 4856 7336
rect 6276 7284 6328 7336
rect 7288 7327 7340 7336
rect 1860 7216 1912 7268
rect 4068 7216 4120 7268
rect 5172 7216 5224 7268
rect 6736 7216 6788 7268
rect 6828 7216 6880 7268
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 8116 7284 8168 7336
rect 2136 7148 2188 7200
rect 3148 7148 3200 7200
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 6460 7148 6512 7200
rect 8760 7216 8812 7268
rect 9036 7216 9088 7268
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 12992 7352 13044 7404
rect 12716 7284 12768 7336
rect 14740 7284 14792 7336
rect 16580 7352 16632 7404
rect 18604 7352 18656 7404
rect 16212 7284 16264 7336
rect 16948 7284 17000 7336
rect 17316 7284 17368 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 18788 7284 18840 7336
rect 19064 7327 19116 7336
rect 19064 7293 19073 7327
rect 19073 7293 19107 7327
rect 19107 7293 19116 7327
rect 19064 7284 19116 7293
rect 19248 7284 19300 7336
rect 21456 7352 21508 7404
rect 19984 7284 20036 7336
rect 7656 7148 7708 7200
rect 12440 7148 12492 7200
rect 16672 7216 16724 7268
rect 17776 7259 17828 7268
rect 17776 7225 17785 7259
rect 17785 7225 17819 7259
rect 17819 7225 17828 7259
rect 17776 7216 17828 7225
rect 19432 7216 19484 7268
rect 21272 7284 21324 7336
rect 24216 7352 24268 7404
rect 21088 7216 21140 7268
rect 24124 7259 24176 7268
rect 24124 7225 24133 7259
rect 24133 7225 24167 7259
rect 24167 7225 24176 7259
rect 24124 7216 24176 7225
rect 20904 7191 20956 7200
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 21364 7148 21416 7200
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1676 6944 1728 6996
rect 2596 6944 2648 6996
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 5632 6944 5684 6996
rect 6000 6944 6052 6996
rect 9128 6987 9180 6996
rect 9128 6953 9137 6987
rect 9137 6953 9171 6987
rect 9171 6953 9180 6987
rect 9128 6944 9180 6953
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 12900 6944 12952 6996
rect 2044 6876 2096 6928
rect 4528 6876 4580 6928
rect 4896 6876 4948 6928
rect 6460 6876 6512 6928
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 12440 6876 12492 6928
rect 13176 6876 13228 6928
rect 14556 6944 14608 6996
rect 18328 6944 18380 6996
rect 18788 6944 18840 6996
rect 19432 6944 19484 6996
rect 15660 6876 15712 6928
rect 16212 6876 16264 6928
rect 5540 6808 5592 6860
rect 7012 6808 7064 6860
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 14464 6808 14516 6860
rect 15844 6808 15896 6860
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 16672 6808 16724 6860
rect 17316 6876 17368 6928
rect 18604 6876 18656 6928
rect 17224 6808 17276 6860
rect 17776 6808 17828 6860
rect 21088 6944 21140 6996
rect 22100 6987 22152 6996
rect 21180 6876 21232 6928
rect 22100 6953 22109 6987
rect 22109 6953 22143 6987
rect 22143 6953 22152 6987
rect 22100 6944 22152 6953
rect 24124 6944 24176 6996
rect 21364 6876 21416 6928
rect 21824 6919 21876 6928
rect 21824 6885 21833 6919
rect 21833 6885 21867 6919
rect 21867 6885 21876 6919
rect 21824 6876 21876 6885
rect 25044 6944 25096 6996
rect 24676 6876 24728 6928
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 2136 6740 2188 6792
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 4620 6740 4672 6792
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10692 6740 10744 6792
rect 11336 6740 11388 6792
rect 21548 6740 21600 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 24768 6740 24820 6749
rect 1216 6672 1268 6724
rect 2504 6672 2556 6724
rect 3056 6672 3108 6724
rect 5448 6672 5500 6724
rect 6736 6715 6788 6724
rect 6736 6681 6745 6715
rect 6745 6681 6779 6715
rect 6779 6681 6788 6715
rect 6736 6672 6788 6681
rect 15568 6672 15620 6724
rect 16948 6672 17000 6724
rect 3976 6604 4028 6656
rect 4344 6604 4396 6656
rect 6184 6604 6236 6656
rect 6828 6604 6880 6656
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 16304 6604 16356 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 20720 6604 20772 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 3240 6400 3292 6452
rect 4896 6443 4948 6452
rect 2504 6264 2556 6316
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 6092 6400 6144 6452
rect 6460 6400 6512 6452
rect 8116 6400 8168 6452
rect 9864 6400 9916 6452
rect 11520 6400 11572 6452
rect 12992 6400 13044 6452
rect 14464 6400 14516 6452
rect 15384 6400 15436 6452
rect 16580 6400 16632 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 18420 6400 18472 6452
rect 4068 6264 4120 6316
rect 9128 6264 9180 6316
rect 9496 6264 9548 6316
rect 9864 6264 9916 6316
rect 6828 6239 6880 6248
rect 2596 6128 2648 6180
rect 3424 6060 3476 6112
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 7196 6196 7248 6248
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 8760 6128 8812 6137
rect 11060 6332 11112 6384
rect 11244 6332 11296 6384
rect 16304 6332 16356 6384
rect 18604 6332 18656 6384
rect 19984 6400 20036 6452
rect 22744 6443 22796 6452
rect 22744 6409 22753 6443
rect 22753 6409 22787 6443
rect 22787 6409 22796 6443
rect 22744 6400 22796 6409
rect 25044 6400 25096 6452
rect 24952 6332 25004 6384
rect 10784 6264 10836 6316
rect 11888 6264 11940 6316
rect 11612 6196 11664 6248
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 15752 6264 15804 6316
rect 16764 6307 16816 6316
rect 16764 6273 16773 6307
rect 16773 6273 16807 6307
rect 16807 6273 16816 6307
rect 16764 6264 16816 6273
rect 18880 6264 18932 6316
rect 23848 6307 23900 6316
rect 16304 6239 16356 6248
rect 16304 6205 16313 6239
rect 16313 6205 16347 6239
rect 16347 6205 16356 6239
rect 16304 6196 16356 6205
rect 16580 6239 16632 6248
rect 16580 6205 16589 6239
rect 16589 6205 16623 6239
rect 16623 6205 16632 6239
rect 16580 6196 16632 6205
rect 17592 6196 17644 6248
rect 17960 6196 18012 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19248 6196 19300 6248
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 23848 6273 23857 6307
rect 23857 6273 23891 6307
rect 23891 6273 23900 6307
rect 23848 6264 23900 6273
rect 24124 6264 24176 6316
rect 24768 6264 24820 6316
rect 10784 6171 10836 6180
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 10968 6128 11020 6180
rect 12992 6171 13044 6180
rect 12992 6137 13001 6171
rect 13001 6137 13035 6171
rect 13035 6137 13044 6171
rect 12992 6128 13044 6137
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 6736 6060 6788 6112
rect 7840 6060 7892 6112
rect 8300 6060 8352 6112
rect 10140 6060 10192 6112
rect 11060 6060 11112 6112
rect 11428 6060 11480 6112
rect 18696 6128 18748 6180
rect 21180 6128 21232 6180
rect 15844 6103 15896 6112
rect 15844 6069 15853 6103
rect 15853 6069 15887 6103
rect 15887 6069 15896 6103
rect 15844 6060 15896 6069
rect 18328 6060 18380 6112
rect 20076 6060 20128 6112
rect 21364 6060 21416 6112
rect 25228 6196 25280 6248
rect 22100 6171 22152 6180
rect 22100 6137 22109 6171
rect 22109 6137 22143 6171
rect 22143 6137 22152 6171
rect 22100 6128 22152 6137
rect 22744 6128 22796 6180
rect 25044 6128 25096 6180
rect 24676 6060 24728 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2228 5856 2280 5908
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 9128 5899 9180 5908
rect 7196 5856 7248 5865
rect 2688 5788 2740 5840
rect 6460 5788 6512 5840
rect 8760 5788 8812 5840
rect 9128 5865 9137 5899
rect 9137 5865 9171 5899
rect 9171 5865 9180 5899
rect 9128 5856 9180 5865
rect 9772 5856 9824 5908
rect 10692 5856 10744 5908
rect 14556 5899 14608 5908
rect 10784 5788 10836 5840
rect 11428 5788 11480 5840
rect 12440 5831 12492 5840
rect 12440 5797 12449 5831
rect 12449 5797 12483 5831
rect 12483 5797 12492 5831
rect 12440 5788 12492 5797
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 13452 5788 13504 5840
rect 1124 5720 1176 5772
rect 4252 5763 4304 5772
rect 4252 5729 4261 5763
rect 4261 5729 4295 5763
rect 4295 5729 4304 5763
rect 4252 5720 4304 5729
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3056 5627 3108 5636
rect 3056 5593 3065 5627
rect 3065 5593 3099 5627
rect 3099 5593 3108 5627
rect 3056 5584 3108 5593
rect 5540 5652 5592 5704
rect 7472 5720 7524 5772
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 9496 5720 9548 5772
rect 10876 5720 10928 5772
rect 11520 5720 11572 5772
rect 15568 5856 15620 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 16120 5720 16172 5772
rect 16580 5856 16632 5908
rect 17132 5856 17184 5908
rect 17224 5856 17276 5908
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 19064 5856 19116 5908
rect 20260 5856 20312 5908
rect 22560 5899 22612 5908
rect 22560 5865 22569 5899
rect 22569 5865 22603 5899
rect 22603 5865 22612 5899
rect 22560 5856 22612 5865
rect 22836 5856 22888 5908
rect 23848 5899 23900 5908
rect 16856 5763 16908 5772
rect 16856 5729 16865 5763
rect 16865 5729 16899 5763
rect 16899 5729 16908 5763
rect 16856 5720 16908 5729
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 17960 5788 18012 5840
rect 18236 5763 18288 5772
rect 18236 5729 18245 5763
rect 18245 5729 18279 5763
rect 18279 5729 18288 5763
rect 18236 5720 18288 5729
rect 21272 5788 21324 5840
rect 23848 5865 23857 5899
rect 23857 5865 23891 5899
rect 23891 5865 23900 5899
rect 23848 5856 23900 5865
rect 25228 5788 25280 5840
rect 9312 5652 9364 5704
rect 11060 5652 11112 5704
rect 5448 5584 5500 5636
rect 8116 5584 8168 5636
rect 10048 5584 10100 5636
rect 13728 5652 13780 5704
rect 15660 5652 15712 5704
rect 17408 5652 17460 5704
rect 19340 5720 19392 5772
rect 20628 5720 20680 5772
rect 21180 5720 21232 5772
rect 22192 5763 22244 5772
rect 22192 5729 22201 5763
rect 22201 5729 22235 5763
rect 22235 5729 22244 5763
rect 22192 5720 22244 5729
rect 22652 5720 22704 5772
rect 24216 5695 24268 5704
rect 22652 5584 22704 5636
rect 24216 5661 24225 5695
rect 24225 5661 24259 5695
rect 24259 5661 24268 5695
rect 24216 5652 24268 5661
rect 24768 5584 24820 5636
rect 2136 5559 2188 5568
rect 2136 5525 2145 5559
rect 2145 5525 2179 5559
rect 2179 5525 2188 5559
rect 2136 5516 2188 5525
rect 5356 5516 5408 5568
rect 6828 5559 6880 5568
rect 6828 5525 6837 5559
rect 6837 5525 6871 5559
rect 6871 5525 6880 5559
rect 6828 5516 6880 5525
rect 8208 5516 8260 5568
rect 10140 5516 10192 5568
rect 10324 5516 10376 5568
rect 11060 5516 11112 5568
rect 12164 5516 12216 5568
rect 21824 5559 21876 5568
rect 21824 5525 21833 5559
rect 21833 5525 21867 5559
rect 21867 5525 21876 5559
rect 21824 5516 21876 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 1124 5312 1176 5364
rect 1860 5312 1912 5364
rect 4252 5312 4304 5364
rect 6368 5312 6420 5364
rect 8024 5312 8076 5364
rect 9496 5312 9548 5364
rect 9864 5312 9916 5364
rect 11520 5355 11572 5364
rect 3148 5244 3200 5296
rect 5632 5244 5684 5296
rect 9772 5244 9824 5296
rect 10876 5244 10928 5296
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 15568 5312 15620 5364
rect 17408 5355 17460 5364
rect 17408 5321 17417 5355
rect 17417 5321 17451 5355
rect 17451 5321 17460 5355
rect 17408 5312 17460 5321
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18788 5355 18840 5364
rect 18788 5321 18797 5355
rect 18797 5321 18831 5355
rect 18831 5321 18840 5355
rect 18788 5312 18840 5321
rect 21088 5355 21140 5364
rect 21088 5321 21097 5355
rect 21097 5321 21131 5355
rect 21131 5321 21140 5355
rect 21088 5312 21140 5321
rect 21272 5312 21324 5364
rect 14648 5287 14700 5296
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 3056 5176 3108 5228
rect 4068 5176 4120 5228
rect 8576 5176 8628 5228
rect 10692 5176 10744 5228
rect 11428 5176 11480 5228
rect 14648 5253 14657 5287
rect 14657 5253 14691 5287
rect 14691 5253 14700 5287
rect 14648 5244 14700 5253
rect 13268 5176 13320 5228
rect 12716 5108 12768 5160
rect 1860 5040 1912 5092
rect 2228 5040 2280 5092
rect 2688 5040 2740 5092
rect 2596 4972 2648 5024
rect 4528 5040 4580 5092
rect 5356 5083 5408 5092
rect 5356 5049 5365 5083
rect 5365 5049 5399 5083
rect 5399 5049 5408 5083
rect 5356 5040 5408 5049
rect 6000 5040 6052 5092
rect 6920 5083 6972 5092
rect 6920 5049 6929 5083
rect 6929 5049 6963 5083
rect 6963 5049 6972 5083
rect 6920 5040 6972 5049
rect 10324 5083 10376 5092
rect 6368 4972 6420 5024
rect 6552 4972 6604 5024
rect 10324 5049 10333 5083
rect 10333 5049 10367 5083
rect 10367 5049 10376 5083
rect 10324 5040 10376 5049
rect 11612 5040 11664 5092
rect 15384 5108 15436 5160
rect 14096 5083 14148 5092
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 9312 5015 9364 5024
rect 9312 4981 9321 5015
rect 9321 4981 9355 5015
rect 9355 4981 9364 5015
rect 9312 4972 9364 4981
rect 14096 5049 14105 5083
rect 14105 5049 14139 5083
rect 14139 5049 14148 5083
rect 14096 5040 14148 5049
rect 16856 5040 16908 5092
rect 17500 5040 17552 5092
rect 19064 5151 19116 5160
rect 19064 5117 19073 5151
rect 19073 5117 19107 5151
rect 19107 5117 19116 5151
rect 19064 5108 19116 5117
rect 19984 5151 20036 5160
rect 19432 5040 19484 5092
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 21824 5219 21876 5228
rect 21824 5185 21833 5219
rect 21833 5185 21867 5219
rect 21867 5185 21876 5219
rect 21824 5176 21876 5185
rect 22560 5312 22612 5364
rect 22744 5355 22796 5364
rect 22744 5321 22753 5355
rect 22753 5321 22787 5355
rect 22787 5321 22796 5355
rect 22744 5312 22796 5321
rect 23388 5312 23440 5364
rect 24216 5312 24268 5364
rect 25228 5355 25280 5364
rect 24400 5244 24452 5296
rect 25228 5321 25237 5355
rect 25237 5321 25271 5355
rect 25271 5321 25280 5355
rect 25228 5312 25280 5321
rect 24768 5219 24820 5228
rect 24768 5185 24777 5219
rect 24777 5185 24811 5219
rect 24811 5185 24820 5219
rect 24768 5176 24820 5185
rect 17776 4972 17828 5024
rect 19984 4972 20036 5024
rect 24400 5083 24452 5092
rect 24400 5049 24409 5083
rect 24409 5049 24443 5083
rect 24443 5049 24452 5083
rect 24400 5040 24452 5049
rect 25136 4972 25188 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 2504 4768 2556 4820
rect 5356 4768 5408 4820
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 5908 4768 5960 4820
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 7840 4811 7892 4820
rect 7840 4777 7849 4811
rect 7849 4777 7883 4811
rect 7883 4777 7892 4811
rect 7840 4768 7892 4777
rect 8576 4768 8628 4820
rect 11244 4768 11296 4820
rect 12900 4811 12952 4820
rect 12900 4777 12909 4811
rect 12909 4777 12943 4811
rect 12943 4777 12952 4811
rect 12900 4768 12952 4777
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 15384 4768 15436 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 17960 4811 18012 4820
rect 17960 4777 17969 4811
rect 17969 4777 18003 4811
rect 18003 4777 18012 4811
rect 17960 4768 18012 4777
rect 18972 4768 19024 4820
rect 19340 4768 19392 4820
rect 20628 4811 20680 4820
rect 20628 4777 20637 4811
rect 20637 4777 20671 4811
rect 20671 4777 20680 4811
rect 20628 4768 20680 4777
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 22192 4811 22244 4820
rect 22192 4777 22201 4811
rect 22201 4777 22235 4811
rect 22235 4777 22244 4811
rect 22192 4768 22244 4777
rect 24124 4811 24176 4820
rect 24124 4777 24133 4811
rect 24133 4777 24167 4811
rect 24167 4777 24176 4811
rect 24124 4768 24176 4777
rect 24676 4811 24728 4820
rect 24676 4777 24685 4811
rect 24685 4777 24719 4811
rect 24719 4777 24728 4811
rect 24676 4768 24728 4777
rect 2596 4743 2648 4752
rect 2596 4709 2605 4743
rect 2605 4709 2639 4743
rect 2639 4709 2648 4743
rect 2596 4700 2648 4709
rect 3148 4743 3200 4752
rect 3148 4709 3157 4743
rect 3157 4709 3191 4743
rect 3191 4709 3200 4743
rect 3148 4700 3200 4709
rect 3976 4700 4028 4752
rect 4620 4700 4672 4752
rect 6460 4700 6512 4752
rect 8116 4743 8168 4752
rect 8116 4709 8125 4743
rect 8125 4709 8159 4743
rect 8159 4709 8168 4743
rect 8116 4700 8168 4709
rect 8208 4743 8260 4752
rect 8208 4709 8217 4743
rect 8217 4709 8251 4743
rect 8251 4709 8260 4743
rect 8208 4700 8260 4709
rect 9312 4700 9364 4752
rect 9772 4700 9824 4752
rect 10784 4700 10836 4752
rect 12716 4700 12768 4752
rect 1768 4632 1820 4684
rect 11704 4675 11756 4684
rect 3148 4564 3200 4616
rect 6644 4564 6696 4616
rect 8760 4607 8812 4616
rect 8760 4573 8769 4607
rect 8769 4573 8803 4607
rect 8803 4573 8812 4607
rect 8760 4564 8812 4573
rect 9496 4564 9548 4616
rect 10048 4607 10100 4616
rect 10048 4573 10057 4607
rect 10057 4573 10091 4607
rect 10091 4573 10100 4607
rect 10048 4564 10100 4573
rect 4528 4496 4580 4548
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 17040 4700 17092 4752
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 15660 4632 15712 4684
rect 18236 4675 18288 4684
rect 15752 4564 15804 4616
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 11336 4496 11388 4548
rect 16580 4496 16632 4548
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 18972 4675 19024 4684
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 17408 4564 17460 4616
rect 18972 4641 18981 4675
rect 18981 4641 19015 4675
rect 19015 4641 19024 4675
rect 18972 4632 19024 4641
rect 21088 4700 21140 4752
rect 21916 4700 21968 4752
rect 22560 4700 22612 4752
rect 22836 4743 22888 4752
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 25044 4632 25096 4684
rect 21088 4564 21140 4616
rect 22008 4564 22060 4616
rect 5356 4428 5408 4480
rect 8300 4428 8352 4480
rect 13084 4428 13136 4480
rect 15752 4471 15804 4480
rect 15752 4437 15761 4471
rect 15761 4437 15795 4471
rect 15795 4437 15804 4471
rect 15752 4428 15804 4437
rect 16304 4428 16356 4480
rect 19156 4428 19208 4480
rect 22468 4496 22520 4548
rect 22652 4496 22704 4548
rect 22836 4428 22888 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 3976 4224 4028 4276
rect 8208 4224 8260 4276
rect 9772 4267 9824 4276
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 11336 4267 11388 4276
rect 11336 4233 11345 4267
rect 11345 4233 11379 4267
rect 11379 4233 11388 4267
rect 11336 4224 11388 4233
rect 11704 4267 11756 4276
rect 11704 4233 11713 4267
rect 11713 4233 11747 4267
rect 11747 4233 11756 4267
rect 11704 4224 11756 4233
rect 13084 4224 13136 4276
rect 15752 4224 15804 4276
rect 16488 4224 16540 4276
rect 17132 4224 17184 4276
rect 17408 4267 17460 4276
rect 17408 4233 17417 4267
rect 17417 4233 17451 4267
rect 17451 4233 17460 4267
rect 17408 4224 17460 4233
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 18236 4267 18288 4276
rect 18236 4233 18245 4267
rect 18245 4233 18279 4267
rect 18279 4233 18288 4267
rect 18236 4224 18288 4233
rect 20168 4224 20220 4276
rect 22468 4224 22520 4276
rect 22560 4224 22612 4276
rect 25044 4267 25096 4276
rect 25044 4233 25053 4267
rect 25053 4233 25087 4267
rect 25087 4233 25096 4267
rect 25044 4224 25096 4233
rect 26148 4267 26200 4276
rect 26148 4233 26157 4267
rect 26157 4233 26191 4267
rect 26191 4233 26200 4267
rect 26148 4224 26200 4233
rect 1768 4156 1820 4208
rect 2228 4156 2280 4208
rect 3424 4199 3476 4208
rect 3424 4165 3433 4199
rect 3433 4165 3467 4199
rect 3467 4165 3476 4199
rect 3424 4156 3476 4165
rect 6460 4156 6512 4208
rect 7748 4199 7800 4208
rect 7748 4165 7757 4199
rect 7757 4165 7791 4199
rect 7791 4165 7800 4199
rect 7748 4156 7800 4165
rect 2320 4088 2372 4140
rect 5540 4131 5592 4140
rect 1860 4020 1912 4072
rect 2320 3884 2372 3936
rect 5540 4097 5549 4131
rect 5549 4097 5583 4131
rect 5583 4097 5592 4131
rect 5540 4088 5592 4097
rect 4436 4020 4488 4072
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 9496 4156 9548 4208
rect 14464 4156 14516 4208
rect 22836 4156 22888 4208
rect 23112 4156 23164 4208
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9772 4088 9824 4140
rect 10140 4088 10192 4140
rect 12256 4063 12308 4072
rect 3608 3952 3660 4004
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5356 3952 5408 3961
rect 7748 3952 7800 4004
rect 3792 3927 3844 3936
rect 3792 3893 3801 3927
rect 3801 3893 3835 3927
rect 3835 3893 3844 3927
rect 3792 3884 3844 3893
rect 7932 3884 7984 3936
rect 9772 3952 9824 4004
rect 12256 4029 12265 4063
rect 12265 4029 12299 4063
rect 12299 4029 12308 4063
rect 18328 4088 18380 4140
rect 12256 4020 12308 4029
rect 14464 4063 14516 4072
rect 10324 3995 10376 4004
rect 10324 3961 10333 3995
rect 10333 3961 10367 3995
rect 10367 3961 10376 3995
rect 10324 3952 10376 3961
rect 10968 3995 11020 4004
rect 10140 3884 10192 3936
rect 10968 3961 10977 3995
rect 10977 3961 11011 3995
rect 11011 3961 11020 3995
rect 10968 3952 11020 3961
rect 11704 3952 11756 4004
rect 14464 4029 14473 4063
rect 14473 4029 14507 4063
rect 14507 4029 14516 4063
rect 14464 4020 14516 4029
rect 16580 4020 16632 4072
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 19064 4088 19116 4140
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 19984 4063 20036 4072
rect 19984 4029 19993 4063
rect 19993 4029 20027 4063
rect 20027 4029 20036 4063
rect 19984 4020 20036 4029
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 14832 3927 14884 3936
rect 13820 3884 13872 3893
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 18880 3927 18932 3936
rect 18880 3893 18889 3927
rect 18889 3893 18923 3927
rect 18923 3893 18932 3927
rect 18880 3884 18932 3893
rect 20720 3884 20772 3936
rect 21180 3884 21232 3936
rect 26148 4020 26200 4072
rect 24768 3995 24820 4004
rect 23756 3884 23808 3936
rect 24768 3961 24777 3995
rect 24777 3961 24811 3995
rect 24811 3961 24820 3995
rect 24768 3952 24820 3961
rect 24676 3884 24728 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 2412 3680 2464 3732
rect 20 3612 72 3664
rect 1584 3612 1636 3664
rect 5080 3680 5132 3732
rect 6552 3723 6604 3732
rect 6552 3689 6561 3723
rect 6561 3689 6595 3723
rect 6595 3689 6604 3723
rect 6552 3680 6604 3689
rect 9128 3723 9180 3732
rect 2688 3612 2740 3664
rect 3148 3655 3200 3664
rect 3148 3621 3157 3655
rect 3157 3621 3191 3655
rect 3191 3621 3200 3655
rect 3148 3612 3200 3621
rect 4160 3655 4212 3664
rect 4160 3621 4169 3655
rect 4169 3621 4203 3655
rect 4203 3621 4212 3655
rect 4160 3612 4212 3621
rect 4436 3612 4488 3664
rect 6368 3612 6420 3664
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 5540 3544 5592 3596
rect 8208 3655 8260 3664
rect 8208 3621 8217 3655
rect 8217 3621 8251 3655
rect 8251 3621 8260 3655
rect 8208 3612 8260 3621
rect 8760 3655 8812 3664
rect 8760 3621 8769 3655
rect 8769 3621 8803 3655
rect 8803 3621 8812 3655
rect 8760 3612 8812 3621
rect 1584 3476 1636 3528
rect 6828 3476 6880 3528
rect 7564 3519 7616 3528
rect 7564 3485 7573 3519
rect 7573 3485 7607 3519
rect 7607 3485 7616 3519
rect 7564 3476 7616 3485
rect 9128 3689 9137 3723
rect 9137 3689 9171 3723
rect 9171 3689 9180 3723
rect 9128 3680 9180 3689
rect 9312 3680 9364 3732
rect 10876 3680 10928 3732
rect 11060 3680 11112 3732
rect 12348 3680 12400 3732
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 13820 3723 13872 3732
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 15752 3723 15804 3732
rect 13820 3680 13872 3689
rect 15752 3689 15761 3723
rect 15761 3689 15795 3723
rect 15795 3689 15804 3723
rect 15752 3680 15804 3689
rect 19248 3680 19300 3732
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 9864 3655 9916 3664
rect 9864 3621 9873 3655
rect 9873 3621 9907 3655
rect 9907 3621 9916 3655
rect 9864 3612 9916 3621
rect 10784 3612 10836 3664
rect 15660 3612 15712 3664
rect 18144 3612 18196 3664
rect 21732 3655 21784 3664
rect 11060 3544 11112 3596
rect 11336 3544 11388 3596
rect 11704 3587 11756 3596
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 13360 3544 13412 3596
rect 14280 3544 14332 3596
rect 16120 3544 16172 3596
rect 17040 3587 17092 3596
rect 17040 3553 17049 3587
rect 17049 3553 17083 3587
rect 17083 3553 17092 3587
rect 17040 3544 17092 3553
rect 17132 3544 17184 3596
rect 17684 3544 17736 3596
rect 4712 3451 4764 3460
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2412 3340 2464 3392
rect 4712 3417 4721 3451
rect 4721 3417 4755 3451
rect 4755 3417 4764 3451
rect 4712 3408 4764 3417
rect 5264 3408 5316 3460
rect 7840 3451 7892 3460
rect 7840 3417 7849 3451
rect 7849 3417 7883 3451
rect 7883 3417 7892 3451
rect 7840 3408 7892 3417
rect 7932 3408 7984 3460
rect 10140 3408 10192 3460
rect 12716 3408 12768 3460
rect 13728 3408 13780 3460
rect 17960 3544 18012 3596
rect 15384 3451 15436 3460
rect 15384 3417 15393 3451
rect 15393 3417 15427 3451
rect 15427 3417 15436 3451
rect 15384 3408 15436 3417
rect 15936 3408 15988 3460
rect 17408 3408 17460 3460
rect 18788 3544 18840 3596
rect 21732 3621 21741 3655
rect 21741 3621 21775 3655
rect 21775 3621 21784 3655
rect 21732 3612 21784 3621
rect 21824 3655 21876 3664
rect 21824 3621 21833 3655
rect 21833 3621 21867 3655
rect 21867 3621 21876 3655
rect 21824 3612 21876 3621
rect 22100 3612 22152 3664
rect 22836 3612 22888 3664
rect 24124 3655 24176 3664
rect 24124 3621 24133 3655
rect 24133 3621 24167 3655
rect 24167 3621 24176 3655
rect 24124 3612 24176 3621
rect 24768 3612 24820 3664
rect 22008 3519 22060 3528
rect 22008 3485 22017 3519
rect 22017 3485 22051 3519
rect 22051 3485 22060 3519
rect 22008 3476 22060 3485
rect 23204 3476 23256 3528
rect 18420 3451 18472 3460
rect 18420 3417 18429 3451
rect 18429 3417 18463 3451
rect 18463 3417 18472 3451
rect 18420 3408 18472 3417
rect 20536 3408 20588 3460
rect 7656 3340 7708 3392
rect 14832 3383 14884 3392
rect 14832 3349 14841 3383
rect 14841 3349 14875 3383
rect 14875 3349 14884 3383
rect 14832 3340 14884 3349
rect 18788 3383 18840 3392
rect 18788 3349 18797 3383
rect 18797 3349 18831 3383
rect 18831 3349 18840 3383
rect 18788 3340 18840 3349
rect 19432 3340 19484 3392
rect 20444 3383 20496 3392
rect 20444 3349 20453 3383
rect 20453 3349 20487 3383
rect 20487 3349 20496 3383
rect 20444 3340 20496 3349
rect 23756 3383 23808 3392
rect 23756 3349 23765 3383
rect 23765 3349 23799 3383
rect 23799 3349 23808 3383
rect 23756 3340 23808 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1400 3136 1452 3188
rect 2688 3136 2740 3188
rect 3608 3179 3660 3188
rect 2136 3111 2188 3120
rect 2136 3077 2145 3111
rect 2145 3077 2179 3111
rect 2179 3077 2188 3111
rect 2136 3068 2188 3077
rect 3608 3145 3617 3179
rect 3617 3145 3651 3179
rect 3651 3145 3660 3179
rect 3608 3136 3660 3145
rect 5080 3179 5132 3188
rect 5080 3145 5089 3179
rect 5089 3145 5123 3179
rect 5123 3145 5132 3179
rect 5080 3136 5132 3145
rect 6460 3136 6512 3188
rect 7564 3136 7616 3188
rect 8208 3136 8260 3188
rect 9864 3136 9916 3188
rect 11060 3136 11112 3188
rect 13360 3136 13412 3188
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 21364 3179 21416 3188
rect 14188 3136 14240 3145
rect 5540 3111 5592 3120
rect 5540 3077 5549 3111
rect 5549 3077 5583 3111
rect 5583 3077 5592 3111
rect 5540 3068 5592 3077
rect 6368 3068 6420 3120
rect 7748 3068 7800 3120
rect 11796 3111 11848 3120
rect 3148 3000 3200 3052
rect 3792 2975 3844 2984
rect 3792 2941 3801 2975
rect 3801 2941 3835 2975
rect 3835 2941 3844 2975
rect 6736 3000 6788 3052
rect 3792 2932 3844 2941
rect 6460 2932 6512 2984
rect 2412 2907 2464 2916
rect 2412 2873 2421 2907
rect 2421 2873 2455 2907
rect 2455 2873 2464 2907
rect 2412 2864 2464 2873
rect 3608 2864 3660 2916
rect 5172 2864 5224 2916
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 14280 3068 14332 3120
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 21732 3136 21784 3188
rect 23204 3136 23256 3188
rect 9128 3000 9180 3052
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 12348 2932 12400 2984
rect 17040 3068 17092 3120
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 15568 3000 15620 3052
rect 16580 3000 16632 3052
rect 17776 3043 17828 3052
rect 17776 3009 17785 3043
rect 17785 3009 17819 3043
rect 17819 3009 17828 3043
rect 17776 3000 17828 3009
rect 15016 2975 15068 2984
rect 9772 2864 9824 2916
rect 3424 2796 3476 2848
rect 3976 2796 4028 2848
rect 12808 2864 12860 2916
rect 15016 2941 15025 2975
rect 15025 2941 15059 2975
rect 15059 2941 15068 2975
rect 15016 2932 15068 2941
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 21824 3000 21876 3052
rect 22560 3000 22612 3052
rect 16304 2864 16356 2916
rect 16856 2864 16908 2916
rect 17132 2907 17184 2916
rect 17132 2873 17141 2907
rect 17141 2873 17175 2907
rect 17175 2873 17184 2907
rect 17132 2864 17184 2873
rect 17684 2864 17736 2916
rect 18788 2932 18840 2984
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 12532 2839 12584 2848
rect 12532 2805 12541 2839
rect 12541 2805 12575 2839
rect 12575 2805 12584 2839
rect 12532 2796 12584 2805
rect 13728 2796 13780 2848
rect 15936 2796 15988 2848
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 17776 2796 17828 2848
rect 18880 2864 18932 2916
rect 20996 2932 21048 2984
rect 23756 2975 23808 2984
rect 23756 2941 23765 2975
rect 23765 2941 23799 2975
rect 23799 2941 23808 2975
rect 23756 2932 23808 2941
rect 24124 3000 24176 3052
rect 18788 2796 18840 2848
rect 20720 2864 20772 2916
rect 21732 2796 21784 2848
rect 27528 2796 27580 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2320 2592 2372 2644
rect 3424 2635 3476 2644
rect 2688 2524 2740 2576
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 4160 2592 4212 2644
rect 4988 2592 5040 2644
rect 7840 2592 7892 2644
rect 3976 2524 4028 2576
rect 7748 2567 7800 2576
rect 7748 2533 7757 2567
rect 7757 2533 7791 2567
rect 7791 2533 7800 2567
rect 7748 2524 7800 2533
rect 1952 2456 2004 2508
rect 3884 2388 3936 2440
rect 4160 2431 4212 2440
rect 4160 2397 4169 2431
rect 4169 2397 4203 2431
rect 4203 2397 4212 2431
rect 4160 2388 4212 2397
rect 4712 2363 4764 2372
rect 4712 2329 4721 2363
rect 4721 2329 4755 2363
rect 4755 2329 4764 2363
rect 4712 2320 4764 2329
rect 7288 2456 7340 2508
rect 12532 2592 12584 2644
rect 15016 2592 15068 2644
rect 16672 2592 16724 2644
rect 17684 2635 17736 2644
rect 9864 2524 9916 2576
rect 10968 2567 11020 2576
rect 10968 2533 10977 2567
rect 10977 2533 11011 2567
rect 11011 2533 11020 2567
rect 10968 2524 11020 2533
rect 11336 2567 11388 2576
rect 11336 2533 11345 2567
rect 11345 2533 11379 2567
rect 11379 2533 11388 2567
rect 11336 2524 11388 2533
rect 12072 2524 12124 2576
rect 9772 2456 9824 2508
rect 14372 2524 14424 2576
rect 15200 2567 15252 2576
rect 15200 2533 15209 2567
rect 15209 2533 15243 2567
rect 15243 2533 15252 2567
rect 15200 2524 15252 2533
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 18972 2592 19024 2644
rect 20628 2592 20680 2644
rect 22652 2635 22704 2644
rect 21364 2567 21416 2576
rect 21364 2533 21373 2567
rect 21373 2533 21407 2567
rect 21407 2533 21416 2567
rect 21364 2524 21416 2533
rect 22652 2601 22661 2635
rect 22661 2601 22695 2635
rect 22695 2601 22704 2635
rect 22652 2592 22704 2601
rect 22836 2592 22888 2644
rect 26148 2635 26200 2644
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 11704 2320 11756 2372
rect 12072 2320 12124 2372
rect 18420 2456 18472 2508
rect 20628 2456 20680 2508
rect 14188 2431 14240 2440
rect 14188 2397 14197 2431
rect 14197 2397 14231 2431
rect 14231 2397 14240 2431
rect 14188 2388 14240 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 26148 2601 26157 2635
rect 26157 2601 26191 2635
rect 26191 2601 26200 2635
rect 26148 2592 26200 2601
rect 16304 2320 16356 2372
rect 16856 2320 16908 2372
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 3884 2252 3936 2304
rect 4988 2252 5040 2304
rect 6000 2295 6052 2304
rect 6000 2261 6009 2295
rect 6009 2261 6043 2295
rect 6043 2261 6052 2295
rect 6000 2252 6052 2261
rect 14740 2252 14792 2304
rect 15752 2295 15804 2304
rect 15752 2261 15761 2295
rect 15761 2261 15795 2295
rect 15795 2261 15804 2295
rect 15752 2252 15804 2261
rect 19340 2252 19392 2304
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 20812 2252 20864 2304
rect 26608 2320 26660 2372
rect 24676 2252 24728 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 2596 2048 2648 2100
rect 2964 2048 3016 2100
rect 7288 2048 7340 2100
rect 10692 2048 10744 2100
rect 19340 2048 19392 2100
rect 8484 76 8536 128
rect 9128 76 9180 128
rect 15752 76 15804 128
rect 19708 76 19760 128
<< metal2 >>
rect 1582 26888 1638 26897
rect 1582 26823 1638 26832
rect 24766 26888 24822 26897
rect 24766 26823 24822 26832
rect 1030 25800 1086 25809
rect 1030 25735 1086 25744
rect 110 20088 166 20097
rect 166 20046 244 20074
rect 110 20023 166 20032
rect 216 19334 244 20046
rect 216 19306 428 19334
rect 296 18148 348 18154
rect 296 18090 348 18096
rect 112 17128 164 17134
rect 112 17070 164 17076
rect 20 15632 72 15638
rect 20 15574 72 15580
rect 32 4154 60 15574
rect 124 6633 152 17070
rect 204 13728 256 13734
rect 204 13670 256 13676
rect 110 6624 166 6633
rect 110 6559 166 6568
rect 110 5672 166 5681
rect 216 5658 244 13670
rect 308 8265 336 18090
rect 400 11082 428 19306
rect 940 18216 992 18222
rect 940 18158 992 18164
rect 952 17785 980 18158
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 1044 16794 1072 25735
rect 1490 24032 1546 24041
rect 1490 23967 1546 23976
rect 1124 21480 1176 21486
rect 1124 21422 1176 21428
rect 1136 18358 1164 21422
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1308 19916 1360 19922
rect 1308 19858 1360 19864
rect 1320 19825 1348 19858
rect 1306 19816 1362 19825
rect 1306 19751 1362 19760
rect 1308 19712 1360 19718
rect 1308 19654 1360 19660
rect 1216 18828 1268 18834
rect 1216 18770 1268 18776
rect 1124 18352 1176 18358
rect 1124 18294 1176 18300
rect 1228 18154 1256 18770
rect 1216 18148 1268 18154
rect 1216 18090 1268 18096
rect 1124 18080 1176 18086
rect 1124 18022 1176 18028
rect 1032 16788 1084 16794
rect 1032 16730 1084 16736
rect 478 12200 534 12209
rect 478 12135 534 12144
rect 388 11076 440 11082
rect 388 11018 440 11024
rect 386 10840 442 10849
rect 492 10826 520 12135
rect 1136 11336 1164 18022
rect 1216 14612 1268 14618
rect 1216 14554 1268 14560
rect 1228 11558 1256 14554
rect 1320 13530 1348 19654
rect 1412 18465 1440 20334
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1400 18352 1452 18358
rect 1400 18294 1452 18300
rect 1308 13524 1360 13530
rect 1308 13466 1360 13472
rect 1320 12850 1348 13466
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1306 11792 1362 11801
rect 1306 11727 1362 11736
rect 1216 11552 1268 11558
rect 1216 11494 1268 11500
rect 1136 11308 1256 11336
rect 1122 11248 1178 11257
rect 1122 11183 1178 11192
rect 442 10798 520 10826
rect 386 10775 442 10784
rect 294 8256 350 8265
rect 294 8191 350 8200
rect 1136 5778 1164 11183
rect 1228 6730 1256 11308
rect 1320 8650 1348 11727
rect 1412 10266 1440 18294
rect 1504 16250 1532 23967
rect 1596 23866 1624 26823
rect 24214 25800 24270 25809
rect 24214 25735 24270 25744
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 1674 24848 1730 24857
rect 1674 24783 1730 24792
rect 23938 24848 23994 24857
rect 23938 24783 23994 24792
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1596 21690 1624 22607
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1582 18592 1638 18601
rect 1582 18527 1638 18536
rect 1596 17882 1624 18527
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1492 16244 1544 16250
rect 1492 16186 1544 16192
rect 1492 15972 1544 15978
rect 1492 15914 1544 15920
rect 1504 15586 1532 15914
rect 1596 15706 1624 16594
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1504 15558 1624 15586
rect 1492 15428 1544 15434
rect 1492 15370 1544 15376
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1320 8622 1440 8650
rect 1308 8560 1360 8566
rect 1308 8502 1360 8508
rect 1216 6724 1268 6730
rect 1216 6666 1268 6672
rect 1124 5772 1176 5778
rect 1124 5714 1176 5720
rect 166 5630 244 5658
rect 110 5607 166 5616
rect 1136 5370 1164 5714
rect 1124 5364 1176 5370
rect 1124 5306 1176 5312
rect 32 4126 152 4154
rect 20 3664 72 3670
rect 20 3606 72 3612
rect 32 3505 60 3606
rect 18 3496 74 3505
rect 18 3431 74 3440
rect 124 82 152 4126
rect 478 82 534 480
rect 124 54 534 82
rect 1320 82 1348 8502
rect 1412 3602 1440 8622
rect 1504 5137 1532 15370
rect 1490 5128 1546 5137
rect 1490 5063 1546 5072
rect 1596 3670 1624 15558
rect 1688 14074 1716 24783
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 23480 23656 23532 23662
rect 23480 23598 23532 23604
rect 2136 23520 2188 23526
rect 2136 23462 2188 23468
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1768 18624 1820 18630
rect 1768 18566 1820 18572
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1780 13814 1808 18566
rect 1872 17649 1900 19246
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1858 17640 1914 17649
rect 1858 17575 1914 17584
rect 1964 16697 1992 19110
rect 1950 16688 2006 16697
rect 1950 16623 2006 16632
rect 2056 16436 2084 19382
rect 1688 13786 1808 13814
rect 1872 16408 2084 16436
rect 1688 9722 1716 13786
rect 1872 12442 1900 16408
rect 2148 16250 2176 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2240 19514 2268 19858
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 2228 19508 2280 19514
rect 2228 19450 2280 19456
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2240 18222 2268 18770
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2056 15570 2084 15642
rect 2044 15564 2096 15570
rect 1964 15524 2044 15552
rect 1964 14618 1992 15524
rect 2044 15506 2096 15512
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2134 14784 2190 14793
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 13530 2084 14758
rect 2134 14719 2190 14728
rect 2148 14074 2176 14719
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1780 11014 1808 11222
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10538 1808 10950
rect 1872 10674 1900 12378
rect 1964 11762 1992 12378
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10532 1820 10538
rect 1768 10474 1820 10480
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1964 9654 1992 9862
rect 1952 9648 2004 9654
rect 1766 9616 1822 9625
rect 1952 9590 2004 9596
rect 1766 9551 1822 9560
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 8090 1716 9318
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1688 7410 1716 8026
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1688 6458 1716 6938
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1780 4690 1808 9551
rect 1964 9518 1992 9590
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 2056 9466 2084 12922
rect 2148 12832 2176 13874
rect 2240 12986 2268 18158
rect 2332 17746 2360 18566
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 2332 17338 2360 17682
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 2596 16652 2648 16658
rect 2596 16594 2648 16600
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2228 12980 2280 12986
rect 2228 12922 2280 12928
rect 2148 12804 2268 12832
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2148 12374 2176 12650
rect 2136 12368 2188 12374
rect 2136 12310 2188 12316
rect 2148 11898 2176 12310
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2056 9438 2176 9466
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 1860 9104 1912 9110
rect 1860 9046 1912 9052
rect 1872 8294 1900 9046
rect 1964 8838 1992 9318
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1872 7274 1900 8230
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1872 5370 1900 7210
rect 1964 6089 1992 8774
rect 2056 6934 2084 9318
rect 2148 7206 2176 9438
rect 2136 7200 2188 7206
rect 2136 7142 2188 7148
rect 2044 6928 2096 6934
rect 2044 6870 2096 6876
rect 2056 6458 2084 6870
rect 2136 6792 2188 6798
rect 2240 6780 2268 12804
rect 2332 12442 2360 15438
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2332 11354 2360 12174
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2332 10266 2360 11086
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 9110 2360 10066
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2332 8498 2360 9046
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2332 7818 2360 8298
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2332 6798 2360 7754
rect 2188 6752 2268 6780
rect 2136 6734 2188 6740
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1950 6080 2006 6089
rect 1950 6015 2006 6024
rect 2240 5914 2268 6752
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2228 5908 2280 5914
rect 2228 5850 2280 5856
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1872 5098 1900 5306
rect 2148 5234 2176 5510
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1860 5092 1912 5098
rect 1860 5034 1912 5040
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1780 4214 1808 4626
rect 1768 4208 1820 4214
rect 1768 4150 1820 4156
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1584 3664 1636 3670
rect 1584 3606 1636 3612
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1412 3194 1440 3538
rect 1584 3528 1636 3534
rect 1584 3470 1636 3476
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1596 2650 1624 3470
rect 1872 3398 1900 4014
rect 2148 3913 2176 5170
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2240 4214 2268 5034
rect 2228 4208 2280 4214
rect 2228 4154 2280 4156
rect 2228 4150 2360 4154
rect 2240 4146 2360 4150
rect 2240 4140 2372 4146
rect 2240 4126 2320 4140
rect 2320 4082 2372 4088
rect 2320 3936 2372 3942
rect 2134 3904 2190 3913
rect 2320 3878 2372 3884
rect 2134 3839 2190 3848
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1872 1057 1900 3334
rect 2134 3224 2190 3233
rect 2134 3159 2190 3168
rect 2148 3126 2176 3159
rect 2136 3120 2188 3126
rect 2136 3062 2188 3068
rect 2332 2650 2360 3878
rect 2424 3738 2452 15846
rect 2516 13530 2544 16390
rect 2608 16028 2636 16594
rect 2688 16040 2740 16046
rect 2608 16000 2688 16028
rect 2688 15982 2740 15988
rect 2700 15638 2728 15982
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2608 13870 2636 14486
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2516 10198 2544 13330
rect 2608 12918 2636 13806
rect 2700 13802 2728 14350
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2700 13190 2728 13738
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2596 12232 2648 12238
rect 2700 12220 2728 13126
rect 2648 12192 2728 12220
rect 2596 12174 2648 12180
rect 2608 10674 2636 12174
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2516 9178 2544 10134
rect 2596 9444 2648 9450
rect 2596 9386 2648 9392
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2504 8016 2556 8022
rect 2608 8004 2636 9386
rect 2700 9382 2728 10134
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2700 8362 2728 8774
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2792 8265 2820 18022
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 16425 2912 17070
rect 2870 16416 2926 16425
rect 2870 16351 2926 16360
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2884 15162 2912 15506
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2884 14958 2912 15098
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14618 2912 14894
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2884 12646 2912 14282
rect 2976 13938 3004 17478
rect 3068 16998 3096 17682
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3068 15502 3096 16934
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3068 14346 3096 15302
rect 3056 14340 3108 14346
rect 3056 14282 3108 14288
rect 3160 14226 3188 17002
rect 3068 14198 3188 14226
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2964 11620 3016 11626
rect 2964 11562 3016 11568
rect 2976 10810 3004 11562
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2976 10538 3004 10746
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2872 8968 2924 8974
rect 3068 8956 3096 14198
rect 3148 13796 3200 13802
rect 3148 13738 3200 13744
rect 3160 13530 3188 13738
rect 3252 13734 3280 19110
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 4344 18148 4396 18154
rect 4344 18090 4396 18096
rect 7288 18148 7340 18154
rect 7288 18090 7340 18096
rect 3424 18080 3476 18086
rect 4356 18057 4384 18090
rect 6828 18080 6880 18086
rect 3424 18022 3476 18028
rect 4342 18048 4398 18057
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 9926 3188 13262
rect 3252 12986 3280 13398
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 2872 8910 2924 8916
rect 2976 8928 3096 8956
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2884 8090 2912 8910
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2556 7976 2636 8004
rect 2504 7958 2556 7964
rect 2608 7546 2636 7976
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2608 7002 2636 7482
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2516 6322 2544 6666
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2608 6186 2636 6938
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 4826 2544 5646
rect 2700 5098 2728 5782
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2608 4758 2636 4966
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2700 3670 2728 5034
rect 2688 3664 2740 3670
rect 2688 3606 2740 3612
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 2424 2922 2452 3334
rect 2700 3194 2728 3606
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2700 2582 2728 3130
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1964 2310 1992 2450
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 1601 1992 2246
rect 2976 2106 3004 8928
rect 3160 8022 3188 9658
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 6322 3096 6666
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 5234 3096 5578
rect 3160 5302 3188 7142
rect 3252 6458 3280 12582
rect 3344 9586 3372 16390
rect 3436 11150 3464 18022
rect 7300 18057 7328 18090
rect 6828 18022 6880 18028
rect 7286 18048 7342 18057
rect 4342 17983 4398 17992
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3516 14476 3568 14482
rect 3516 14418 3568 14424
rect 3528 13530 3556 14418
rect 3516 13524 3568 13530
rect 3516 13466 3568 13472
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3528 12442 3556 13262
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3514 12336 3570 12345
rect 3514 12271 3570 12280
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3436 9586 3464 9998
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3344 9178 3372 9522
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3528 8906 3556 12271
rect 3620 10674 3648 14758
rect 3712 13258 3740 16934
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 12442 3740 12786
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3700 12300 3752 12306
rect 3700 12242 3752 12248
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3620 10266 3648 10610
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9178 3648 9862
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3712 7562 3740 12242
rect 3804 11762 3832 17478
rect 3988 17066 4016 17682
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 3976 17060 4028 17066
rect 3976 17002 4028 17008
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4160 16176 4212 16182
rect 4160 16118 4212 16124
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3884 15904 3936 15910
rect 3988 15881 4016 15914
rect 3884 15846 3936 15852
rect 3974 15872 4030 15881
rect 3896 13394 3924 15846
rect 3974 15807 4030 15816
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 11354 3832 11698
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11200 3924 13194
rect 3988 12850 4016 13738
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3988 11762 4016 12786
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11286 4016 11698
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 3804 11172 3924 11200
rect 3804 10198 3832 11172
rect 4080 11132 4108 15370
rect 4172 14482 4200 16118
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 14822 4292 15506
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4172 13734 4200 14418
rect 4160 13728 4212 13734
rect 4160 13670 4212 13676
rect 4172 13433 4200 13670
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 4264 13326 4292 14758
rect 4356 13938 4384 15982
rect 4448 15910 4476 16594
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4342 13832 4398 13841
rect 4342 13767 4398 13776
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4172 12714 4200 12922
rect 4160 12708 4212 12714
rect 4160 12650 4212 12656
rect 4172 11830 4200 12650
rect 4250 12472 4306 12481
rect 4250 12407 4306 12416
rect 4264 12170 4292 12407
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3896 11104 4108 11132
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3804 9722 3832 10134
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3896 9518 3924 11104
rect 4172 10538 4200 11222
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 4264 9024 4292 11698
rect 4080 8996 4292 9024
rect 4080 8566 4108 8996
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 4356 8480 4384 13767
rect 4448 11762 4476 15846
rect 4632 14793 4660 17138
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4618 14784 4674 14793
rect 4618 14719 4674 14728
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4436 10192 4488 10198
rect 4436 10134 4488 10140
rect 4448 9382 4476 10134
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4172 8452 4384 8480
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3804 7886 3832 8230
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3344 7534 3740 7562
rect 3804 7546 3832 7822
rect 3988 7546 4016 7958
rect 3792 7540 3844 7546
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3160 4758 3188 5238
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3160 3670 3188 4558
rect 3344 4154 3372 7534
rect 3792 7482 3844 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3620 7002 3648 7346
rect 4080 7274 4108 8230
rect 4068 7268 4120 7274
rect 4068 7210 4120 7216
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 4214 3464 6054
rect 3988 4758 4016 6598
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4080 5234 4108 6258
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 3976 4752 4028 4758
rect 3976 4694 4028 4700
rect 3988 4282 4016 4694
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3252 4126 3372 4154
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3160 3058 3188 3606
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2596 2100 2648 2106
rect 2596 2042 2648 2048
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 1950 1592 2006 1601
rect 1950 1527 2006 1536
rect 1858 1048 1914 1057
rect 1858 983 1914 992
rect 1398 82 1454 480
rect 1320 54 1454 82
rect 478 0 534 54
rect 1398 0 1454 54
rect 2318 82 2374 480
rect 2608 82 2636 2042
rect 2318 54 2636 82
rect 3252 82 3280 4126
rect 3436 2854 3464 4150
rect 3608 4004 3660 4010
rect 3608 3946 3660 3952
rect 3620 3194 3648 3946
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3641 3832 3878
rect 4172 3670 4200 8452
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7886 4384 8298
rect 4448 8022 4476 9318
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4540 7410 4568 14214
rect 4632 13802 4660 14214
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10470 4660 11154
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4632 9625 4660 10406
rect 4618 9616 4674 9625
rect 4618 9551 4674 9560
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4632 8634 4660 8978
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 6934 4568 7142
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4620 6792 4672 6798
rect 4724 6780 4752 16934
rect 4816 10742 4844 16934
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4908 14822 4936 15506
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4908 9330 4936 14758
rect 5000 13394 5028 14758
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12986 5028 13330
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4986 12336 5042 12345
rect 4986 12271 4988 12280
rect 5040 12271 5042 12280
rect 4988 12242 5040 12248
rect 5000 11558 5028 12242
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 5000 10713 5028 11494
rect 5092 11354 5120 17478
rect 5276 16998 5304 17682
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6368 17264 6420 17270
rect 6368 17206 6420 17212
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5184 14618 5212 14894
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5184 14074 5212 14350
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5184 13530 5212 13738
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5184 12986 5212 13330
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4986 10704 5042 10713
rect 5092 10674 5120 11290
rect 5184 10674 5212 12582
rect 4986 10639 5042 10648
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5170 10160 5226 10169
rect 5170 10095 5226 10104
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4816 9302 4936 9330
rect 4816 7342 4844 9302
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4908 7818 4936 9114
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4672 6752 4752 6780
rect 4620 6734 4672 6740
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4264 5370 4292 5714
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4160 3664 4212 3670
rect 3790 3632 3846 3641
rect 4160 3606 4212 3612
rect 3790 3567 3846 3576
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3620 2922 3648 3130
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3436 2650 3464 2790
rect 3804 2650 3832 2926
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3988 2582 4016 2790
rect 4160 2644 4212 2650
rect 4160 2586 4212 2592
rect 3976 2576 4028 2582
rect 3976 2518 4028 2524
rect 4172 2446 4200 2586
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 3896 2310 3924 2382
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3330 82 3386 480
rect 3252 54 3386 82
rect 2318 0 2374 54
rect 3330 0 3386 54
rect 4250 82 4306 480
rect 4356 82 4384 6598
rect 4434 6080 4490 6089
rect 4434 6015 4490 6024
rect 4448 5914 4476 6015
rect 4724 5914 4752 6752
rect 4908 6458 4936 6870
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4448 4536 4476 5850
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4540 5001 4568 5034
rect 4526 4992 4582 5001
rect 4526 4927 4582 4936
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4528 4548 4580 4554
rect 4448 4508 4528 4536
rect 4528 4490 4580 4496
rect 4436 4072 4488 4078
rect 4632 4060 4660 4694
rect 4488 4032 4660 4060
rect 4436 4014 4488 4020
rect 4448 3670 4476 4014
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4724 2378 4752 3402
rect 5000 2650 5028 9454
rect 5092 9178 5120 9522
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5184 9042 5212 10095
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 7954 5120 8230
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5172 7744 5224 7750
rect 5172 7686 5224 7692
rect 5184 7274 5212 7686
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5276 4154 5304 16934
rect 5368 12918 5396 16934
rect 6196 16726 6224 16934
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15366 5580 15846
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 14940 5580 15302
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5632 14952 5684 14958
rect 5552 14912 5632 14940
rect 5632 14894 5684 14900
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12306 5396 12650
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5460 11218 5488 14554
rect 5644 14482 5672 14894
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5552 13938 5580 14418
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5644 13814 5672 13942
rect 6012 13841 6040 16458
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 5552 13786 5672 13814
rect 5998 13832 6054 13841
rect 5552 12850 5580 13786
rect 5998 13767 6054 13776
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 6012 12374 6040 12922
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11898 5580 12174
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11898 6040 12310
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6012 11286 6040 11834
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 6012 10538 6040 11222
rect 6104 11014 6132 16390
rect 6196 16153 6224 16662
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6182 16144 6238 16153
rect 6288 16114 6316 16594
rect 6182 16079 6238 16088
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6288 16017 6316 16050
rect 6274 16008 6330 16017
rect 6274 15943 6330 15952
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6196 14006 6224 14826
rect 6274 14512 6330 14521
rect 6274 14447 6330 14456
rect 6288 14113 6316 14447
rect 6274 14104 6330 14113
rect 6274 14039 6330 14048
rect 6184 14000 6236 14006
rect 6184 13942 6236 13948
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 6196 10690 6224 13942
rect 6288 11898 6316 14039
rect 6380 11914 6408 17206
rect 6748 16998 6776 17682
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6472 15162 6500 15506
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6472 14822 6500 14962
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 12050 6500 14758
rect 6564 12170 6592 15846
rect 6656 15570 6684 16390
rect 6644 15564 6696 15570
rect 6644 15506 6696 15512
rect 6656 14618 6684 15506
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 12646 6684 13738
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6748 12170 6776 16934
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6472 12022 6776 12050
rect 6276 11892 6328 11898
rect 6380 11886 6592 11914
rect 6276 11834 6328 11840
rect 6288 11694 6316 11834
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6380 11626 6408 11766
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6380 11354 6408 11562
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6368 11348 6420 11354
rect 6368 11290 6420 11296
rect 6472 11150 6500 11494
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6104 10662 6224 10690
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9450 5396 9862
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 5368 9178 5396 9386
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 9042 5488 10202
rect 6104 10198 6132 10662
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 6012 9722 6040 10066
rect 6104 9722 6132 10134
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5460 8634 5488 8978
rect 5920 8974 5948 9386
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 8022 5396 8298
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7750 5396 7958
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5460 6730 5488 8434
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 8022 5672 8230
rect 6012 8022 6040 9046
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 7002 5672 7142
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5448 6724 5500 6730
rect 5448 6666 5500 6672
rect 5552 6458 5580 6802
rect 5920 6644 5948 7346
rect 6012 7002 6040 7822
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5920 6616 6040 6644
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5368 5098 5396 5510
rect 5356 5092 5408 5098
rect 5356 5034 5408 5040
rect 5368 4826 5396 5034
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5184 4126 5304 4154
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5092 3194 5120 3674
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5184 2922 5212 4126
rect 5368 4010 5396 4422
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5276 3466 5304 3946
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5172 2916 5224 2922
rect 5172 2858 5224 2864
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4712 2372 4764 2378
rect 4712 2314 4764 2320
rect 5000 2310 5028 2586
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4250 54 4384 82
rect 5184 82 5212 2858
rect 5460 1873 5488 5578
rect 5552 4826 5580 5646
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 4706 5672 5238
rect 6012 5098 6040 6616
rect 6104 6458 6132 9658
rect 6196 6662 6224 10542
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5908 4820 5960 4826
rect 5960 4780 6040 4808
rect 5908 4762 5960 4768
rect 5552 4678 5672 4706
rect 5552 4146 5580 4678
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 6012 3641 6040 4780
rect 5998 3632 6054 3641
rect 5540 3596 5592 3602
rect 5998 3567 6054 3576
rect 5540 3538 5592 3544
rect 5552 3126 5580 3538
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5446 1864 5502 1873
rect 5446 1799 5502 1808
rect 6012 1465 6040 2246
rect 5998 1456 6054 1465
rect 5998 1391 6054 1400
rect 5262 82 5318 480
rect 5184 54 5318 82
rect 4250 0 4306 54
rect 5262 0 5318 54
rect 6182 82 6238 480
rect 6288 82 6316 7278
rect 6380 5370 6408 11018
rect 6458 9616 6514 9625
rect 6458 9551 6514 9560
rect 6472 8537 6500 9551
rect 6458 8528 6514 8537
rect 6458 8463 6514 8472
rect 6564 8294 6592 11886
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6656 8090 6684 9318
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6472 7206 6500 7958
rect 6748 7410 6776 12022
rect 6840 11830 6868 18022
rect 7286 17983 7342 17992
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 13452 17740 13504 17746
rect 13452 17682 13504 17688
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7116 15910 7144 16594
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 12238 6960 13670
rect 7024 12850 7052 15438
rect 7116 13512 7144 15846
rect 7208 13682 7236 17478
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13870 7328 14214
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7208 13654 7328 13682
rect 7116 13484 7236 13512
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 12986 7144 13330
rect 7208 12986 7236 13484
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6840 11354 6868 11766
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8090 6868 8230
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6932 7886 6960 10950
rect 7024 8906 7052 12582
rect 7116 11762 7144 12650
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7300 10130 7328 13654
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9518 7328 10066
rect 7104 9512 7156 9518
rect 7104 9454 7156 9460
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6828 7268 6880 7274
rect 6828 7210 6880 7216
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6472 6934 6500 7142
rect 6460 6928 6512 6934
rect 6460 6870 6512 6876
rect 6472 6458 6500 6870
rect 6748 6730 6776 7210
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6840 6662 6868 7210
rect 7024 6866 7052 8026
rect 7116 7750 7144 9454
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 8498 7236 9386
rect 7300 9110 7328 9454
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7300 8022 7328 9046
rect 7392 9042 7420 16934
rect 7668 16590 7696 16934
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7472 16040 7524 16046
rect 7472 15982 7524 15988
rect 7484 15026 7512 15982
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7392 8634 7420 8978
rect 7380 8628 7432 8634
rect 7380 8570 7432 8576
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 5846 6500 6394
rect 6840 6254 6868 6598
rect 7208 6254 7236 7822
rect 7300 7342 7328 7958
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6368 5024 6420 5030
rect 6472 5012 6500 5782
rect 6656 5137 6684 6054
rect 6642 5128 6698 5137
rect 6642 5063 6698 5072
rect 6420 4984 6500 5012
rect 6368 4966 6420 4972
rect 6472 4758 6500 4984
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6472 4214 6500 4694
rect 6460 4208 6512 4214
rect 6460 4154 6512 4156
rect 6380 4150 6512 4154
rect 6380 4126 6500 4150
rect 6380 3670 6408 4126
rect 6564 3738 6592 4966
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4078 6684 4558
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6380 3126 6408 3606
rect 6656 3505 6684 4014
rect 6642 3496 6698 3505
rect 6642 3431 6698 3440
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6368 3120 6420 3126
rect 6368 3062 6420 3068
rect 6472 2990 6500 3130
rect 6748 3058 6776 6054
rect 6840 5574 6868 6190
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6840 3534 6868 5510
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 6932 4826 6960 5034
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6840 3233 6868 3470
rect 6826 3224 6882 3233
rect 6826 3159 6882 3168
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6460 2984 6512 2990
rect 6458 2952 6460 2961
rect 6512 2952 6514 2961
rect 6458 2887 6514 2896
rect 6472 2861 6500 2887
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7300 2106 7328 2450
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 6182 54 6316 82
rect 7194 82 7250 480
rect 7392 82 7420 8570
rect 7484 5778 7512 14758
rect 7576 13546 7604 15030
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7668 13734 7696 13874
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7576 13518 7696 13546
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7576 12374 7604 12582
rect 7564 12368 7616 12374
rect 7564 12310 7616 12316
rect 7576 11354 7604 12310
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 11234 7696 13518
rect 7576 11206 7696 11234
rect 7760 11218 7788 16730
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7852 15978 7880 16594
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8220 16046 8248 16526
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 7840 15972 7892 15978
rect 7840 15914 7892 15920
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 8024 15904 8076 15910
rect 8024 15846 8076 15852
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7944 14958 7972 15642
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7944 13870 7972 14554
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7840 13728 7892 13734
rect 7944 13705 7972 13806
rect 7840 13670 7892 13676
rect 7930 13696 7986 13705
rect 7852 12322 7880 13670
rect 7930 13631 7986 13640
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12442 7972 13330
rect 7932 12436 7984 12442
rect 7932 12378 7984 12384
rect 7852 12294 7972 12322
rect 7748 11212 7800 11218
rect 7576 9586 7604 11206
rect 7748 11154 7800 11160
rect 7760 10266 7788 11154
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7668 9178 7696 9862
rect 7838 9344 7894 9353
rect 7838 9279 7894 9288
rect 7852 9178 7880 9279
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7746 9072 7802 9081
rect 7746 9007 7802 9016
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7668 7206 7696 7890
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7576 3194 7604 3470
rect 7668 3398 7696 7142
rect 7760 4214 7788 9007
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7852 6866 7880 8842
rect 7944 7954 7972 12294
rect 8036 10674 8064 15846
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 14890 8156 15506
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8312 14482 8340 15914
rect 8404 15570 8432 15982
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8404 14618 8432 15506
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8128 14074 8156 14418
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8312 13734 8340 14418
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8128 10198 8156 13126
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 8220 11898 8248 12310
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8312 11286 8340 12854
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8312 10810 8340 11222
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8312 10538 8340 10746
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8220 10198 8248 10406
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8128 9722 8156 10134
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8220 9586 8248 10134
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8312 8634 8340 9046
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8022 7168 8078 7177
rect 8022 7103 8078 7112
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 6118 7880 6802
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 4826 7880 5714
rect 8036 5370 8064 7103
rect 8128 6866 8156 7278
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8128 6458 8156 6802
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8404 6225 8432 12038
rect 8390 6216 8446 6225
rect 8390 6151 8446 6160
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7748 4004 7800 4010
rect 7800 3964 7880 3992
rect 7748 3946 7800 3952
rect 7852 3466 7880 3964
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7944 3466 7972 3878
rect 7840 3460 7892 3466
rect 7840 3402 7892 3408
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7760 2582 7788 3062
rect 7852 2650 7880 3402
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7194 54 7420 82
rect 8036 82 8064 5306
rect 8128 4758 8156 5578
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 4758 8248 5510
rect 8312 5001 8340 6054
rect 8298 4992 8354 5001
rect 8298 4927 8354 4936
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 8220 4282 8248 4694
rect 8312 4486 8340 4927
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8220 3194 8248 3606
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8114 82 8170 480
rect 8496 134 8524 12582
rect 8588 5234 8616 15438
rect 8680 10985 8708 17274
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 8772 13870 8800 17206
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9048 14550 9076 14758
rect 9036 14544 9088 14550
rect 9036 14486 9088 14492
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8864 13462 8892 13806
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 8864 12986 8892 13398
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12442 8892 12786
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8666 10976 8722 10985
rect 8666 10911 8722 10920
rect 8772 9110 8800 11630
rect 8864 10198 8892 12242
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8772 7274 8800 8230
rect 8864 7546 8892 9998
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8772 6186 8800 7210
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5846 8800 6122
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8588 4826 8616 5170
rect 8772 5030 8800 5782
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8772 4146 8800 4558
rect 8956 4154 8984 14350
rect 9048 14278 9076 14486
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13841 9076 14214
rect 9034 13832 9090 13841
rect 9034 13767 9090 13776
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 9048 11762 9076 13670
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 9722 9076 11494
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 9048 9450 9076 9658
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9048 7546 9076 9386
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 7274 9076 7482
rect 9140 7478 9168 16934
rect 9232 9586 9260 17070
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 9784 16046 9812 16594
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9312 15904 9364 15910
rect 9312 15846 9364 15852
rect 9324 13394 9352 15846
rect 9784 15638 9812 15982
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9312 13388 9364 13394
rect 9312 13330 9364 13336
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9324 12442 9352 12582
rect 9312 12436 9364 12442
rect 9312 12378 9364 12384
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 9324 11914 9352 12271
rect 9416 12220 9444 14758
rect 9692 14074 9720 14758
rect 9864 14544 9916 14550
rect 9864 14486 9916 14492
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9784 13920 9812 14350
rect 9600 13892 9812 13920
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 12345 9536 13670
rect 9600 13462 9628 13892
rect 9876 13530 9904 14486
rect 9968 13938 9996 16730
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 15910 10088 16526
rect 10888 16454 10916 17206
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16046 10916 16390
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10060 15094 10088 15846
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10140 15088 10192 15094
rect 10140 15030 10192 15036
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9954 13832 10010 13841
rect 9954 13767 10010 13776
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9494 12336 9550 12345
rect 9600 12306 9628 13398
rect 9494 12271 9550 12280
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9416 12192 9536 12220
rect 9324 11886 9444 11914
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 9178 9260 9522
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9232 7954 9260 8434
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9232 7857 9260 7890
rect 9218 7848 9274 7857
rect 9218 7783 9274 7792
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9140 7002 9168 7414
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5914 9168 6258
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9324 5710 9352 11766
rect 9416 10130 9444 11886
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4758 9352 4966
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9416 4154 9444 9862
rect 9508 6322 9536 12192
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9600 9722 9628 10066
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9692 6769 9720 12106
rect 9784 11082 9812 13398
rect 9968 12170 9996 13767
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10060 11558 10088 14894
rect 10152 13705 10180 15030
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10138 13696 10194 13705
rect 10138 13631 10194 13640
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10704 13462 10732 13738
rect 10784 13728 10836 13734
rect 10784 13670 10836 13676
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10152 12374 10180 13262
rect 10520 12986 10548 13262
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10704 12918 10732 13398
rect 10796 13190 10824 13670
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10796 12714 10824 13126
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10152 11898 10180 12310
rect 10704 12238 10732 12650
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10704 11762 10732 12174
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9876 9654 9904 11494
rect 10152 11354 10180 11698
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 10060 11014 10088 11222
rect 10704 11150 10732 11698
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10538 10088 10950
rect 10520 10810 10548 11086
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 10048 10532 10100 10538
rect 10048 10474 10100 10480
rect 9968 10062 9996 10474
rect 10152 10198 10180 10610
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10192 10192 10198
rect 10140 10134 10192 10140
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9784 7478 9812 8910
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9876 8022 9904 8570
rect 9968 8566 9996 8978
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9876 7546 9904 7958
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6792 9824 6798
rect 9678 6760 9734 6769
rect 9772 6734 9824 6740
rect 9678 6695 9734 6704
rect 9496 6316 9548 6322
rect 9496 6258 9548 6264
rect 9784 5914 9812 6734
rect 9876 6458 9904 6870
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 5370 9536 5714
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9784 5302 9812 5850
rect 9876 5370 9904 6258
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 9508 4214 9536 4558
rect 9784 4282 9812 4694
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 8760 4140 8812 4146
rect 8956 4126 9168 4154
rect 8760 4082 8812 4088
rect 8772 3670 8800 4082
rect 9140 3738 9168 4126
rect 9324 4126 9444 4154
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9772 4140 9824 4146
rect 9324 3738 9352 4126
rect 9772 4082 9824 4088
rect 9784 4010 9812 4082
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 9140 3058 9168 3674
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 9784 2922 9812 3946
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9876 3194 9904 3606
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 2916 9824 2922
rect 9772 2858 9824 2864
rect 9784 2514 9812 2858
rect 9876 2582 9904 3130
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 8036 54 8170 82
rect 8484 128 8536 134
rect 8484 70 8536 76
rect 9126 128 9182 480
rect 9126 76 9128 128
rect 9180 76 9182 128
rect 6182 0 6238 54
rect 7194 0 7250 54
rect 8114 0 8170 54
rect 9126 0 9182 76
rect 9968 82 9996 7958
rect 10060 7886 10088 9386
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8498 10732 8910
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10692 6792 10744 6798
rect 10796 6780 10824 11494
rect 10888 10146 10916 15982
rect 10980 15570 11008 17274
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10980 15162 11008 15506
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10980 14958 11008 15098
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10980 14618 11008 14894
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10980 12850 11008 14350
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 10980 12442 11008 12786
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 10888 10118 11008 10146
rect 10874 10024 10930 10033
rect 10874 9959 10930 9968
rect 10888 9926 10916 9959
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9586 10916 9862
rect 10980 9654 11008 10118
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 11072 9160 11100 16934
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11164 13326 11192 15438
rect 11256 13530 11284 15438
rect 11334 14648 11390 14657
rect 11334 14583 11390 14592
rect 11348 14414 11376 14583
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 13938 11376 14350
rect 11440 14074 11468 14486
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11256 11801 11284 13262
rect 11336 13184 11388 13190
rect 11336 13126 11388 13132
rect 11242 11792 11298 11801
rect 11348 11778 11376 13126
rect 11440 12374 11468 14010
rect 11428 12368 11480 12374
rect 11428 12310 11480 12316
rect 11440 11898 11468 12310
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11348 11750 11468 11778
rect 11242 11727 11298 11736
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 10198 11376 10474
rect 11336 10192 11388 10198
rect 11336 10134 11388 10140
rect 11348 9722 11376 10134
rect 11336 9716 11388 9722
rect 11336 9658 11388 9664
rect 11072 9132 11284 9160
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11072 8090 11100 8978
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8362 11192 8910
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11256 6780 11284 9132
rect 11336 6792 11388 6798
rect 10796 6752 10916 6780
rect 10692 6734 10744 6740
rect 10060 5642 10088 6734
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 5817 10180 6054
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5914 10732 6734
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10796 6322 10824 6598
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10796 5953 10824 6122
rect 10782 5944 10838 5953
rect 10692 5908 10744 5914
rect 10782 5879 10838 5888
rect 10692 5850 10744 5856
rect 10138 5808 10194 5817
rect 10138 5743 10194 5752
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10060 4622 10088 5578
rect 10152 5574 10180 5743
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5098 10364 5510
rect 10704 5234 10732 5850
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10796 4758 10824 5782
rect 10888 5778 10916 6752
rect 11256 6752 11336 6780
rect 11256 6390 11284 6752
rect 11336 6734 11388 6740
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10980 5692 11008 6122
rect 11072 6118 11100 6326
rect 11440 6236 11468 11750
rect 11532 11354 11560 15914
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11532 9586 11560 10134
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8634 11560 9046
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11532 7478 11560 8570
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11532 6458 11560 7210
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11624 6254 11652 17614
rect 13464 17338 13492 17682
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11716 14278 11744 15506
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 11830 11744 14214
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11808 11642 11836 17070
rect 11992 16250 12020 17070
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11886 13968 11942 13977
rect 11992 13938 12020 14350
rect 11886 13903 11942 13912
rect 11980 13932 12032 13938
rect 11900 12306 11928 13903
rect 11980 13874 12032 13880
rect 12084 13814 12112 16186
rect 12268 16114 12296 16390
rect 12728 16182 12756 16594
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12268 15434 12296 16050
rect 12624 16040 12676 16046
rect 12452 16000 12624 16028
rect 12452 15910 12480 16000
rect 12624 15982 12676 15988
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15570 12480 15846
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12268 14618 12296 15370
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12360 14550 12388 15506
rect 12452 14958 12480 15506
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 11992 13786 12112 13814
rect 11992 12617 12020 13786
rect 12164 13456 12216 13462
rect 12164 13398 12216 13404
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 12084 12646 12112 13330
rect 12176 12918 12204 13398
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12072 12640 12124 12646
rect 11978 12608 12034 12617
rect 12072 12582 12124 12588
rect 11978 12543 12034 12552
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11900 11898 11928 12242
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11716 11614 11836 11642
rect 11716 8090 11744 11614
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 7002 11744 7822
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11164 6208 11468 6236
rect 11612 6248 11664 6254
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11060 5704 11112 5710
rect 10980 5664 11060 5692
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10140 4140 10192 4146
rect 10888 4128 10916 5238
rect 10140 4082 10192 4088
rect 10796 4100 10916 4128
rect 10152 3942 10180 4082
rect 10324 4004 10376 4010
rect 10376 3964 10732 3992
rect 10324 3946 10376 3952
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10152 3058 10180 3402
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10336 1057 10364 2382
rect 10704 2106 10732 3964
rect 10796 3670 10824 4100
rect 10980 4010 11008 5664
rect 11060 5646 11112 5652
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 10796 3058 10824 3606
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10888 1601 10916 3674
rect 10980 2582 11008 3946
rect 11072 3738 11100 5510
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 11072 3194 11100 3538
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 10322 1048 10378 1057
rect 10322 983 10378 992
rect 10046 82 10102 480
rect 9968 54 10102 82
rect 10046 0 10102 54
rect 11058 82 11114 480
rect 11164 82 11192 6208
rect 11612 6190 11664 6196
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5846 11468 6054
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11440 5234 11468 5782
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11532 5370 11560 5714
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11256 3369 11284 4762
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4282 11376 4490
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11624 3641 11652 5034
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11716 4282 11744 4626
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11716 4010 11744 4218
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11610 3632 11666 3641
rect 11336 3596 11388 3602
rect 11716 3602 11744 3946
rect 11610 3567 11666 3576
rect 11704 3596 11756 3602
rect 11336 3538 11388 3544
rect 11704 3538 11756 3544
rect 11242 3360 11298 3369
rect 11242 3295 11298 3304
rect 11348 2582 11376 3538
rect 11808 3346 11836 11494
rect 11992 11218 12020 12543
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 10674 12020 11154
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11992 10577 12020 10610
rect 11978 10568 12034 10577
rect 11978 10503 12034 10512
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11900 8906 11928 9415
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 7818 11928 8298
rect 11992 8022 12020 8978
rect 11980 8016 12032 8022
rect 11980 7958 12032 7964
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11992 7546 12020 7958
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11716 3318 11836 3346
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11716 2378 11744 3318
rect 11794 3224 11850 3233
rect 11794 3159 11850 3168
rect 11808 3126 11836 3159
rect 11796 3120 11848 3126
rect 11900 3097 11928 6258
rect 11796 3062 11848 3068
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 12084 2961 12112 12582
rect 12268 11762 12296 14350
rect 12360 14074 12388 14486
rect 12728 14346 12756 16118
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12544 13938 12572 14214
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13530 12480 13670
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12256 11552 12308 11558
rect 12176 11512 12256 11540
rect 12176 5574 12204 11512
rect 12256 11494 12308 11500
rect 12360 10266 12388 12038
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9382 12296 9998
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8401 12296 9318
rect 12452 8945 12480 12106
rect 12544 10198 12572 13874
rect 12728 13734 12756 14282
rect 12820 14074 12848 14894
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12820 12782 12848 13874
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12102 12664 12582
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11694 12664 12038
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12438 8936 12494 8945
rect 12360 8894 12438 8922
rect 12254 8392 12310 8401
rect 12254 8327 12310 8336
rect 12256 7744 12308 7750
rect 12256 7686 12308 7692
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12268 4078 12296 7686
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12360 3738 12388 8894
rect 12438 8871 12494 8880
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12544 8498 12572 8842
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7206 12480 8230
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 6934 12480 7142
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12452 5846 12480 6870
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 12544 3942 12572 3975
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12360 2990 12388 3674
rect 12348 2984 12400 2990
rect 12070 2952 12126 2961
rect 12348 2926 12400 2932
rect 12070 2887 12126 2896
rect 12084 2582 12112 2887
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 2650 12572 2790
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11058 54 11192 82
rect 11978 82 12034 480
rect 12084 82 12112 2314
rect 11978 54 12112 82
rect 12636 82 12664 11630
rect 12820 11014 12848 11698
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12728 8634 12756 10134
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12728 7342 12756 7686
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12728 4758 12756 5102
rect 12716 4752 12768 4758
rect 12716 4694 12768 4700
rect 12820 4154 12848 10950
rect 12912 8022 12940 15914
rect 13004 10674 13032 17138
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13096 14822 13124 15506
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13096 12288 13124 14758
rect 13188 14482 13216 14826
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13188 13394 13216 14010
rect 13372 13870 13400 14418
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13188 12646 13216 13330
rect 13280 13258 13308 13670
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12646 13308 13194
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13096 12260 13216 12288
rect 13084 12164 13136 12170
rect 13084 12106 13136 12112
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13096 9722 13124 12106
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13096 9518 13124 9658
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9178 13124 9318
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12992 8016 13044 8022
rect 13188 7970 13216 12260
rect 13280 11762 13308 12582
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 12992 7958 13044 7964
rect 12912 7002 12940 7958
rect 13004 7410 13032 7958
rect 13096 7942 13216 7970
rect 13096 7818 13124 7942
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13004 6458 13032 7346
rect 13188 6934 13216 7822
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13004 6186 13032 6394
rect 13280 6322 13308 8298
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 13280 5234 13308 6258
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13266 5128 13322 5137
rect 13266 5063 13322 5072
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12728 4126 12848 4154
rect 12728 3466 12756 4126
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12820 2961 12848 3538
rect 12912 3505 12940 4762
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 13096 4486 13124 4626
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13280 3738 13308 5063
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13372 3602 13400 13806
rect 13556 13308 13584 15846
rect 13648 15706 13676 16594
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13556 13280 13676 13308
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13556 12306 13584 12718
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13464 11354 13492 11834
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13464 10470 13492 11290
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13464 10198 13492 10406
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13464 8634 13492 8978
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13556 7546 13584 11766
rect 13648 11150 13676 13280
rect 13740 12238 13768 16730
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13648 9586 13676 10678
rect 13740 9722 13768 10950
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 9178 13676 9522
rect 13740 9450 13768 9658
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13832 8498 13860 17138
rect 13924 16998 13952 17682
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16658 13952 16934
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 13190 13952 14758
rect 14004 13728 14056 13734
rect 14004 13670 14056 13676
rect 14016 13530 14044 13670
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 14016 12918 14044 13466
rect 14108 13394 14136 17614
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14200 16522 14228 17070
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14016 12714 14044 12854
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 14016 12374 14044 12650
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11286 13952 12038
rect 14016 11898 14044 12310
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13912 11280 13964 11286
rect 13912 11222 13964 11228
rect 13924 10198 13952 11222
rect 14016 10810 14044 11494
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14016 10198 14044 10746
rect 14108 10470 14136 10950
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 13924 9654 13952 10134
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13924 9042 13952 9590
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13464 5370 13492 5782
rect 13728 5704 13780 5710
rect 13634 5672 13690 5681
rect 13690 5652 13728 5658
rect 13690 5646 13780 5652
rect 13690 5630 13768 5646
rect 13634 5607 13690 5616
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 14096 5092 14148 5098
rect 14096 5034 14148 5040
rect 14108 4826 14136 5034
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3738 13860 3878
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 13372 3194 13400 3538
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12806 2952 12862 2961
rect 12806 2887 12808 2896
rect 12860 2887 12862 2896
rect 12808 2858 12860 2864
rect 12820 2827 12848 2858
rect 13740 2854 13768 3402
rect 14200 3194 14228 16458
rect 14292 15638 14320 16594
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14280 15632 14332 15638
rect 14280 15574 14332 15580
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14292 13376 14320 15370
rect 14384 14278 14412 15370
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 13530 14412 14214
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14292 13348 14412 13376
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 11234 14320 13194
rect 14384 12186 14412 13348
rect 14476 13326 14504 13806
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12374 14504 12582
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14384 12158 14504 12186
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14384 11354 14412 11562
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14292 11206 14412 11234
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14292 9586 14320 9930
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 14292 8090 14320 8298
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14292 7886 14320 8026
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14384 4154 14412 11206
rect 14476 8974 14504 12158
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14568 7426 14596 16526
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15212 15434 15240 16050
rect 15200 15428 15252 15434
rect 15200 15370 15252 15376
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14660 14113 14688 15098
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14646 14104 14702 14113
rect 14646 14039 14702 14048
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14660 10742 14688 13466
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14660 9722 14688 9998
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14660 9382 14688 9658
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14476 7398 14596 7426
rect 14476 6866 14504 7398
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14476 6458 14504 6802
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14568 6322 14596 6938
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14568 5914 14596 6258
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14660 5302 14688 8434
rect 14752 7546 14780 14962
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14844 14550 14872 14826
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14844 13814 14872 14486
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14844 13786 14964 13814
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14844 12986 14872 13330
rect 14936 13258 14964 13786
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15304 12889 15332 17478
rect 15580 17202 15608 17682
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15660 17128 15712 17134
rect 15660 17070 15712 17076
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15396 16250 15424 16594
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 15488 15910 15516 16594
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15396 14482 15424 15506
rect 15488 14482 15516 15846
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 14958 15608 15302
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15476 14476 15528 14482
rect 15476 14418 15528 14424
rect 15488 13802 15516 14418
rect 15476 13796 15528 13802
rect 15476 13738 15528 13744
rect 15290 12880 15346 12889
rect 15290 12815 15346 12824
rect 15488 12782 15516 13738
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15476 12776 15528 12782
rect 15476 12718 15528 12724
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14752 7342 14780 7482
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14292 4126 14412 4154
rect 14464 4208 14516 4214
rect 14464 4154 14516 4156
rect 14844 4154 14872 12718
rect 15384 12708 15436 12714
rect 15304 12668 15384 12696
rect 15304 12102 15332 12668
rect 15384 12650 15436 12656
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15304 11762 15332 12038
rect 15396 11898 15424 12310
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15488 11354 15516 12174
rect 15580 11830 15608 14894
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 10266 15148 10474
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14464 4150 14872 4154
rect 14476 4126 14872 4150
rect 15304 4154 15332 10746
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15396 9722 15424 10134
rect 15488 10062 15516 11290
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15580 10674 15608 11086
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15476 10056 15528 10062
rect 15476 9998 15528 10004
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15396 8634 15424 9658
rect 15672 9024 15700 17070
rect 15844 17060 15896 17066
rect 15896 17020 15976 17048
rect 15844 17002 15896 17008
rect 15844 16040 15896 16046
rect 15750 16008 15806 16017
rect 15844 15982 15896 15988
rect 15750 15943 15806 15952
rect 15764 15706 15792 15943
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15752 14952 15804 14958
rect 15856 14940 15884 15982
rect 15804 14912 15884 14940
rect 15752 14894 15804 14900
rect 15764 14822 15792 14894
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15948 14346 15976 17020
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 12714 15792 13806
rect 15856 13258 15884 13942
rect 15948 13734 15976 14282
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15844 13252 15896 13258
rect 15844 13194 15896 13200
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11694 15792 12038
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15488 8996 15700 9024
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15384 8288 15436 8294
rect 15384 8230 15436 8236
rect 15396 6458 15424 8230
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15396 5166 15424 6394
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15396 4826 15424 5102
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15304 4126 15424 4154
rect 14292 3602 14320 4126
rect 14476 4078 14504 4126
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14292 3126 14320 3538
rect 14370 3496 14426 3505
rect 14370 3431 14426 3440
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12990 82 13046 480
rect 12636 54 13046 82
rect 13740 82 13768 2790
rect 14384 2582 14412 3431
rect 14372 2576 14424 2582
rect 14372 2518 14424 2524
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 14200 1873 14228 2382
rect 14186 1864 14242 1873
rect 14186 1799 14242 1808
rect 13910 82 13966 480
rect 13740 54 13966 82
rect 14476 82 14504 4014
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3398 14872 3878
rect 15396 3466 15424 4126
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 2972 14872 3334
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15488 3058 15516 8996
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15672 7954 15700 8230
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15580 6730 15608 7686
rect 15672 6934 15700 7686
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15672 6372 15700 6870
rect 15580 6344 15700 6372
rect 15580 5914 15608 6344
rect 15764 6322 15792 10678
rect 15856 10033 15884 11018
rect 15948 10810 15976 13670
rect 16040 11880 16068 16934
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 16856 16652 16908 16658
rect 16856 16594 16908 16600
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16684 16250 16712 16458
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16132 14550 16160 16186
rect 16868 15910 16896 16594
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 13530 16252 14214
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16408 13462 16436 14350
rect 16500 13870 16528 14554
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16396 13456 16448 13462
rect 16396 13398 16448 13404
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16040 11852 16160 11880
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16040 11150 16068 11698
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 16040 10742 16068 11086
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 15842 10024 15898 10033
rect 15842 9959 15898 9968
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9489 15976 9522
rect 15934 9480 15990 9489
rect 15934 9415 15990 9424
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8362 15884 8774
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15948 8362 15976 8570
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15856 7818 15884 8298
rect 16132 8090 16160 11852
rect 16224 11626 16252 13126
rect 16394 13016 16450 13025
rect 16394 12951 16450 12960
rect 16408 12918 16436 12951
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16408 12374 16436 12854
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11642 16344 12038
rect 16408 11762 16436 12310
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16212 11620 16264 11626
rect 16316 11614 16436 11642
rect 16212 11562 16264 11568
rect 16408 10742 16436 11614
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16224 9024 16252 9930
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9450 16344 9862
rect 16408 9586 16436 10678
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16304 9444 16356 9450
rect 16304 9386 16356 9392
rect 16304 9036 16356 9042
rect 16224 8996 16304 9024
rect 16304 8978 16356 8984
rect 16316 8838 16344 8978
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 8412 16344 8774
rect 16408 8566 16436 9522
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16316 8384 16436 8412
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 16132 7324 16160 8026
rect 16316 7857 16344 8026
rect 16408 7886 16436 8384
rect 16396 7880 16448 7886
rect 16302 7848 16358 7857
rect 16396 7822 16448 7828
rect 16302 7783 16358 7792
rect 16408 7546 16436 7822
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16212 7336 16264 7342
rect 16132 7296 16212 7324
rect 16212 7278 16264 7284
rect 16224 6934 16252 7278
rect 16212 6928 16264 6934
rect 16212 6870 16264 6876
rect 15844 6860 15896 6866
rect 15844 6802 15896 6808
rect 15752 6316 15804 6322
rect 15672 6276 15752 6304
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15580 5370 15608 5850
rect 15672 5710 15700 6276
rect 15752 6258 15804 6264
rect 15750 6216 15806 6225
rect 15750 6151 15806 6160
rect 15764 5914 15792 6151
rect 15856 6118 15884 6802
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 6390 16344 6598
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16316 6254 16344 6326
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15672 4808 15700 5646
rect 15672 4780 15792 4808
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15580 3942 15608 4626
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15580 3058 15608 3878
rect 15672 3670 15700 4626
rect 15764 4622 15792 4780
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15764 4282 15792 4422
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15856 4154 15884 6054
rect 16120 5772 16172 5778
rect 16120 5714 16172 5720
rect 16132 4622 16160 5714
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 15764 4126 15884 4154
rect 15764 3738 15792 4126
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15660 3664 15712 3670
rect 15660 3606 15712 3612
rect 16132 3602 16160 4558
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15016 2984 15068 2990
rect 14844 2944 15016 2972
rect 15016 2926 15068 2932
rect 15028 2650 15056 2926
rect 15948 2854 15976 3402
rect 16316 2922 16344 4422
rect 16500 4282 16528 13126
rect 16592 12238 16620 13670
rect 16684 13394 16712 14758
rect 16868 14006 16896 15846
rect 16856 14000 16908 14006
rect 16856 13942 16908 13948
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16592 9042 16620 9590
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16592 7954 16620 8978
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 16592 7546 16620 7890
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16592 7410 16620 7482
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16592 6866 16620 7346
rect 16684 7274 16712 12854
rect 16776 9722 16804 13806
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 12918 16896 13670
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16764 9716 16816 9722
rect 16764 9658 16816 9664
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6866 16712 7210
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16592 6458 16620 6802
rect 16762 6760 16818 6769
rect 16762 6695 16818 6704
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16776 6322 16804 6695
rect 16764 6316 16816 6322
rect 16764 6258 16816 6264
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5914 16620 6190
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16868 5778 16896 12650
rect 16960 9178 16988 13942
rect 17052 13734 17080 16390
rect 17592 16176 17644 16182
rect 17592 16118 17644 16124
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17236 14822 17264 15506
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17052 13394 17080 13466
rect 17040 13388 17092 13394
rect 17236 13376 17264 14758
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17328 13938 17356 14214
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 13530 17356 13874
rect 17512 13814 17540 14418
rect 17420 13786 17540 13814
rect 17420 13734 17448 13786
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17316 13388 17368 13394
rect 17092 13348 17172 13376
rect 17236 13348 17316 13376
rect 17040 13330 17092 13336
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17052 12646 17080 13194
rect 17144 12986 17172 13348
rect 17316 13330 17368 13336
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 9172 17000 9178
rect 16948 9114 17000 9120
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16960 8634 16988 8978
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16960 7954 16988 8570
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16960 7478 16988 7890
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 6730 16988 7278
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16868 5098 16896 5714
rect 16856 5092 16908 5098
rect 16856 5034 16908 5040
rect 17052 4758 17080 12582
rect 17144 9042 17172 12922
rect 17328 12714 17356 13330
rect 17420 13161 17448 13670
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17406 13152 17462 13161
rect 17406 13087 17462 13096
rect 17420 12753 17448 13087
rect 17406 12744 17462 12753
rect 17316 12708 17368 12714
rect 17406 12679 17462 12688
rect 17316 12650 17368 12656
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17236 11558 17264 12174
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17236 11354 17264 11494
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17420 9518 17448 11766
rect 17512 11286 17540 13466
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17512 10810 17540 11222
rect 17604 11218 17632 16118
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17788 13870 17816 15438
rect 17868 14816 17920 14822
rect 17868 14758 17920 14764
rect 17776 13864 17828 13870
rect 17696 13812 17776 13814
rect 17696 13806 17828 13812
rect 17696 13786 17816 13806
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17696 10962 17724 13786
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17604 10934 17724 10962
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17512 10198 17540 10746
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9586 17540 10134
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17132 9036 17184 9042
rect 17132 8978 17184 8984
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17236 8634 17264 8978
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17144 5914 17172 8502
rect 17236 8090 17264 8570
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 17236 6866 17264 8026
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17328 7342 17356 7890
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 5914 17264 6802
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17224 5908 17276 5914
rect 17224 5850 17276 5856
rect 17328 5846 17356 6870
rect 17604 6254 17632 10934
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17696 10130 17724 10746
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17696 9654 17724 10066
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17788 8430 17816 13262
rect 17880 12442 17908 14758
rect 18064 14618 18092 15982
rect 18420 15972 18472 15978
rect 18420 15914 18472 15920
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17972 12714 18000 14214
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 17972 11898 18000 12310
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17972 11626 18000 11834
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10130 17908 11154
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17880 7954 17908 9114
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17788 7274 17816 7822
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 6866 17816 7210
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17788 6458 17816 6802
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17972 6254 18000 10950
rect 18064 7342 18092 13398
rect 18156 11150 18184 15846
rect 18236 15632 18288 15638
rect 18236 15574 18288 15580
rect 18248 14958 18276 15574
rect 18432 15570 18460 15914
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18248 14278 18276 14894
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14550 18368 14826
rect 18432 14822 18460 15506
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 18248 12918 18276 14214
rect 18236 12912 18288 12918
rect 18236 12854 18288 12860
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18156 10810 18184 11086
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18234 8936 18290 8945
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 5370 17448 5646
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17420 4622 17448 5306
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 16488 4276 16540 4282
rect 16488 4218 16540 4224
rect 16592 4078 16620 4490
rect 17132 4276 17184 4282
rect 17132 4218 17184 4224
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16672 3936 16724 3942
rect 16672 3878 16724 3884
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15198 2680 15254 2689
rect 15016 2644 15068 2650
rect 15198 2615 15254 2624
rect 15016 2586 15068 2592
rect 15212 2582 15240 2615
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 14752 1193 14780 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14738 1184 14794 1193
rect 14738 1119 14794 1128
rect 14922 82 14978 480
rect 15764 134 15792 2246
rect 14476 54 14978 82
rect 15752 128 15804 134
rect 15752 70 15804 76
rect 15842 82 15898 480
rect 15948 82 15976 2790
rect 16316 2378 16344 2858
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 11058 0 11114 54
rect 11978 0 12034 54
rect 12990 0 13046 54
rect 13910 0 13966 54
rect 14922 0 14978 54
rect 15842 54 15976 82
rect 16592 82 16620 2994
rect 16684 2650 16712 3878
rect 16868 2922 16896 4014
rect 17144 3602 17172 4218
rect 17328 4049 17356 4558
rect 17420 4282 17448 4558
rect 17408 4276 17460 4282
rect 17408 4218 17460 4224
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17052 3126 17080 3538
rect 17408 3460 17460 3466
rect 17408 3402 17460 3408
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 16868 2378 16896 2858
rect 17144 2446 17172 2858
rect 17420 2854 17448 3402
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 16856 2372 16908 2378
rect 16856 2314 16908 2320
rect 17420 1465 17448 2790
rect 17406 1456 17462 1465
rect 17406 1391 17462 1400
rect 16854 82 16910 480
rect 16592 54 16910 82
rect 17512 82 17540 5034
rect 17696 4826 17724 5850
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17788 4282 17816 4966
rect 17972 4826 18000 5782
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17972 3602 18000 4762
rect 18156 3670 18184 8910
rect 18234 8871 18290 8880
rect 18248 8634 18276 8871
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18340 7002 18368 14486
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18432 6458 18460 14758
rect 18616 14657 18644 16390
rect 20442 16144 20498 16153
rect 20442 16079 20498 16088
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18602 14648 18658 14657
rect 18602 14583 18658 14592
rect 18510 14512 18566 14521
rect 18510 14447 18566 14456
rect 18524 13530 18552 14447
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18616 12986 18644 14214
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18524 12753 18552 12786
rect 18510 12744 18566 12753
rect 18510 12679 18566 12688
rect 18616 12646 18644 12922
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18708 12306 18736 12650
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 18800 10130 18828 15302
rect 18972 15088 19024 15094
rect 18972 15030 19024 15036
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18892 14074 18920 14418
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18892 13462 18920 14010
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 18892 12442 18920 13398
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18892 11014 18920 11630
rect 18984 11218 19012 15030
rect 19248 13252 19300 13258
rect 19248 13194 19300 13200
rect 19260 12918 19288 13194
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 11898 19196 12582
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 19352 11762 19380 15438
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19444 13870 19472 14214
rect 20364 14006 20392 14894
rect 20456 14385 20484 16079
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20442 14376 20498 14385
rect 20442 14311 20498 14320
rect 20536 14340 20588 14346
rect 20352 14000 20404 14006
rect 20350 13968 20352 13977
rect 20404 13968 20406 13977
rect 20350 13903 20406 13912
rect 20364 13877 20392 13903
rect 20456 13870 20484 14311
rect 20536 14282 20588 14288
rect 19432 13864 19484 13870
rect 20444 13864 20496 13870
rect 19484 13812 19564 13814
rect 19432 13806 19564 13812
rect 20444 13806 20496 13812
rect 19444 13786 19564 13806
rect 19432 13728 19484 13734
rect 19432 13670 19484 13676
rect 19444 11898 19472 13670
rect 19536 12646 19564 13786
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19996 13326 20024 13670
rect 20076 13456 20128 13462
rect 20076 13398 20128 13404
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 12986 20024 13262
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 20088 12306 20116 13398
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19904 11830 19932 12242
rect 20180 12186 20208 12922
rect 20442 12880 20498 12889
rect 20442 12815 20498 12824
rect 20456 12714 20484 12815
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20088 12158 20208 12186
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 18972 11212 19024 11218
rect 19024 11172 19104 11200
rect 18972 11154 19024 11160
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18892 10198 18920 10950
rect 19076 10538 19104 11172
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10713 19380 10950
rect 19536 10810 19564 11562
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19338 10704 19394 10713
rect 19338 10639 19340 10648
rect 19392 10639 19394 10648
rect 19340 10610 19392 10616
rect 19352 10579 19380 10610
rect 19536 10538 19564 10746
rect 19064 10532 19116 10538
rect 19064 10474 19116 10480
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18880 10192 18932 10198
rect 18880 10134 18932 10140
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18524 9042 18552 9454
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18524 8566 18552 8978
rect 18512 8560 18564 8566
rect 18512 8502 18564 8508
rect 18616 7410 18644 10066
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 8022 18736 9318
rect 18800 9178 18828 10066
rect 18880 10056 18932 10062
rect 18880 9998 18932 10004
rect 18892 9518 18920 9998
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18892 9042 18920 9454
rect 18984 9382 19012 10406
rect 19076 10266 19104 10474
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19076 9586 19104 10202
rect 19156 10056 19208 10062
rect 19156 9998 19208 10004
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18800 7954 18828 8366
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 8022 18920 8230
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18616 6934 18644 7346
rect 18800 7342 18828 7890
rect 18892 7478 18920 7958
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18616 6390 18644 6870
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18696 6180 18748 6186
rect 18696 6122 18748 6128
rect 18328 6112 18380 6118
rect 18328 6054 18380 6060
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18248 5370 18276 5714
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18248 4690 18276 5306
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18248 4282 18276 4626
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18340 4146 18368 6054
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17696 2922 17724 3538
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 2961 17816 2994
rect 17774 2952 17830 2961
rect 17684 2916 17736 2922
rect 17774 2887 17830 2896
rect 17684 2858 17736 2864
rect 17696 2650 17724 2858
rect 17788 2854 17816 2887
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 18432 2514 18460 3402
rect 18708 2836 18736 6122
rect 18800 5370 18828 6938
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18788 5364 18840 5370
rect 18788 5306 18840 5312
rect 18800 3602 18828 5306
rect 18892 3942 18920 6258
rect 19076 6254 19104 7278
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19076 5914 19104 6190
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 19076 5166 19104 5850
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18984 4690 19012 4762
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 2990 18828 3334
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 18892 2922 18920 3878
rect 18984 2990 19012 4626
rect 19076 4146 19104 5102
rect 19168 4486 19196 9998
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19352 9042 19380 9386
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 19260 7886 19288 8366
rect 19340 8084 19392 8090
rect 19340 8026 19392 8032
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19260 7342 19288 7822
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19260 6254 19288 7278
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19352 5778 19380 8026
rect 19536 7954 19564 9046
rect 19996 8430 20024 9454
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19996 8090 20024 8366
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19444 7002 19472 7210
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19996 6458 20024 7278
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19996 6254 20024 6394
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20088 6118 20116 12158
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20180 11626 20208 11834
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20272 11354 20300 11698
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 4826 19380 5714
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 19156 4480 19208 4486
rect 19156 4422 19208 4428
rect 19064 4140 19116 4146
rect 19116 4100 19288 4128
rect 19064 4082 19116 4088
rect 19260 3738 19288 4100
rect 19444 4078 19472 5034
rect 19996 5030 20024 5102
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19996 4078 20024 4966
rect 20180 4282 20208 10950
rect 20272 7562 20300 10950
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 9382 20392 10066
rect 20456 9926 20484 11154
rect 20444 9920 20496 9926
rect 20444 9862 20496 9868
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 9081 20392 9318
rect 20350 9072 20406 9081
rect 20350 9007 20406 9016
rect 20364 8906 20392 9007
rect 20352 8900 20404 8906
rect 20352 8842 20404 8848
rect 20272 7534 20392 7562
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20272 5914 20300 6598
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19984 4072 20036 4078
rect 19984 4014 20036 4020
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19444 3398 19472 4014
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20364 3505 20392 7534
rect 20456 4154 20484 9862
rect 20548 9058 20576 14282
rect 20640 13802 20668 14418
rect 20628 13796 20680 13802
rect 20628 13738 20680 13744
rect 20640 12850 20668 13738
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 11830 20668 12786
rect 20732 12442 20760 13330
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20732 11286 20760 12378
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20732 10810 20760 11222
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20548 9030 20668 9058
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20548 8498 20576 8910
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20640 5778 20668 9030
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 6662 20760 7686
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20628 5772 20680 5778
rect 20628 5714 20680 5720
rect 20640 4826 20668 5714
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 20456 4126 20668 4154
rect 20350 3496 20406 3505
rect 20350 3431 20406 3440
rect 20536 3460 20588 3466
rect 20536 3402 20588 3408
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20456 3058 20484 3334
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18788 2848 18840 2854
rect 18708 2808 18788 2836
rect 18708 2650 18736 2808
rect 18788 2790 18840 2796
rect 18984 2650 19012 2926
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17774 82 17830 480
rect 17512 54 17830 82
rect 18708 82 18736 2586
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19352 2106 19380 2246
rect 19340 2100 19392 2106
rect 19340 2042 19392 2048
rect 18786 82 18842 480
rect 18708 54 18842 82
rect 15842 0 15898 54
rect 16854 0 16910 54
rect 17774 0 17830 54
rect 18786 0 18842 54
rect 19706 128 19762 480
rect 19706 76 19708 128
rect 19760 76 19762 128
rect 19706 0 19762 76
rect 20548 82 20576 3402
rect 20640 2650 20668 4126
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20732 2922 20760 3878
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20640 2310 20668 2450
rect 20824 2310 20852 16526
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20904 14272 20956 14278
rect 20904 14214 20956 14220
rect 20916 13814 20944 14214
rect 20916 13786 21036 13814
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20916 11150 20944 12038
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9654 20944 9998
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20916 9110 20944 9590
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20916 7206 20944 7890
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 20640 785 20668 2246
rect 20916 2009 20944 7142
rect 21008 2990 21036 13786
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 11898 21128 12242
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21100 10810 21128 11834
rect 21088 10804 21140 10810
rect 21088 10746 21140 10752
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21100 10198 21128 10474
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 21100 9722 21128 10134
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21100 9178 21128 9658
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 21100 7546 21128 9114
rect 21192 8566 21220 15302
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21456 14884 21508 14890
rect 21456 14826 21508 14832
rect 21468 13274 21496 14826
rect 21284 13246 21496 13274
rect 21180 8560 21232 8566
rect 21180 8502 21232 8508
rect 21284 8498 21312 13246
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 11898 21404 13126
rect 21456 12096 21508 12102
rect 21456 12038 21508 12044
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21376 11558 21404 11834
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21468 9722 21496 12038
rect 21560 11830 21588 14894
rect 21548 11824 21600 11830
rect 21548 11766 21600 11772
rect 21560 11354 21588 11766
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21456 9716 21508 9722
rect 21456 9658 21508 9664
rect 21468 9450 21496 9658
rect 21652 9654 21680 15438
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21652 9178 21680 9590
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21548 8560 21600 8566
rect 21548 8502 21600 8508
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21100 7274 21128 7482
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21100 5370 21128 6938
rect 21192 6934 21220 8230
rect 21284 8090 21312 8434
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 21364 7744 21416 7750
rect 21284 7704 21364 7732
rect 21284 7342 21312 7704
rect 21364 7686 21416 7692
rect 21468 7410 21496 7890
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21180 6928 21232 6934
rect 21180 6870 21232 6876
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21192 5778 21220 6122
rect 21284 5846 21312 7278
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21376 6934 21404 7142
rect 21364 6928 21416 6934
rect 21364 6870 21416 6876
rect 21560 6798 21588 8502
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21180 5772 21232 5778
rect 21180 5714 21232 5720
rect 21088 5364 21140 5370
rect 21088 5306 21140 5312
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 21100 4758 21128 5306
rect 21284 4826 21312 5306
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 21100 3738 21128 4558
rect 21284 4154 21312 4762
rect 21192 4126 21312 4154
rect 21192 3942 21220 4126
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 21376 3194 21404 6054
rect 21744 3670 21772 15846
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 12646 21864 13194
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21928 11286 21956 11698
rect 22020 11336 22048 16118
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22100 15564 22152 15570
rect 22100 15506 22152 15512
rect 22112 14822 22140 15506
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22112 13433 22140 14758
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22296 13734 22324 14418
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22098 13424 22154 13433
rect 22098 13359 22154 13368
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22020 11308 22140 11336
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21928 10674 21956 11222
rect 22008 11212 22060 11218
rect 22008 11154 22060 11160
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21836 10266 21864 10474
rect 21928 10266 21956 10610
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 22020 9926 22048 11154
rect 22008 9920 22060 9926
rect 22008 9862 22060 9868
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 6934 21864 8434
rect 21824 6928 21876 6934
rect 21876 6888 21956 6916
rect 21824 6870 21876 6876
rect 21824 5568 21876 5574
rect 21824 5510 21876 5516
rect 21836 5234 21864 5510
rect 21824 5228 21876 5234
rect 21824 5170 21876 5176
rect 21928 4758 21956 6888
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 22020 4622 22048 9862
rect 22112 8106 22140 11308
rect 22204 10577 22232 13262
rect 22190 10568 22246 10577
rect 22296 10538 22324 13670
rect 22374 13424 22430 13433
rect 22374 13359 22430 13368
rect 22388 13161 22416 13359
rect 22374 13152 22430 13161
rect 22374 13087 22430 13096
rect 22480 11234 22508 15846
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22388 11206 22508 11234
rect 22190 10503 22246 10512
rect 22284 10532 22336 10538
rect 22284 10474 22336 10480
rect 22296 9654 22324 10474
rect 22284 9648 22336 9654
rect 22284 9590 22336 9596
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22296 8634 22324 9046
rect 22284 8628 22336 8634
rect 22284 8570 22336 8576
rect 22112 8078 22324 8106
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 22112 7002 22140 7822
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22100 6180 22152 6186
rect 22100 6122 22152 6128
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 21822 4040 21878 4049
rect 21822 3975 21878 3984
rect 21836 3670 21864 3975
rect 21732 3664 21784 3670
rect 21732 3606 21784 3612
rect 21824 3664 21876 3670
rect 21824 3606 21876 3612
rect 21744 3194 21772 3606
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 20996 2984 21048 2990
rect 20996 2926 21048 2932
rect 21376 2582 21404 3130
rect 21836 3058 21864 3606
rect 22020 3534 22048 4558
rect 22112 3670 22140 6122
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22204 4826 22232 5714
rect 22296 5681 22324 8078
rect 22388 7546 22416 11206
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22480 10810 22508 11086
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22572 9042 22600 13670
rect 22652 13388 22704 13394
rect 22652 13330 22704 13336
rect 22664 12646 22692 13330
rect 22756 13326 22784 16050
rect 22744 13320 22796 13326
rect 22744 13262 22796 13268
rect 22836 13184 22888 13190
rect 22756 13144 22836 13172
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22282 5672 22338 5681
rect 22282 5607 22338 5616
rect 22192 4820 22244 4826
rect 22192 4762 22244 4768
rect 22480 4554 22508 8774
rect 22560 8628 22612 8634
rect 22560 8570 22612 8576
rect 22572 8022 22600 8570
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22572 7478 22600 7958
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22572 5914 22600 7414
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22572 5370 22600 5850
rect 22664 5778 22692 12582
rect 22756 9058 22784 13144
rect 22836 13126 22888 13132
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22848 10441 22876 12922
rect 22834 10432 22890 10441
rect 22834 10367 22890 10376
rect 22940 10033 22968 16934
rect 23112 15972 23164 15978
rect 23112 15914 23164 15920
rect 23020 13728 23072 13734
rect 23020 13670 23072 13676
rect 23032 12986 23060 13670
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 23124 11540 23152 15914
rect 23296 15564 23348 15570
rect 23296 15506 23348 15512
rect 23308 14822 23336 15506
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23032 11512 23152 11540
rect 23032 10198 23060 11512
rect 23308 11268 23336 14758
rect 23492 12753 23520 23598
rect 23662 20904 23718 20913
rect 23662 20839 23718 20848
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 16182 23612 16594
rect 23572 16176 23624 16182
rect 23572 16118 23624 16124
rect 23676 12918 23704 20839
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23768 13734 23796 14418
rect 23952 14006 23980 24783
rect 24122 23760 24178 23769
rect 24122 23695 24178 23704
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 24044 14618 24072 21422
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23768 13025 23796 13670
rect 24136 13530 24164 23695
rect 24228 15162 24256 25735
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24780 23866 24808 26823
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24766 22672 24822 22681
rect 24766 22607 24822 22616
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24780 21690 24808 22607
rect 25410 21720 25466 21729
rect 24768 21684 24820 21690
rect 25410 21655 25466 21664
rect 24768 21626 24820 21632
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24766 18592 24822 18601
rect 24289 18524 24585 18544
rect 24766 18527 24822 18536
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24780 17882 24808 18527
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24584 16992 24636 16998
rect 24688 16980 24716 17682
rect 24766 17504 24822 17513
rect 24766 17439 24822 17448
rect 24636 16952 24716 16980
rect 24584 16934 24636 16940
rect 24596 16794 24624 16934
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24780 16658 24808 17439
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24780 16250 24808 16594
rect 25226 16552 25282 16561
rect 25226 16487 25282 16496
rect 25240 16250 25268 16487
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25240 16046 25268 16186
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24674 15464 24730 15473
rect 24674 15399 24730 15408
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24688 14482 24716 15399
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14418
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 24214 13424 24270 13433
rect 23940 13388 23992 13394
rect 24214 13359 24216 13368
rect 23940 13330 23992 13336
rect 24268 13359 24270 13368
rect 24216 13330 24268 13336
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23754 13016 23810 13025
rect 23754 12951 23810 12960
rect 23664 12912 23716 12918
rect 23664 12854 23716 12860
rect 23478 12744 23534 12753
rect 23478 12679 23534 12688
rect 23572 12300 23624 12306
rect 23572 12242 23624 12248
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23216 11240 23336 11268
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23124 10810 23152 11154
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23020 10192 23072 10198
rect 23020 10134 23072 10140
rect 22926 10024 22982 10033
rect 22926 9959 22982 9968
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 23032 9874 23060 10134
rect 23124 9994 23152 10746
rect 23216 10169 23244 11240
rect 23296 11144 23348 11150
rect 23296 11086 23348 11092
rect 23202 10160 23258 10169
rect 23202 10095 23258 10104
rect 23204 10056 23256 10062
rect 23204 9998 23256 10004
rect 23112 9988 23164 9994
rect 23112 9930 23164 9936
rect 22940 9178 22968 9862
rect 23032 9846 23152 9874
rect 23018 9752 23074 9761
rect 23124 9722 23152 9846
rect 23018 9687 23074 9696
rect 23112 9716 23164 9722
rect 22928 9172 22980 9178
rect 22928 9114 22980 9120
rect 22756 9030 22876 9058
rect 22744 8968 22796 8974
rect 22744 8910 22796 8916
rect 22756 8634 22784 8910
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22848 7478 22876 9030
rect 23032 8566 23060 9687
rect 23112 9658 23164 9664
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23020 8356 23072 8362
rect 23020 8298 23072 8304
rect 23032 8090 23060 8298
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22756 6458 22784 6802
rect 22744 6452 22796 6458
rect 22796 6412 22876 6440
rect 22744 6394 22796 6400
rect 22744 6180 22796 6186
rect 22744 6122 22796 6128
rect 22652 5772 22704 5778
rect 22652 5714 22704 5720
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22560 5364 22612 5370
rect 22560 5306 22612 5312
rect 22664 4842 22692 5578
rect 22756 5370 22784 6122
rect 22848 5914 22876 6412
rect 22836 5908 22888 5914
rect 22836 5850 22888 5856
rect 22744 5364 22796 5370
rect 22744 5306 22796 5312
rect 22664 4814 22784 4842
rect 22560 4752 22612 4758
rect 22560 4694 22612 4700
rect 22468 4548 22520 4554
rect 22468 4490 22520 4496
rect 22572 4282 22600 4694
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 22480 4154 22508 4218
rect 22480 4126 22600 4154
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22572 3058 22600 4126
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21364 2576 21416 2582
rect 21364 2518 21416 2524
rect 20902 2000 20958 2009
rect 20902 1935 20958 1944
rect 20626 776 20682 785
rect 20626 711 20682 720
rect 20718 82 20774 480
rect 20548 54 20774 82
rect 20718 0 20774 54
rect 21638 82 21694 480
rect 21744 82 21772 2790
rect 22664 2650 22692 4490
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 21638 54 21772 82
rect 22650 82 22706 480
rect 22756 82 22784 4814
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 22848 4486 22876 4694
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22848 4214 22876 4422
rect 23124 4214 23152 9046
rect 23216 8498 23244 9998
rect 23308 9450 23336 11086
rect 23492 10810 23520 12174
rect 23584 11898 23612 12242
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23492 10470 23520 10746
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23386 10296 23442 10305
rect 23386 10231 23442 10240
rect 23400 9586 23428 10231
rect 23584 10180 23612 11834
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23664 10192 23716 10198
rect 23584 10152 23664 10180
rect 23584 9926 23612 10152
rect 23664 10134 23716 10140
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23584 9722 23612 9862
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 9444 23348 9450
rect 23296 9386 23348 9392
rect 23768 8634 23796 11630
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23204 8492 23256 8498
rect 23204 8434 23256 8440
rect 23216 8090 23244 8434
rect 23768 8362 23796 8570
rect 23756 8356 23808 8362
rect 23756 8298 23808 8304
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23400 5370 23428 6734
rect 23860 6322 23888 13126
rect 23952 12646 23980 13330
rect 24228 12986 24256 13330
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 23952 9110 23980 9930
rect 24044 9722 24072 11086
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 23940 9104 23992 9110
rect 23940 9046 23992 9052
rect 23952 8634 23980 9046
rect 24032 8968 24084 8974
rect 24032 8910 24084 8916
rect 23940 8628 23992 8634
rect 23940 8570 23992 8576
rect 24044 6882 24072 8910
rect 24136 7274 24164 11494
rect 24228 8616 24256 12582
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24320 10198 24348 10610
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24596 8974 24624 9522
rect 24688 9489 24716 9862
rect 24674 9480 24730 9489
rect 24674 9415 24730 9424
rect 24584 8968 24636 8974
rect 24584 8910 24636 8916
rect 24780 8906 24808 15302
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24872 10554 24900 14214
rect 24964 10810 24992 15846
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25226 12336 25282 12345
rect 25136 12300 25188 12306
rect 25226 12271 25282 12280
rect 25136 12242 25188 12248
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24952 10804 25004 10810
rect 24952 10746 25004 10752
rect 24872 10526 24992 10554
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24768 8900 24820 8906
rect 24768 8842 24820 8848
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24768 8628 24820 8634
rect 24228 8588 24348 8616
rect 24320 8537 24348 8588
rect 24768 8570 24820 8576
rect 24306 8528 24362 8537
rect 24216 8492 24268 8498
rect 24306 8463 24362 8472
rect 24216 8434 24268 8440
rect 24228 7410 24256 8434
rect 24780 8090 24808 8570
rect 24872 8401 24900 10406
rect 24964 10305 24992 10526
rect 24950 10296 25006 10305
rect 24950 10231 24952 10240
rect 25004 10231 25006 10240
rect 24952 10202 25004 10208
rect 24964 10171 24992 10202
rect 24858 8392 24914 8401
rect 24858 8327 24914 8336
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24964 7546 24992 7822
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 24124 7268 24176 7274
rect 24124 7210 24176 7216
rect 24136 7002 24164 7210
rect 25056 7002 25084 12038
rect 25148 11626 25176 12242
rect 25240 11694 25268 12271
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 25136 11620 25188 11626
rect 25136 11562 25188 11568
rect 25332 10248 25360 15438
rect 25424 11898 25452 21655
rect 26146 19544 26202 19553
rect 26146 19479 26202 19488
rect 25412 11892 25464 11898
rect 25412 11834 25464 11840
rect 25412 11212 25464 11218
rect 25412 11154 25464 11160
rect 25424 10674 25452 11154
rect 25502 10704 25558 10713
rect 25412 10668 25464 10674
rect 25502 10639 25558 10648
rect 25412 10610 25464 10616
rect 25148 10220 25360 10248
rect 24124 6996 24176 7002
rect 24124 6938 24176 6944
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 24676 6928 24728 6934
rect 24044 6854 24256 6882
rect 24676 6870 24728 6876
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 23860 5914 23888 6258
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23388 5364 23440 5370
rect 23388 5306 23440 5312
rect 24136 4826 24164 6258
rect 24228 5710 24256 6854
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6118 24716 6870
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24780 6322 24808 6734
rect 25056 6458 25084 6938
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 24216 5704 24268 5710
rect 24216 5646 24268 5652
rect 24228 5370 24256 5646
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24412 5098 24440 5238
rect 24400 5092 24452 5098
rect 24400 5034 24452 5040
rect 24688 4826 24716 6054
rect 24768 5636 24820 5642
rect 24768 5578 24820 5584
rect 24780 5234 24808 5578
rect 24768 5228 24820 5234
rect 24768 5170 24820 5176
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24676 4820 24728 4826
rect 24676 4762 24728 4768
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 23112 4208 23164 4214
rect 23112 4150 23164 4156
rect 24136 4146 24164 4762
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 24768 4004 24820 4010
rect 24768 3946 24820 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 22836 3664 22888 3670
rect 22836 3606 22888 3612
rect 23202 3632 23258 3641
rect 22848 2650 22876 3606
rect 23202 3567 23258 3576
rect 23216 3534 23244 3567
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23216 3194 23244 3470
rect 23768 3398 23796 3878
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23768 2990 23796 3334
rect 24136 3058 24164 3606
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3097 24716 3878
rect 24780 3670 24808 3946
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 24674 3088 24730 3097
rect 24124 3052 24176 3058
rect 24674 3023 24730 3032
rect 24124 2994 24176 3000
rect 23756 2984 23808 2990
rect 23756 2926 23808 2932
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 24676 2304 24728 2310
rect 24676 2246 24728 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23662 1184 23718 1193
rect 23662 1119 23718 1128
rect 22650 54 22784 82
rect 23570 82 23626 480
rect 23676 82 23704 1119
rect 24688 1057 24716 2246
rect 24674 1048 24730 1057
rect 24674 983 24730 992
rect 23570 54 23704 82
rect 24582 82 24638 480
rect 24964 82 24992 6326
rect 25044 6180 25096 6186
rect 25044 6122 25096 6128
rect 25056 4690 25084 6122
rect 25148 5030 25176 10220
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25332 9382 25360 10066
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25228 8900 25280 8906
rect 25228 8842 25280 8848
rect 25240 6254 25268 8842
rect 25332 8265 25360 9318
rect 25516 9178 25544 10639
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25504 9172 25556 9178
rect 25504 9114 25556 9120
rect 25780 9036 25832 9042
rect 25780 8978 25832 8984
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25424 8430 25452 8774
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 25792 8294 25820 8978
rect 25780 8288 25832 8294
rect 25318 8256 25374 8265
rect 25780 8230 25832 8236
rect 25318 8191 25374 8200
rect 25688 7200 25740 7206
rect 25688 7142 25740 7148
rect 25228 6248 25280 6254
rect 25228 6190 25280 6196
rect 25228 5840 25280 5846
rect 25228 5782 25280 5788
rect 25240 5370 25268 5782
rect 25228 5364 25280 5370
rect 25228 5306 25280 5312
rect 25136 5024 25188 5030
rect 25136 4966 25188 4972
rect 25044 4684 25096 4690
rect 25044 4626 25096 4632
rect 25056 4282 25084 4626
rect 25044 4276 25096 4282
rect 25044 4218 25096 4224
rect 24582 54 24992 82
rect 25502 82 25558 480
rect 25700 82 25728 7142
rect 25792 5137 25820 8230
rect 26068 5953 26096 10406
rect 26160 8634 26188 19479
rect 27618 13968 27674 13977
rect 27618 13903 27674 13912
rect 27632 13462 27660 13903
rect 27620 13456 27672 13462
rect 27620 13398 27672 13404
rect 27618 11792 27674 11801
rect 27618 11727 27674 11736
rect 27632 11626 27660 11727
rect 27620 11620 27672 11626
rect 27620 11562 27672 11568
rect 27712 10668 27764 10674
rect 27712 10610 27764 10616
rect 26148 8628 26200 8634
rect 26148 8570 26200 8576
rect 26146 6080 26202 6089
rect 26146 6015 26202 6024
rect 26054 5944 26110 5953
rect 26054 5879 26110 5888
rect 25778 5128 25834 5137
rect 25778 5063 25834 5072
rect 26160 4282 26188 6015
rect 26148 4276 26200 4282
rect 26148 4218 26200 4224
rect 26160 4078 26188 4218
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 26146 2952 26202 2961
rect 26146 2887 26202 2896
rect 26160 2650 26188 2887
rect 27528 2848 27580 2854
rect 27528 2790 27580 2796
rect 26148 2644 26200 2650
rect 26148 2586 26200 2592
rect 26608 2372 26660 2378
rect 26608 2314 26660 2320
rect 25502 54 25728 82
rect 26514 82 26570 480
rect 26620 82 26648 2314
rect 26514 54 26648 82
rect 27434 82 27490 480
rect 27540 82 27568 2790
rect 27724 2553 27752 10610
rect 27710 2544 27766 2553
rect 27710 2479 27766 2488
rect 27434 54 27568 82
rect 21638 0 21694 54
rect 22650 0 22706 54
rect 23570 0 23626 54
rect 24582 0 24638 54
rect 25502 0 25558 54
rect 26514 0 26570 54
rect 27434 0 27490 54
<< via2 >>
rect 1582 26832 1638 26888
rect 24766 26832 24822 26888
rect 1030 25744 1086 25800
rect 110 20032 166 20088
rect 110 6568 166 6624
rect 110 5616 166 5672
rect 938 17720 994 17776
rect 1490 23976 1546 24032
rect 1306 19760 1362 19816
rect 478 12144 534 12200
rect 386 10784 442 10840
rect 1398 18400 1454 18456
rect 1306 11736 1362 11792
rect 1122 11192 1178 11248
rect 294 8200 350 8256
rect 24214 25744 24270 25800
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 1674 24792 1730 24848
rect 23938 24792 23994 24848
rect 1582 22616 1638 22672
rect 1582 18536 1638 18592
rect 18 3440 74 3496
rect 1490 5072 1546 5128
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 1858 17584 1914 17640
rect 1950 16632 2006 16688
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 2134 14728 2190 14784
rect 1766 9560 1822 9616
rect 1950 6024 2006 6080
rect 2134 3848 2190 3904
rect 2134 3168 2190 3224
rect 2870 16360 2926 16416
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 2778 8200 2834 8256
rect 4342 17992 4398 18048
rect 3514 12280 3570 12336
rect 3974 15816 4030 15872
rect 4158 13368 4214 13424
rect 4342 13776 4398 13832
rect 4250 12416 4306 12472
rect 4618 14728 4674 14784
rect 1950 1536 2006 1592
rect 1858 992 1914 1048
rect 4618 9560 4674 9616
rect 4986 12300 5042 12336
rect 4986 12280 4988 12300
rect 4988 12280 5040 12300
rect 5040 12280 5042 12300
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 4986 10648 5042 10704
rect 5170 10104 5226 10160
rect 3790 3576 3846 3632
rect 4434 6024 4490 6080
rect 4526 4936 4582 4992
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5998 13776 6054 13832
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 6182 16088 6238 16144
rect 6274 15952 6330 16008
rect 6274 14456 6330 14512
rect 6274 14048 6330 14104
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5998 3576 6054 3632
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5446 1808 5502 1864
rect 5998 1400 6054 1456
rect 6458 9560 6514 9616
rect 6458 8472 6514 8528
rect 7286 17992 7342 18048
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 6642 5072 6698 5128
rect 6642 3440 6698 3496
rect 6826 3168 6882 3224
rect 6458 2932 6460 2952
rect 6460 2932 6512 2952
rect 6512 2932 6514 2952
rect 6458 2896 6514 2932
rect 7930 13640 7986 13696
rect 7838 9288 7894 9344
rect 7746 9016 7802 9072
rect 8022 7112 8078 7168
rect 8390 6160 8446 6216
rect 8298 4936 8354 4992
rect 8666 10920 8722 10976
rect 9034 13776 9090 13832
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9310 12280 9366 12336
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9954 13776 10010 13832
rect 9494 12280 9550 12336
rect 9218 7792 9274 7848
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 13640 10194 13696
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 9678 6704 9734 6760
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10874 9968 10930 10024
rect 11334 14592 11390 14648
rect 11242 11736 11298 11792
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5888 10838 5944
rect 10138 5752 10194 5808
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 11886 13912 11942 13968
rect 11978 12552 12034 12608
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 1536 10930 1592
rect 10322 992 10378 1048
rect 11610 3576 11666 3632
rect 11242 3304 11298 3360
rect 11978 10512 12034 10568
rect 11886 9424 11942 9480
rect 11794 3168 11850 3224
rect 11886 3032 11942 3088
rect 12254 8336 12310 8392
rect 12438 8880 12494 8936
rect 12530 3984 12586 4040
rect 12070 2896 12126 2952
rect 13266 5072 13322 5128
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 13634 5616 13690 5672
rect 12898 3440 12954 3496
rect 12806 2916 12862 2952
rect 12806 2896 12808 2916
rect 12808 2896 12860 2916
rect 12860 2896 12862 2916
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14646 14048 14702 14104
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15290 12824 15346 12880
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15750 15952 15806 16008
rect 14370 3440 14426 3496
rect 14186 1808 14242 1864
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 15842 9968 15898 10024
rect 15934 9424 15990 9480
rect 16394 12960 16450 13016
rect 16302 7792 16358 7848
rect 15750 6160 15806 6216
rect 16762 6704 16818 6760
rect 17406 13096 17462 13152
rect 17406 12688 17462 12744
rect 15198 2624 15254 2680
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14738 1128 14794 1184
rect 17314 3984 17370 4040
rect 17406 1400 17462 1456
rect 18234 8880 18290 8936
rect 20442 16088 20498 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 18602 14592 18658 14648
rect 18510 14456 18566 14512
rect 18510 12688 18566 12744
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 20442 14320 20498 14376
rect 20350 13948 20352 13968
rect 20352 13948 20404 13968
rect 20404 13948 20406 13968
rect 20350 13912 20406 13948
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 20442 12824 20498 12880
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19338 10668 19394 10704
rect 19338 10648 19340 10668
rect 19340 10648 19392 10668
rect 19392 10648 19394 10668
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 17774 2896 17830 2952
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 20350 9016 20406 9072
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20350 3440 20406 3496
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22098 13368 22154 13424
rect 22190 10512 22246 10568
rect 22374 13368 22430 13424
rect 22374 13096 22430 13152
rect 21822 3984 21878 4040
rect 22282 5616 22338 5672
rect 22834 10376 22890 10432
rect 23662 20848 23718 20904
rect 24122 23704 24178 23760
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 22616 24822 22672
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 25410 21664 25466 21720
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24766 18536 24822 18592
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24766 17448 24822 17504
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25226 16496 25282 16552
rect 24674 15408 24730 15464
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24214 13388 24270 13424
rect 24214 13368 24216 13388
rect 24216 13368 24268 13388
rect 24268 13368 24270 13388
rect 23754 12960 23810 13016
rect 23478 12688 23534 12744
rect 22926 9968 22982 10024
rect 23202 10104 23258 10160
rect 23018 9696 23074 9752
rect 20902 1944 20958 2000
rect 20626 720 20682 776
rect 23386 10240 23442 10296
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24674 9424 24730 9480
rect 25226 12280 25282 12336
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24306 8472 24362 8528
rect 24950 10260 25006 10296
rect 24950 10240 24952 10260
rect 24952 10240 25004 10260
rect 25004 10240 25006 10260
rect 24858 8336 24914 8392
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 26146 19488 26202 19544
rect 25502 10648 25558 10704
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23202 3576 23258 3632
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24674 3032 24730 3088
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23662 1128 23718 1184
rect 24674 992 24730 1048
rect 25318 8200 25374 8256
rect 27618 13912 27674 13968
rect 27618 11736 27674 11792
rect 26146 6024 26202 6080
rect 26054 5888 26110 5944
rect 25778 5072 25834 5128
rect 26146 2896 26202 2952
rect 27710 2488 27766 2544
<< metal3 >>
rect 0 27344 480 27464
rect 27520 27344 28000 27464
rect 62 26890 122 27344
rect 1577 26890 1643 26893
rect 62 26888 1643 26890
rect 62 26832 1582 26888
rect 1638 26832 1643 26888
rect 62 26830 1643 26832
rect 1577 26827 1643 26830
rect 24761 26890 24827 26893
rect 27662 26890 27722 27344
rect 24761 26888 27722 26890
rect 24761 26832 24766 26888
rect 24822 26832 27722 26888
rect 24761 26830 27722 26832
rect 24761 26827 24827 26830
rect 0 26256 480 26376
rect 27520 26256 28000 26376
rect 62 25802 122 26256
rect 1025 25802 1091 25805
rect 62 25800 1091 25802
rect 62 25744 1030 25800
rect 1086 25744 1091 25800
rect 62 25742 1091 25744
rect 1025 25739 1091 25742
rect 24209 25802 24275 25805
rect 27662 25802 27722 26256
rect 24209 25800 27722 25802
rect 24209 25744 24214 25800
rect 24270 25744 27722 25800
rect 24209 25742 27722 25744
rect 24209 25739 24275 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25396 480 25424
rect 0 25332 60 25396
rect 124 25332 480 25396
rect 0 25304 480 25332
rect 27520 25304 28000 25424
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 54 24788 60 24852
rect 124 24850 130 24852
rect 1669 24850 1735 24853
rect 124 24848 1735 24850
rect 124 24792 1674 24848
rect 1730 24792 1735 24848
rect 124 24790 1735 24792
rect 124 24788 130 24790
rect 1669 24787 1735 24790
rect 23933 24850 23999 24853
rect 27662 24850 27722 25304
rect 23933 24848 27722 24850
rect 23933 24792 23938 24848
rect 23994 24792 27722 24848
rect 23933 24790 27722 24792
rect 23933 24787 23999 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24216 480 24336
rect 27520 24308 28000 24336
rect 27520 24244 27660 24308
rect 27724 24244 28000 24308
rect 27520 24216 28000 24244
rect 62 24034 122 24216
rect 1485 24034 1551 24037
rect 62 24032 1551 24034
rect 62 23976 1490 24032
rect 1546 23976 1551 24032
rect 62 23974 1551 23976
rect 1485 23971 1551 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24117 23762 24183 23765
rect 27654 23762 27660 23764
rect 24117 23760 27660 23762
rect 24117 23704 24122 23760
rect 24178 23704 27660 23760
rect 24117 23702 27660 23704
rect 24117 23699 24183 23702
rect 27654 23700 27660 23702
rect 27724 23700 27730 23764
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 0 23128 480 23248
rect 27520 23128 28000 23248
rect 62 22674 122 23128
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 1577 22674 1643 22677
rect 62 22672 1643 22674
rect 62 22616 1582 22672
rect 1638 22616 1643 22672
rect 62 22614 1643 22616
rect 1577 22611 1643 22614
rect 24761 22674 24827 22677
rect 27662 22674 27722 23128
rect 24761 22672 27722 22674
rect 24761 22616 24766 22672
rect 24822 22616 27722 22672
rect 24761 22614 27722 22616
rect 24761 22611 24827 22614
rect 10277 22336 10597 22337
rect 0 22176 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 27520 22176 28000 22296
rect 62 21722 122 22176
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 2262 21722 2268 21724
rect 62 21662 2268 21722
rect 2262 21660 2268 21662
rect 2332 21660 2338 21724
rect 25405 21722 25471 21725
rect 27662 21722 27722 22176
rect 25405 21720 27722 21722
rect 25405 21664 25410 21720
rect 25466 21664 27722 21720
rect 25405 21662 27722 21664
rect 25405 21659 25471 21662
rect 10277 21248 10597 21249
rect 0 21088 480 21208
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 27520 21088 28000 21208
rect 62 20634 122 21088
rect 23657 20906 23723 20909
rect 27662 20906 27722 21088
rect 23657 20904 27722 20906
rect 23657 20848 23662 20904
rect 23718 20848 27722 20904
rect 23657 20846 27722 20848
rect 23657 20843 23723 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 2630 20634 2636 20636
rect 62 20574 2636 20634
rect 2630 20572 2636 20574
rect 2700 20572 2706 20636
rect 10277 20160 10597 20161
rect 0 20088 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20032 110 20088
rect 166 20032 480 20088
rect 0 20000 480 20032
rect 27520 20000 28000 20120
rect 54 19756 60 19820
rect 124 19818 130 19820
rect 1301 19818 1367 19821
rect 124 19816 1367 19818
rect 124 19760 1306 19816
rect 1362 19760 1367 19816
rect 124 19758 1367 19760
rect 124 19756 130 19758
rect 1301 19755 1367 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 26141 19546 26207 19549
rect 27662 19546 27722 20000
rect 26141 19544 27722 19546
rect 26141 19488 26146 19544
rect 26202 19488 27722 19544
rect 26141 19486 27722 19488
rect 26141 19483 26207 19486
rect 0 19048 480 19168
rect 10277 19072 10597 19073
rect 62 18594 122 19048
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19168
rect 19610 19007 19930 19008
rect 1577 18594 1643 18597
rect 62 18592 1643 18594
rect 62 18536 1582 18592
rect 1638 18536 1643 18592
rect 62 18534 1643 18536
rect 1577 18531 1643 18534
rect 24761 18594 24827 18597
rect 27662 18594 27722 19048
rect 24761 18592 27722 18594
rect 24761 18536 24766 18592
rect 24822 18536 27722 18592
rect 24761 18534 27722 18536
rect 24761 18531 24827 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 1393 18458 1459 18461
rect 62 18456 1459 18458
rect 62 18400 1398 18456
rect 1454 18400 1459 18456
rect 62 18398 1459 18400
rect 62 18080 122 18398
rect 1393 18395 1459 18398
rect 0 17960 480 18080
rect 4337 18050 4403 18053
rect 4470 18050 4476 18052
rect 4337 18048 4476 18050
rect 4337 17992 4342 18048
rect 4398 17992 4476 18048
rect 4337 17990 4476 17992
rect 4337 17987 4403 17990
rect 4470 17988 4476 17990
rect 4540 17988 4546 18052
rect 7281 18050 7347 18053
rect 7414 18050 7420 18052
rect 7281 18048 7420 18050
rect 7281 17992 7286 18048
rect 7342 17992 7420 18048
rect 7281 17990 7420 17992
rect 7281 17987 7347 17990
rect 7414 17988 7420 17990
rect 7484 17988 7490 18052
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 18080
rect 19610 17919 19930 17920
rect 238 17716 244 17780
rect 308 17778 314 17780
rect 933 17778 999 17781
rect 308 17776 999 17778
rect 308 17720 938 17776
rect 994 17720 999 17776
rect 308 17718 999 17720
rect 308 17716 314 17718
rect 933 17715 999 17718
rect 1853 17642 1919 17645
rect 62 17640 1919 17642
rect 62 17584 1858 17640
rect 1914 17584 1919 17640
rect 62 17582 1919 17584
rect 62 17128 122 17582
rect 1853 17579 1919 17582
rect 24761 17506 24827 17509
rect 27662 17506 27722 17960
rect 24761 17504 27722 17506
rect 24761 17448 24766 17504
rect 24822 17448 27722 17504
rect 24761 17446 27722 17448
rect 24761 17443 24827 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 0 17008 480 17128
rect 27520 17008 28000 17128
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 1945 16690 2011 16693
rect 2078 16690 2084 16692
rect 1945 16688 2084 16690
rect 1945 16632 1950 16688
rect 2006 16632 2084 16688
rect 1945 16630 2084 16632
rect 1945 16627 2011 16630
rect 2078 16628 2084 16630
rect 2148 16628 2154 16692
rect 25221 16554 25287 16557
rect 27662 16554 27722 17008
rect 25221 16552 27722 16554
rect 25221 16496 25226 16552
rect 25282 16496 27722 16552
rect 25221 16494 27722 16496
rect 25221 16491 25287 16494
rect 2865 16418 2931 16421
rect 62 16416 2931 16418
rect 62 16360 2870 16416
rect 2926 16360 2931 16416
rect 62 16358 2931 16360
rect 62 16040 122 16358
rect 2865 16355 2931 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 6177 16146 6243 16149
rect 20437 16146 20503 16149
rect 6177 16144 20503 16146
rect 6177 16088 6182 16144
rect 6238 16088 20442 16144
rect 20498 16088 20503 16144
rect 6177 16086 20503 16088
rect 6177 16083 6243 16086
rect 20437 16083 20503 16086
rect 0 15920 480 16040
rect 6269 16010 6335 16013
rect 15745 16010 15811 16013
rect 6269 16008 15811 16010
rect 6269 15952 6274 16008
rect 6330 15952 15750 16008
rect 15806 15952 15811 16008
rect 6269 15950 15811 15952
rect 6269 15947 6335 15950
rect 15745 15947 15811 15950
rect 27520 15920 28000 16040
rect 3969 15874 4035 15877
rect 4102 15874 4108 15876
rect 3969 15872 4108 15874
rect 3969 15816 3974 15872
rect 4030 15816 4108 15872
rect 3969 15814 4108 15816
rect 3969 15811 4035 15814
rect 4102 15812 4108 15814
rect 4172 15812 4178 15876
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 24669 15466 24735 15469
rect 27662 15466 27722 15920
rect 24669 15464 27722 15466
rect 24669 15408 24674 15464
rect 24730 15408 27722 15464
rect 24669 15406 27722 15408
rect 24669 15403 24735 15406
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 0 14832 480 14952
rect 27520 14832 28000 14952
rect 62 14514 122 14832
rect 2129 14786 2195 14789
rect 4613 14786 4679 14789
rect 2129 14784 7344 14786
rect 2129 14728 2134 14784
rect 2190 14728 4618 14784
rect 4674 14728 7344 14784
rect 2129 14726 7344 14728
rect 2129 14723 2195 14726
rect 4613 14723 4679 14726
rect 6269 14514 6335 14517
rect 62 14512 6335 14514
rect 62 14456 6274 14512
rect 6330 14456 6335 14512
rect 62 14454 6335 14456
rect 7284 14514 7344 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 11329 14650 11395 14653
rect 18597 14650 18663 14653
rect 11329 14648 18663 14650
rect 11329 14592 11334 14648
rect 11390 14592 18602 14648
rect 18658 14592 18663 14648
rect 11329 14590 18663 14592
rect 11329 14587 11395 14590
rect 18597 14587 18663 14590
rect 18505 14514 18571 14517
rect 7284 14512 18571 14514
rect 7284 14456 18510 14512
rect 18566 14456 18571 14512
rect 7284 14454 18571 14456
rect 6269 14451 6335 14454
rect 18505 14451 18571 14454
rect 20437 14378 20503 14381
rect 27662 14378 27722 14832
rect 20437 14376 27722 14378
rect 20437 14320 20442 14376
rect 20498 14320 27722 14376
rect 20437 14318 27722 14320
rect 20437 14315 20503 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6269 14106 6335 14109
rect 14641 14106 14707 14109
rect 6269 14104 14707 14106
rect 6269 14048 6274 14104
rect 6330 14048 14646 14104
rect 14702 14048 14707 14104
rect 6269 14046 14707 14048
rect 6269 14043 6335 14046
rect 14641 14043 14707 14046
rect 0 13880 480 14000
rect 11881 13970 11947 13973
rect 20345 13970 20411 13973
rect 3972 13968 20411 13970
rect 3972 13912 11886 13968
rect 11942 13912 20350 13968
rect 20406 13912 20411 13968
rect 3972 13910 20411 13912
rect 62 13698 122 13880
rect 3972 13698 4032 13910
rect 11881 13907 11947 13910
rect 20345 13907 20411 13910
rect 27520 13968 28000 14000
rect 27520 13912 27618 13968
rect 27674 13912 28000 13968
rect 27520 13880 28000 13912
rect 4337 13834 4403 13837
rect 5993 13834 6059 13837
rect 4337 13832 6059 13834
rect 4337 13776 4342 13832
rect 4398 13776 5998 13832
rect 6054 13776 6059 13832
rect 4337 13774 6059 13776
rect 4337 13771 4403 13774
rect 5993 13771 6059 13774
rect 9029 13834 9095 13837
rect 9949 13834 10015 13837
rect 9029 13832 10015 13834
rect 9029 13776 9034 13832
rect 9090 13776 9954 13832
rect 10010 13776 10015 13832
rect 9029 13774 10015 13776
rect 9029 13771 9095 13774
rect 9949 13771 10015 13774
rect 62 13638 4032 13698
rect 7925 13698 7991 13701
rect 10133 13698 10199 13701
rect 7925 13696 10199 13698
rect 7925 13640 7930 13696
rect 7986 13640 10138 13696
rect 10194 13640 10199 13696
rect 7925 13638 10199 13640
rect 7925 13635 7991 13638
rect 10133 13635 10199 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4153 13426 4219 13429
rect 22093 13426 22159 13429
rect 4153 13424 22159 13426
rect 4153 13368 4158 13424
rect 4214 13368 22098 13424
rect 22154 13368 22159 13424
rect 4153 13366 22159 13368
rect 4153 13363 4219 13366
rect 22093 13363 22159 13366
rect 22369 13426 22435 13429
rect 24209 13426 24275 13429
rect 22369 13424 24275 13426
rect 22369 13368 22374 13424
rect 22430 13368 24214 13424
rect 24270 13368 24275 13424
rect 22369 13366 24275 13368
rect 22369 13363 22435 13366
rect 24209 13363 24275 13366
rect 22096 13290 22156 13363
rect 22096 13230 27722 13290
rect 17401 13154 17467 13157
rect 22369 13154 22435 13157
rect 17401 13152 22435 13154
rect 17401 13096 17406 13152
rect 17462 13096 22374 13152
rect 22430 13096 22435 13152
rect 17401 13094 22435 13096
rect 17401 13091 17467 13094
rect 22369 13091 22435 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 16389 13018 16455 13021
rect 23749 13018 23815 13021
rect 16389 13016 23815 13018
rect 16389 12960 16394 13016
rect 16450 12960 23754 13016
rect 23810 12960 23815 13016
rect 16389 12958 23815 12960
rect 16389 12955 16455 12958
rect 23749 12955 23815 12958
rect 27662 12912 27722 13230
rect 0 12882 480 12912
rect 0 12822 9690 12882
rect 0 12792 480 12822
rect 9630 12746 9690 12822
rect 14774 12820 14780 12884
rect 14844 12882 14850 12884
rect 15285 12882 15351 12885
rect 20437 12882 20503 12885
rect 14844 12880 15351 12882
rect 14844 12824 15290 12880
rect 15346 12824 15351 12880
rect 14844 12822 15351 12824
rect 14844 12820 14850 12822
rect 15285 12819 15351 12822
rect 18278 12880 20503 12882
rect 18278 12824 20442 12880
rect 20498 12824 20503 12880
rect 18278 12822 20503 12824
rect 17401 12746 17467 12749
rect 9262 12744 17467 12746
rect 9262 12688 17406 12744
rect 17462 12688 17467 12744
rect 9262 12686 17467 12688
rect 2262 12412 2268 12476
rect 2332 12474 2338 12476
rect 4245 12474 4311 12477
rect 2332 12472 4311 12474
rect 2332 12416 4250 12472
rect 4306 12416 4311 12472
rect 2332 12414 4311 12416
rect 2332 12412 2338 12414
rect 4245 12411 4311 12414
rect 9262 12341 9322 12686
rect 17401 12683 17467 12686
rect 11973 12610 12039 12613
rect 18278 12610 18338 12822
rect 20437 12819 20503 12822
rect 27520 12792 28000 12912
rect 18505 12746 18571 12749
rect 23473 12746 23539 12749
rect 18505 12744 23539 12746
rect 18505 12688 18510 12744
rect 18566 12688 23478 12744
rect 23534 12688 23539 12744
rect 18505 12686 23539 12688
rect 18505 12683 18571 12686
rect 23473 12683 23539 12686
rect 11973 12608 18338 12610
rect 11973 12552 11978 12608
rect 12034 12552 18338 12608
rect 11973 12550 18338 12552
rect 11973 12547 12039 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 2630 12276 2636 12340
rect 2700 12338 2706 12340
rect 3509 12338 3575 12341
rect 2700 12336 3575 12338
rect 2700 12280 3514 12336
rect 3570 12280 3575 12336
rect 2700 12278 3575 12280
rect 2700 12276 2706 12278
rect 3509 12275 3575 12278
rect 4470 12276 4476 12340
rect 4540 12338 4546 12340
rect 4981 12338 5047 12341
rect 4540 12336 5047 12338
rect 4540 12280 4986 12336
rect 5042 12280 5047 12336
rect 4540 12278 5047 12280
rect 9262 12336 9371 12341
rect 9262 12280 9310 12336
rect 9366 12280 9371 12336
rect 9262 12278 9371 12280
rect 4540 12276 4546 12278
rect 4981 12275 5047 12278
rect 9305 12275 9371 12278
rect 9489 12338 9555 12341
rect 25221 12338 25287 12341
rect 9489 12336 25287 12338
rect 9489 12280 9494 12336
rect 9550 12280 25226 12336
rect 25282 12280 25287 12336
rect 9489 12278 25287 12280
rect 9489 12275 9555 12278
rect 473 12202 539 12205
rect 9630 12202 9690 12278
rect 25221 12275 25287 12278
rect 473 12200 9690 12202
rect 473 12144 478 12200
rect 534 12144 9690 12200
rect 473 12142 9690 12144
rect 473 12139 539 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11704 480 11824
rect 1301 11794 1367 11797
rect 11237 11794 11303 11797
rect 1301 11792 11303 11794
rect 1301 11736 1306 11792
rect 1362 11736 11242 11792
rect 11298 11736 11303 11792
rect 1301 11734 11303 11736
rect 1301 11731 1367 11734
rect 11237 11731 11303 11734
rect 27520 11792 28000 11824
rect 27520 11736 27618 11792
rect 27674 11736 28000 11792
rect 27520 11704 28000 11736
rect 62 11250 122 11704
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 1117 11250 1183 11253
rect 62 11248 1183 11250
rect 62 11192 1122 11248
rect 1178 11192 1183 11248
rect 62 11190 1183 11192
rect 1117 11187 1183 11190
rect 8661 10978 8727 10981
rect 9622 10978 9628 10980
rect 8661 10976 9628 10978
rect 8661 10920 8666 10976
rect 8722 10920 9628 10976
rect 8661 10918 9628 10920
rect 8661 10915 8727 10918
rect 9622 10916 9628 10918
rect 9692 10916 9698 10980
rect 5610 10912 5930 10913
rect 0 10840 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10784 386 10840
rect 442 10784 480 10840
rect 0 10752 480 10784
rect 27520 10752 28000 10872
rect 4981 10706 5047 10709
rect 19333 10706 19399 10709
rect 25497 10706 25563 10709
rect 4981 10704 13830 10706
rect 4981 10648 4986 10704
rect 5042 10648 13830 10704
rect 4981 10646 13830 10648
rect 4981 10643 5047 10646
rect 11973 10570 12039 10573
rect 62 10568 12039 10570
rect 62 10512 11978 10568
rect 12034 10512 12039 10568
rect 62 10510 12039 10512
rect 13770 10570 13830 10646
rect 19333 10704 25563 10706
rect 19333 10648 19338 10704
rect 19394 10648 25502 10704
rect 25558 10648 25563 10704
rect 19333 10646 25563 10648
rect 19333 10643 19399 10646
rect 25497 10643 25563 10646
rect 22185 10570 22251 10573
rect 27662 10570 27722 10752
rect 13770 10568 27722 10570
rect 13770 10512 22190 10568
rect 22246 10512 27722 10568
rect 13770 10510 27722 10512
rect 62 9784 122 10510
rect 11973 10507 12039 10510
rect 22185 10507 22251 10510
rect 22829 10434 22895 10437
rect 20716 10432 27722 10434
rect 20716 10376 22834 10432
rect 22890 10376 27722 10432
rect 20716 10374 27722 10376
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 4102 10100 4108 10164
rect 4172 10162 4178 10164
rect 5165 10162 5231 10165
rect 20716 10162 20776 10374
rect 22829 10371 22895 10374
rect 23381 10298 23447 10301
rect 24945 10298 25011 10301
rect 23381 10296 25011 10298
rect 23381 10240 23386 10296
rect 23442 10240 24950 10296
rect 25006 10240 25011 10296
rect 23381 10238 25011 10240
rect 23381 10235 23447 10238
rect 24945 10235 25011 10238
rect 4172 10160 20776 10162
rect 4172 10104 5170 10160
rect 5226 10104 20776 10160
rect 4172 10102 20776 10104
rect 23197 10162 23263 10165
rect 23197 10160 23306 10162
rect 23197 10104 23202 10160
rect 23258 10104 23306 10160
rect 4172 10100 4178 10102
rect 5165 10099 5231 10102
rect 23197 10099 23306 10104
rect 10869 10026 10935 10029
rect 15837 10026 15903 10029
rect 10869 10024 15903 10026
rect 10869 9968 10874 10024
rect 10930 9968 15842 10024
rect 15898 9968 15903 10024
rect 10869 9966 15903 9968
rect 10869 9963 10935 9966
rect 15837 9963 15903 9966
rect 22686 9964 22692 10028
rect 22756 10026 22762 10028
rect 22921 10026 22987 10029
rect 22756 10024 22987 10026
rect 22756 9968 22926 10024
rect 22982 9968 22987 10024
rect 22756 9966 22987 9968
rect 22756 9964 22762 9966
rect 22921 9963 22987 9966
rect 5610 9824 5930 9825
rect 0 9664 480 9784
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 23013 9754 23079 9757
rect 23246 9754 23306 10099
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 27662 9784 27722 10374
rect 24277 9759 24597 9760
rect 23013 9752 23306 9754
rect 23013 9696 23018 9752
rect 23074 9696 23306 9752
rect 23013 9694 23306 9696
rect 23013 9691 23079 9694
rect 27520 9664 28000 9784
rect 1761 9618 1827 9621
rect 4613 9618 4679 9621
rect 6453 9618 6519 9621
rect 1761 9616 6519 9618
rect 1761 9560 1766 9616
rect 1822 9560 4618 9616
rect 4674 9560 6458 9616
rect 6514 9560 6519 9616
rect 1761 9558 6519 9560
rect 1761 9555 1827 9558
rect 4613 9555 4679 9558
rect 6453 9555 6519 9558
rect 9622 9420 9628 9484
rect 9692 9482 9698 9484
rect 11881 9482 11947 9485
rect 9692 9480 11947 9482
rect 9692 9424 11886 9480
rect 11942 9424 11947 9480
rect 9692 9422 11947 9424
rect 9692 9420 9698 9422
rect 11881 9419 11947 9422
rect 15929 9482 15995 9485
rect 24669 9482 24735 9485
rect 15929 9480 24735 9482
rect 15929 9424 15934 9480
rect 15990 9424 24674 9480
rect 24730 9424 24735 9480
rect 15929 9422 24735 9424
rect 15929 9419 15995 9422
rect 24669 9419 24735 9422
rect 2078 9284 2084 9348
rect 2148 9346 2154 9348
rect 7833 9346 7899 9349
rect 2148 9344 7899 9346
rect 2148 9288 7838 9344
rect 7894 9288 7899 9344
rect 2148 9286 7899 9288
rect 2148 9284 2154 9286
rect 7833 9283 7899 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 7741 9074 7807 9077
rect 20345 9074 20411 9077
rect 62 9072 20411 9074
rect 62 9016 7746 9072
rect 7802 9016 20350 9072
rect 20406 9016 20411 9072
rect 62 9014 20411 9016
rect 62 8832 122 9014
rect 7741 9011 7807 9014
rect 20345 9011 20411 9014
rect 12433 8938 12499 8941
rect 18229 8938 18295 8941
rect 12433 8936 18295 8938
rect 12433 8880 12438 8936
rect 12494 8880 18234 8936
rect 18290 8880 18295 8936
rect 12433 8878 18295 8880
rect 12433 8875 12499 8878
rect 18229 8875 18295 8878
rect 0 8712 480 8832
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8832
rect 24277 8671 24597 8672
rect 6453 8530 6519 8533
rect 24301 8530 24367 8533
rect 27662 8530 27722 8712
rect 6453 8528 27722 8530
rect 6453 8472 6458 8528
rect 6514 8472 24306 8528
rect 24362 8472 27722 8528
rect 6453 8470 27722 8472
rect 6453 8467 6519 8470
rect 24301 8467 24367 8470
rect 12249 8394 12315 8397
rect 24853 8394 24919 8397
rect 12249 8392 24919 8394
rect 12249 8336 12254 8392
rect 12310 8336 24858 8392
rect 24914 8336 24919 8392
rect 12249 8334 24919 8336
rect 12249 8331 12315 8334
rect 24853 8331 24919 8334
rect 289 8258 355 8261
rect 62 8256 355 8258
rect 62 8200 294 8256
rect 350 8200 355 8256
rect 62 8198 355 8200
rect 62 7744 122 8198
rect 289 8195 355 8198
rect 2446 8196 2452 8260
rect 2516 8258 2522 8260
rect 2773 8258 2839 8261
rect 2516 8256 2839 8258
rect 2516 8200 2778 8256
rect 2834 8200 2839 8256
rect 2516 8198 2839 8200
rect 2516 8196 2522 8198
rect 2773 8195 2839 8198
rect 25313 8258 25379 8261
rect 25313 8256 27722 8258
rect 25313 8200 25318 8256
rect 25374 8200 27722 8256
rect 25313 8198 27722 8200
rect 25313 8195 25379 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 9213 7850 9279 7853
rect 16297 7850 16363 7853
rect 9213 7848 16363 7850
rect 9213 7792 9218 7848
rect 9274 7792 16302 7848
rect 16358 7792 16363 7848
rect 9213 7790 16363 7792
rect 9213 7787 9279 7790
rect 16297 7787 16363 7790
rect 27662 7744 27722 8198
rect 0 7624 480 7744
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7744
rect 24277 7583 24597 7584
rect 7414 7108 7420 7172
rect 7484 7170 7490 7172
rect 8017 7170 8083 7173
rect 7484 7168 8083 7170
rect 7484 7112 8022 7168
rect 8078 7112 8083 7168
rect 7484 7110 8083 7112
rect 7484 7108 7490 7110
rect 8017 7107 8083 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 9673 6762 9739 6765
rect 16757 6762 16823 6765
rect 9673 6760 16823 6762
rect 9673 6704 9678 6760
rect 9734 6704 16762 6760
rect 16818 6704 16823 6760
rect 9673 6702 16823 6704
rect 9673 6699 9739 6702
rect 16757 6699 16823 6702
rect 0 6624 480 6656
rect 0 6568 110 6624
rect 166 6568 480 6624
rect 0 6536 480 6568
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6656
rect 24277 6495 24597 6496
rect 8385 6218 8451 6221
rect 15745 6218 15811 6221
rect 8385 6216 15811 6218
rect 8385 6160 8390 6216
rect 8446 6160 15750 6216
rect 15806 6160 15811 6216
rect 8385 6158 15811 6160
rect 8385 6155 8451 6158
rect 15745 6155 15811 6158
rect 1945 6082 2011 6085
rect 4429 6082 4495 6085
rect 1945 6080 4495 6082
rect 1945 6024 1950 6080
rect 2006 6024 4434 6080
rect 4490 6024 4495 6080
rect 1945 6022 4495 6024
rect 1945 6019 2011 6022
rect 4429 6019 4495 6022
rect 26141 6082 26207 6085
rect 27662 6082 27722 6536
rect 26141 6080 27722 6082
rect 26141 6024 26146 6080
rect 26202 6024 27722 6080
rect 26141 6022 27722 6024
rect 26141 6019 26207 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 10777 5946 10843 5949
rect 10734 5944 10843 5946
rect 10734 5888 10782 5944
rect 10838 5888 10843 5944
rect 10734 5883 10843 5888
rect 26049 5946 26115 5949
rect 26049 5944 27722 5946
rect 26049 5888 26054 5944
rect 26110 5888 27722 5944
rect 26049 5886 27722 5888
rect 26049 5883 26115 5886
rect 10133 5810 10199 5813
rect 10734 5810 10794 5883
rect 10133 5808 10794 5810
rect 10133 5752 10138 5808
rect 10194 5752 10794 5808
rect 10133 5750 10794 5752
rect 10133 5747 10199 5750
rect 27662 5704 27722 5886
rect 0 5672 480 5704
rect 0 5616 110 5672
rect 166 5616 480 5672
rect 0 5584 480 5616
rect 13629 5674 13695 5677
rect 22277 5674 22343 5677
rect 13629 5672 22343 5674
rect 13629 5616 13634 5672
rect 13690 5616 22282 5672
rect 22338 5616 22343 5672
rect 13629 5614 22343 5616
rect 13629 5611 13695 5614
rect 22277 5611 22343 5614
rect 27520 5584 28000 5704
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 1485 5130 1551 5133
rect 62 5128 1551 5130
rect 62 5072 1490 5128
rect 1546 5072 1551 5128
rect 62 5070 1551 5072
rect 62 4616 122 5070
rect 1485 5067 1551 5070
rect 6637 5130 6703 5133
rect 13261 5130 13327 5133
rect 6637 5128 13327 5130
rect 6637 5072 6642 5128
rect 6698 5072 13266 5128
rect 13322 5072 13327 5128
rect 6637 5070 13327 5072
rect 6637 5067 6703 5070
rect 13261 5067 13327 5070
rect 25773 5130 25839 5133
rect 25773 5128 27722 5130
rect 25773 5072 25778 5128
rect 25834 5072 27722 5128
rect 25773 5070 27722 5072
rect 25773 5067 25839 5070
rect 4521 4994 4587 4997
rect 8293 4994 8359 4997
rect 4521 4992 8359 4994
rect 4521 4936 4526 4992
rect 4582 4936 8298 4992
rect 8354 4936 8359 4992
rect 4521 4934 8359 4936
rect 4521 4931 4587 4934
rect 8293 4931 8359 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 27662 4616 27722 5070
rect 0 4496 480 4616
rect 27520 4496 28000 4616
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 12525 4042 12591 4045
rect 4110 4040 12591 4042
rect 4110 3984 12530 4040
rect 12586 3984 12591 4040
rect 4110 3982 12591 3984
rect 2129 3906 2195 3909
rect 4110 3906 4170 3982
rect 12525 3979 12591 3982
rect 17309 4042 17375 4045
rect 21817 4042 21883 4045
rect 17309 4040 21883 4042
rect 17309 3984 17314 4040
rect 17370 3984 21822 4040
rect 21878 3984 21883 4040
rect 17309 3982 21883 3984
rect 17309 3979 17375 3982
rect 21817 3979 21883 3982
rect 2129 3904 4170 3906
rect 2129 3848 2134 3904
rect 2190 3848 4170 3904
rect 2129 3846 4170 3848
rect 2129 3843 2195 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3785 3634 3851 3637
rect 5993 3634 6059 3637
rect 11605 3634 11671 3637
rect 3785 3632 4170 3634
rect 3785 3576 3790 3632
rect 3846 3576 4170 3632
rect 3785 3574 4170 3576
rect 3785 3571 3851 3574
rect 0 3496 480 3528
rect 0 3440 18 3496
rect 74 3440 480 3496
rect 0 3408 480 3440
rect 4110 3498 4170 3574
rect 5993 3632 11671 3634
rect 5993 3576 5998 3632
rect 6054 3576 11610 3632
rect 11666 3576 11671 3632
rect 5993 3574 11671 3576
rect 5993 3571 6059 3574
rect 11605 3571 11671 3574
rect 22686 3572 22692 3636
rect 22756 3634 22762 3636
rect 23197 3634 23263 3637
rect 22756 3632 23263 3634
rect 22756 3576 23202 3632
rect 23258 3576 23263 3632
rect 22756 3574 23263 3576
rect 22756 3572 22762 3574
rect 23197 3571 23263 3574
rect 6637 3498 6703 3501
rect 12893 3498 12959 3501
rect 4110 3438 6056 3498
rect 5996 3362 6056 3438
rect 6637 3496 12959 3498
rect 6637 3440 6642 3496
rect 6698 3440 12898 3496
rect 12954 3440 12959 3496
rect 6637 3438 12959 3440
rect 6637 3435 6703 3438
rect 12893 3435 12959 3438
rect 14365 3498 14431 3501
rect 20345 3498 20411 3501
rect 14365 3496 20411 3498
rect 14365 3440 14370 3496
rect 14426 3440 20350 3496
rect 20406 3440 20411 3496
rect 14365 3438 20411 3440
rect 14365 3435 14431 3438
rect 20345 3435 20411 3438
rect 27520 3408 28000 3528
rect 11237 3362 11303 3365
rect 5996 3360 11303 3362
rect 5996 3304 11242 3360
rect 11298 3304 11303 3360
rect 5996 3302 11303 3304
rect 11237 3299 11303 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2129 3226 2195 3229
rect 2446 3226 2452 3228
rect 2129 3224 2452 3226
rect 2129 3168 2134 3224
rect 2190 3168 2452 3224
rect 2129 3166 2452 3168
rect 2129 3163 2195 3166
rect 2446 3164 2452 3166
rect 2516 3164 2522 3228
rect 6821 3226 6887 3229
rect 11789 3226 11855 3229
rect 6821 3224 11855 3226
rect 6821 3168 6826 3224
rect 6882 3168 11794 3224
rect 11850 3168 11855 3224
rect 6821 3166 11855 3168
rect 6821 3163 6887 3166
rect 11789 3163 11855 3166
rect 11881 3090 11947 3093
rect 24669 3090 24735 3093
rect 11881 3088 24735 3090
rect 11881 3032 11886 3088
rect 11942 3032 24674 3088
rect 24730 3032 24735 3088
rect 11881 3030 24735 3032
rect 11881 3027 11947 3030
rect 24669 3027 24735 3030
rect 6453 2954 6519 2957
rect 12065 2954 12131 2957
rect 6453 2952 12131 2954
rect 6453 2896 6458 2952
rect 6514 2896 12070 2952
rect 12126 2896 12131 2952
rect 6453 2894 12131 2896
rect 6453 2891 6519 2894
rect 12065 2891 12131 2894
rect 12801 2954 12867 2957
rect 17769 2954 17835 2957
rect 12801 2952 17835 2954
rect 12801 2896 12806 2952
rect 12862 2896 17774 2952
rect 17830 2896 17835 2952
rect 12801 2894 17835 2896
rect 12801 2891 12867 2894
rect 17769 2891 17835 2894
rect 26141 2954 26207 2957
rect 27662 2954 27722 3408
rect 26141 2952 27722 2954
rect 26141 2896 26146 2952
rect 26202 2896 27722 2952
rect 26141 2894 27722 2896
rect 26141 2891 26207 2894
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 14774 2620 14780 2684
rect 14844 2682 14850 2684
rect 15193 2682 15259 2685
rect 14844 2680 15259 2682
rect 14844 2624 15198 2680
rect 15254 2624 15259 2680
rect 14844 2622 15259 2624
rect 14844 2620 14850 2622
rect 15193 2619 15259 2622
rect 0 2548 480 2576
rect 0 2484 60 2548
rect 124 2484 480 2548
rect 0 2456 480 2484
rect 27520 2544 28000 2576
rect 27520 2488 27710 2544
rect 27766 2488 28000 2544
rect 27520 2456 28000 2488
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 20897 2002 20963 2005
rect 20897 2000 27722 2002
rect 20897 1944 20902 2000
rect 20958 1944 27722 2000
rect 20897 1942 27722 1944
rect 20897 1939 20963 1942
rect 5441 1866 5507 1869
rect 14181 1866 14247 1869
rect 5441 1864 14247 1866
rect 5441 1808 5446 1864
rect 5502 1808 14186 1864
rect 14242 1808 14247 1864
rect 5441 1806 14247 1808
rect 5441 1803 5507 1806
rect 14181 1803 14247 1806
rect 1945 1594 2011 1597
rect 10869 1594 10935 1597
rect 1945 1592 10935 1594
rect 1945 1536 1950 1592
rect 2006 1536 10874 1592
rect 10930 1536 10935 1592
rect 1945 1534 10935 1536
rect 1945 1531 2011 1534
rect 10869 1531 10935 1534
rect 27662 1488 27722 1942
rect 0 1460 480 1488
rect 0 1396 60 1460
rect 124 1396 480 1460
rect 0 1368 480 1396
rect 5993 1458 6059 1461
rect 17401 1458 17467 1461
rect 5993 1456 17467 1458
rect 5993 1400 5998 1456
rect 6054 1400 17406 1456
rect 17462 1400 17467 1456
rect 5993 1398 17467 1400
rect 5993 1395 6059 1398
rect 17401 1395 17467 1398
rect 27520 1368 28000 1488
rect 14733 1186 14799 1189
rect 23657 1186 23723 1189
rect 14733 1184 23723 1186
rect 14733 1128 14738 1184
rect 14794 1128 23662 1184
rect 23718 1128 23723 1184
rect 14733 1126 23723 1128
rect 14733 1123 14799 1126
rect 23657 1123 23723 1126
rect 1853 1050 1919 1053
rect 62 1048 1919 1050
rect 62 992 1858 1048
rect 1914 992 1919 1048
rect 62 990 1919 992
rect 62 536 122 990
rect 1853 987 1919 990
rect 10317 1050 10383 1053
rect 24669 1050 24735 1053
rect 10317 1048 24735 1050
rect 10317 992 10322 1048
rect 10378 992 24674 1048
rect 24730 992 24735 1048
rect 10317 990 24735 992
rect 10317 987 10383 990
rect 24669 987 24735 990
rect 20621 778 20687 781
rect 20621 776 27722 778
rect 20621 720 20626 776
rect 20682 720 27722 776
rect 20621 718 27722 720
rect 20621 715 20687 718
rect 27662 536 27722 718
rect 0 416 480 536
rect 27520 416 28000 536
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 60 25332 124 25396
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 60 24788 124 24852
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 27660 24244 27724 24308
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 27660 23700 27724 23764
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 2268 21660 2332 21724
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 2636 20572 2700 20636
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 60 19756 124 19820
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 4476 17988 4540 18052
rect 7420 17988 7484 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 244 17716 308 17780
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 2084 16628 2148 16692
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 4108 15812 4172 15876
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 14780 12820 14844 12884
rect 2268 12412 2332 12476
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 2636 12276 2700 12340
rect 4476 12276 4540 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 9628 10916 9692 10980
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 4108 10100 4172 10164
rect 22692 9964 22756 10028
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 9628 9420 9692 9484
rect 2084 9284 2148 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 2452 8196 2516 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 7420 7108 7484 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 22692 3572 22756 3636
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 2452 3164 2516 3228
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 14780 2620 14844 2684
rect 60 2484 124 2548
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 60 1396 124 1460
<< metal4 >>
rect 59 25396 125 25397
rect 59 25332 60 25396
rect 124 25332 125 25396
rect 59 25331 125 25332
rect 62 24853 122 25331
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 59 24852 125 24853
rect 59 24788 60 24852
rect 124 24788 125 24852
rect 59 24787 125 24788
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 2267 21724 2333 21725
rect 2267 21660 2268 21724
rect 2332 21660 2333 21724
rect 2267 21659 2333 21660
rect 59 19820 125 19821
rect 59 19756 60 19820
rect 124 19756 125 19820
rect 59 19755 125 19756
rect 62 2549 122 19755
rect 243 17780 309 17781
rect 243 17716 244 17780
rect 308 17716 309 17780
rect 243 17715 309 17716
rect 59 2548 125 2549
rect 59 2484 60 2548
rect 124 2484 125 2548
rect 59 2483 125 2484
rect 59 1460 125 1461
rect 59 1396 60 1460
rect 124 1458 125 1460
rect 246 1458 306 17715
rect 2083 16692 2149 16693
rect 2083 16628 2084 16692
rect 2148 16628 2149 16692
rect 2083 16627 2149 16628
rect 2086 9349 2146 16627
rect 2270 12477 2330 21659
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 2635 20636 2701 20637
rect 2635 20572 2636 20636
rect 2700 20572 2701 20636
rect 2635 20571 2701 20572
rect 2267 12476 2333 12477
rect 2267 12412 2268 12476
rect 2332 12412 2333 12476
rect 2267 12411 2333 12412
rect 2638 12341 2698 20571
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 4475 18052 4541 18053
rect 4475 17988 4476 18052
rect 4540 17988 4541 18052
rect 4475 17987 4541 17988
rect 4107 15876 4173 15877
rect 4107 15812 4108 15876
rect 4172 15812 4173 15876
rect 4107 15811 4173 15812
rect 2635 12340 2701 12341
rect 2635 12276 2636 12340
rect 2700 12276 2701 12340
rect 2635 12275 2701 12276
rect 4110 10165 4170 15811
rect 4478 12341 4538 17987
rect 5610 17440 5931 18464
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 7419 18052 7485 18053
rect 7419 17988 7420 18052
rect 7484 17988 7485 18052
rect 7419 17987 7485 17988
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 4475 12340 4541 12341
rect 4475 12276 4476 12340
rect 4540 12276 4541 12340
rect 4475 12275 4541 12276
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 4107 10164 4173 10165
rect 4107 10100 4108 10164
rect 4172 10100 4173 10164
rect 4107 10099 4173 10100
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 2083 9348 2149 9349
rect 2083 9284 2084 9348
rect 2148 9284 2149 9348
rect 2083 9283 2149 9284
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 2451 8260 2517 8261
rect 2451 8196 2452 8260
rect 2516 8196 2517 8260
rect 2451 8195 2517 8196
rect 2454 3229 2514 8195
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 7422 7173 7482 17987
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14779 12884 14845 12885
rect 14779 12820 14780 12884
rect 14844 12820 14845 12884
rect 14779 12819 14845 12820
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 9627 10980 9693 10981
rect 9627 10916 9628 10980
rect 9692 10916 9693 10980
rect 9627 10915 9693 10916
rect 9630 9485 9690 10915
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 9627 9484 9693 9485
rect 9627 9420 9628 9484
rect 9692 9420 9693 9484
rect 9627 9419 9693 9420
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 7419 7172 7485 7173
rect 7419 7108 7420 7172
rect 7484 7108 7485 7172
rect 7419 7107 7485 7108
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 2451 3228 2517 3229
rect 2451 3164 2452 3228
rect 2516 3164 2517 3228
rect 2451 3163 2517 3164
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14782 2685 14842 12819
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14779 2684 14845 2685
rect 14779 2620 14780 2684
rect 14844 2620 14845 2684
rect 14779 2619 14845 2620
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 27659 24308 27725 24309
rect 27659 24244 27660 24308
rect 27724 24244 27725 24308
rect 27659 24243 27725 24244
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 27662 23765 27722 24243
rect 27659 23764 27725 23765
rect 27659 23700 27660 23764
rect 27724 23700 27725 23764
rect 27659 23699 27725 23700
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 22691 10028 22757 10029
rect 22691 9964 22692 10028
rect 22756 9964 22757 10028
rect 22691 9963 22757 9964
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 22694 3637 22754 9963
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 22691 3636 22757 3637
rect 22691 3572 22692 3636
rect 22756 3572 22757 3636
rect 22691 3571 22757 3572
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 124 1398 306 1458
rect 124 1396 125 1398
rect 59 1395 125 1396
use scs8hd_decap_3  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_1  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_25
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3772 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_44 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_45
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _085_
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_4_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_65
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_89
timestamp 1586364061
transform 1 0 9292 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_93
timestamp 1586364061
transform 1 0 9660 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9476 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_106
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_112
timestamp 1586364061
transform 1 0 11408 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_112 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__C
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_nor2_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_136
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_139
timestamp 1586364061
transform 1 0 13892 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _084_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_144
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _242_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_156 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 406 592
use scs8hd_or3_4  _163_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_165
timestamp 1586364061
transform 1 0 16284 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_161
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_165
timestamp 1586364061
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_161
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16468 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_178
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor4_4  _185_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18124 0 1 2720
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_1_202
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_202
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_198
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 19872 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_231
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_227
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_237
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_233
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_241
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_254
timestamp 1586364061
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_258
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_266
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_269
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_270 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25944 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_276
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_10
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_71
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_119
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 406 592
use scs8hd_or3_4  _099_
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_136
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_140
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 406 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 16468 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 19872 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_212
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21068 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_219
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_232 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_2_244
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_247
timestamp 1586364061
transform 1 0 23828 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_257
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_269
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_26
timestamp 1586364061
transform 1 0 3496 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_30
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_70
timestamp 1586364061
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8280 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_108
timestamp 1586364061
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_112
timestamp 1586364061
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_116
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 406 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_163
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 21804 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25576 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_262
timestamp 1586364061
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_273
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_46
timestamp 1586364061
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_88
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_136
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_1  _112_
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_146
timestamp 1586364061
transform 1 0 14536 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_164
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 18124 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 17940 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 17572 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22172 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_231
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_243
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_260
timestamp 1586364061
transform 1 0 25024 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_272
timestamp 1586364061
transform 1 0 26128 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_22
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_26
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_107
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_111
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_115
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_119
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_132
timestamp 1586364061
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_136
timestamp 1586364061
transform 1 0 13616 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _187_
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__C
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_149
timestamp 1586364061
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_153
timestamp 1586364061
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_166
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 406 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 18952 0 1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_211
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21620 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_215
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_219
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_260
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_264
timestamp 1586364061
transform 1 0 25392 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_268
timestamp 1586364061
transform 1 0 25760 0 1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_5_276
timestamp 1586364061
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_6
timestamp 1586364061
transform 1 0 1656 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_13
timestamp 1586364061
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_10
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_22
timestamp 1586364061
transform 1 0 3128 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_buf_1  _103_
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_37
timestamp 1586364061
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _100_
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_decap_3  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__148__B
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_88
timestamp 1586364061
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_84
timestamp 1586364061
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 8832 0 1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 5984
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10948 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_118
timestamp 1586364061
transform 1 0 11960 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_124
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_135
timestamp 1586364061
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_139
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_4  FILLER_7_136
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_148
timestamp 1586364061
transform 1 0 14720 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_157
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 1050 592
use scs8hd_or3_4  _153_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__145__C
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 17296 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 314 592
use scs8hd_or3_4  _145_
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_182
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 20792 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_203
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_207
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_211
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_212
timestamp 1586364061
transform 1 0 20608 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_221
timestamp 1586364061
transform 1 0 21436 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 21068 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_229
timestamp 1586364061
transform 1 0 22172 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_233
timestamp 1586364061
transform 1 0 22540 0 1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_240
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_248
timestamp 1586364061
transform 1 0 23920 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23736 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23736 0 1 5984
box -38 -48 866 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_259
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_255
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_259
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_7_271
timestamp 1586364061
transform 1 0 26036 0 1 5984
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_22
timestamp 1586364061
transform 1 0 3128 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_26
timestamp 1586364061
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_29
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_49
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _148_
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_66
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 406 592
use scs8hd_conb_1  _217_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12328 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_113
timestamp 1586364061
transform 1 0 11500 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _126_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_131
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__D
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_157
timestamp 1586364061
transform 1 0 15548 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_161
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_182
timestamp 1586364061
transform 1 0 17848 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_193
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21068 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_226
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_230
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 22632 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23920 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_247
timestamp 1586364061
transform 1 0 23828 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 866 592
use scs8hd_fill_1  FILLER_8_250
timestamp 1586364061
transform 1 0 24104 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_260
timestamp 1586364061
transform 1 0 25024 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_19
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_42
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_46
timestamp 1586364061
transform 1 0 5336 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_71
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_75
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_79
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 590 592
use scs8hd_inv_8  _188_
timestamp 1586364061
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _128_
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 314 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__171__C
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_151
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _090_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_nor4_4  _182_
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_212
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_216
timestamp 1586364061
transform 1 0 20976 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_231
timestamp 1586364061
transform 1 0 22356 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_235
timestamp 1586364061
transform 1 0 22724 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 314 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 25484 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_261
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_273
timestamp 1586364061
transform 1 0 26220 0 1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_81
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_86
timestamp 1586364061
transform 1 0 9016 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_136
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_144
timestamp 1586364061
transform 1 0 14352 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _171_
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 16008 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_185
timestamp 1586364061
transform 1 0 18124 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__D
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_206
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 1050 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21068 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21528 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_220
timestamp 1586364061
transform 1 0 21344 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_224
timestamp 1586364061
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_258
timestamp 1586364061
transform 1 0 24840 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_270
timestamp 1586364061
transform 1 0 25944 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  FILLER_11_9
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 314 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_32
timestamp 1586364061
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_36
timestamp 1586364061
transform 1 0 4416 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_40
timestamp 1586364061
transform 1 0 4784 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_71
timestamp 1586364061
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8832 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_75
timestamp 1586364061
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_79
timestamp 1586364061
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_99
timestamp 1586364061
transform 1 0 10212 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_151
timestamp 1586364061
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_155
timestamp 1586364061
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_168
timestamp 1586364061
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_172
timestamp 1586364061
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_176
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 406 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_nor4_4  _180_
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__C
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_187
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_191
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_229
timestamp 1586364061
transform 1 0 22172 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22724 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_233
timestamp 1586364061
transform 1 0 22540 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_241
timestamp 1586364061
transform 1 0 23276 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 25944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_268
timestamp 1586364061
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_272
timestamp 1586364061
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 1050 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_18
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_26
timestamp 1586364061
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_36
timestamp 1586364061
transform 1 0 4416 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_42
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_6  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_136
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_140
timestamp 1586364061
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_144
timestamp 1586364061
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_152
timestamp 1586364061
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_160
timestamp 1586364061
transform 1 0 15824 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 16192 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__D
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_210
timestamp 1586364061
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20976 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_219
timestamp 1586364061
transform 1 0 21252 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_225
timestamp 1586364061
transform 1 0 21804 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_238
timestamp 1586364061
transform 1 0 23000 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_244
timestamp 1586364061
transform 1 0 23552 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_256
timestamp 1586364061
transform 1 0 24656 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_8  FILLER_12_267
timestamp 1586364061
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_12
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_34
timestamp 1586364061
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_38
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_41
timestamp 1586364061
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_46
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 314 592
use scs8hd_nor2_4  _147_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_58
timestamp 1586364061
transform 1 0 6440 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_77
timestamp 1586364061
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_96
timestamp 1586364061
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_96
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_107
timestamp 1586364061
transform 1 0 10948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_104
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_100
timestamp 1586364061
transform 1 0 10304 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_100
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 12512 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_118
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_128
timestamp 1586364061
transform 1 0 12880 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_131
timestamp 1586364061
transform 1 0 13156 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_127
timestamp 1586364061
transform 1 0 12788 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 866 592
use scs8hd_fill_1  FILLER_14_150
timestamp 1586364061
transform 1 0 14904 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_6  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_13_148
timestamp 1586364061
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_144
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_152
timestamp 1586364061
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_167
timestamp 1586364061
transform 1 0 16468 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_176
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__B
timestamp 1586364061
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__C
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_nor4_4  _172_
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 1602 592
use scs8hd_nor4_4  _175_
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_194
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_198
timestamp 1586364061
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21620 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_226
timestamp 1586364061
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_230
timestamp 1586364061
transform 1 0 22264 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_235
timestamp 1586364061
transform 1 0 22724 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22540 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23460 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24196 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_264
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_256
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_276
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_14
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5888 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_50
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_54
timestamp 1586364061
transform 1 0 6072 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_58
timestamp 1586364061
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_69
timestamp 1586364061
transform 1 0 7452 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_112
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 590 592
use scs8hd_fill_1  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13064 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_127
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_141
timestamp 1586364061
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_145
timestamp 1586364061
transform 1 0 14444 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_151
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__173__C
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__D
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_168
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_199
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_231
timestamp 1586364061
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_235
timestamp 1586364061
transform 1 0 22724 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_261
timestamp 1586364061
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_268
timestamp 1586364061
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_272
timestamp 1586364061
transform 1 0 26128 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_276
timestamp 1586364061
transform 1 0 26496 0 1 10336
box -38 -48 130 592
use scs8hd_conb_1  _215_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_30
timestamp 1586364061
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_58
timestamp 1586364061
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_6  FILLER_16_64
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_16_70
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_118
timestamp 1586364061
transform 1 0 11960 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13064 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_126
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _173_
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 1602 592
use scs8hd_decap_8  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_173
timestamp 1586364061
transform 1 0 17020 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_191
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_195
timestamp 1586364061
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_199
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_210
timestamp 1586364061
transform 1 0 20424 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20976 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_225
timestamp 1586364061
transform 1 0 21804 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_229
timestamp 1586364061
transform 1 0 22172 0 -1 11424
box -38 -48 406 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 23736 0 -1 11424
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_255
timestamp 1586364061
transform 1 0 24564 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_266
timestamp 1586364061
transform 1 0 25576 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_274
timestamp 1586364061
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 1050 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3680 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_24
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_41
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_71
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 406 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_77
timestamp 1586364061
transform 1 0 8188 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_81
timestamp 1586364061
transform 1 0 8556 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _108_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_140
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_152
timestamp 1586364061
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_169
timestamp 1586364061
transform 1 0 16652 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18216 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_214
timestamp 1586364061
transform 1 0 20792 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21528 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_218
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_231
timestamp 1586364061
transform 1 0 22356 0 1 11424
box -38 -48 590 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_237
timestamp 1586364061
transform 1 0 22908 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_240
timestamp 1586364061
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_254
timestamp 1586364061
transform 1 0 24472 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_266
timestamp 1586364061
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_270
timestamp 1586364061
transform 1 0 25944 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_276
timestamp 1586364061
transform 1 0 26496 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_7
timestamp 1586364061
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_46
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_59
timestamp 1586364061
transform 1 0 6532 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_71
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_right_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11960 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_18_121
timestamp 1586364061
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_140
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_144
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_150
timestamp 1586364061
transform 1 0 14904 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_163
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_167
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_179
timestamp 1586364061
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_192
timestamp 1586364061
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_196
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_200
timestamp 1586364061
transform 1 0 19504 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_18_206
timestamp 1586364061
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 21160 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 23460 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_4  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_8
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_23
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_19
timestamp 1586364061
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4784 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_36
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_40
timestamp 1586364061
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_53
timestamp 1586364061
transform 1 0 5980 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_61
timestamp 1586364061
transform 1 0 6716 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_65
timestamp 1586364061
transform 1 0 7084 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_73
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_88
timestamp 1586364061
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 10120 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_96
timestamp 1586364061
transform 1 0 9936 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_92
timestamp 1586364061
transform 1 0 9568 0 1 12512
box -38 -48 406 592
use scs8hd_decap_4  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_101
timestamp 1586364061
transform 1 0 10396 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_99
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_120
timestamp 1586364061
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_right_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11132 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_131
timestamp 1586364061
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1050 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_1  FILLER_20_150
timestamp 1586364061
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_19_146
timestamp 1586364061
transform 1 0 14536 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__C
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_156
timestamp 1586364061
transform 1 0 15456 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_152
timestamp 1586364061
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_169
timestamp 1586364061
transform 1 0 16652 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_166
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_170
timestamp 1586364061
transform 1 0 16744 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 17020 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use scs8hd_decap_8  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_203
timestamp 1586364061
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_199
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19964 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_213
timestamp 1586364061
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_209
timestamp 1586364061
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20148 0 1 12512
box -38 -48 866 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 866 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 21160 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_216
timestamp 1586364061
transform 1 0 20976 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_8  FILLER_20_236
timestamp 1586364061
transform 1 0 22816 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_237
timestamp 1586364061
transform 1 0 22908 0 1 12512
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_233
timestamp 1586364061
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_247
timestamp 1586364061
transform 1 0 23828 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_4  FILLER_19_249
timestamp 1586364061
transform 1 0 24012 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_19_243
timestamp 1586364061
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_259
timestamp 1586364061
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_263
timestamp 1586364061
transform 1 0 25300 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_275
timestamp 1586364061
transform 1 0 26404 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _156_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_55
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_75
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_79
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_85
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_89
timestamp 1586364061
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_104
timestamp 1586364061
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__102__C
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_108
timestamp 1586364061
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_140
timestamp 1586364061
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_right_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 14352 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_155
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use scs8hd_or3_4  _116_
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_172
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 406 592
use scs8hd_decap_4  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 406 592
use scs8hd_buf_1  _178_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_187
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_191
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_195
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_205
timestamp 1586364061
transform 1 0 19964 0 1 13600
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21528 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21896 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_216
timestamp 1586364061
transform 1 0 20976 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_224
timestamp 1586364061
transform 1 0 21712 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_228
timestamp 1586364061
transform 1 0 22080 0 1 13600
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_21_236
timestamp 1586364061
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_240
timestamp 1586364061
transform 1 0 23184 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_249
timestamp 1586364061
transform 1 0 24012 0 1 13600
box -38 -48 406 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 25116 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_259
timestamp 1586364061
transform 1 0 24932 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_263
timestamp 1586364061
transform 1 0 25300 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_275
timestamp 1586364061
transform 1 0 26404 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  FILLER_22_9
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_21
timestamp 1586364061
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_25
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_28
timestamp 1586364061
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 5060 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_41
timestamp 1586364061
transform 1 0 4876 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_45
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_55
timestamp 1586364061
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_59
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_22_64
timestamp 1586364061
transform 1 0 6992 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_82
timestamp 1586364061
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_119
timestamp 1586364061
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_or3_4  _102_
timestamp 1586364061
transform 1 0 12788 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_136
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 590 592
use scs8hd_or3_4  _089_
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_146
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_149
timestamp 1586364061
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__C
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_8  _192_
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_179
timestamp 1586364061
transform 1 0 17572 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_186
timestamp 1586364061
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_196
timestamp 1586364061
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21896 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_218
timestamp 1586364061
transform 1 0 21160 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_229
timestamp 1586364061
transform 1 0 22172 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_right_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_241
timestamp 1586364061
transform 1 0 23276 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_247
timestamp 1586364061
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_258
timestamp 1586364061
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_270
timestamp 1586364061
transform 1 0 25944 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_274
timestamp 1586364061
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _155_
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 866 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_35
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 5060 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_58
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_66
timestamp 1586364061
transform 1 0 7176 0 1 14688
box -38 -48 130 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_78
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_82
timestamp 1586364061
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_95
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_99
timestamp 1586364061
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _098_
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_112
timestamp 1586364061
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_inv_8  _088_
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_136
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_or3_4  _127_
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_149
timestamp 1586364061
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_166
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_23_173
timestamp 1586364061
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20792 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_217
timestamp 1586364061
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23828 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_249
timestamp 1586364061
transform 1 0 24012 0 1 14688
box -38 -48 590 592
use scs8hd_buf_2  _230_
timestamp 1586364061
transform 1 0 24564 0 1 14688
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_259
timestamp 1586364061
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_263
timestamp 1586364061
transform 1 0 25300 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_275
timestamp 1586364061
transform 1 0 26404 0 1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__221__A
timestamp 1586364061
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_16
timestamp 1586364061
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_35
timestamp 1586364061
transform 1 0 4324 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_46
timestamp 1586364061
transform 1 0 5336 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_50
timestamp 1586364061
transform 1 0 5704 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_65
timestamp 1586364061
transform 1 0 7084 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_71
timestamp 1586364061
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 7820 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_82
timestamp 1586364061
transform 1 0 8648 0 -1 15776
box -38 -48 590 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 10580 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_90
timestamp 1586364061
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 590 592
use scs8hd_or3_4  _095_
timestamp 1586364061
transform 1 0 12144 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_112
timestamp 1586364061
transform 1 0 11408 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13708 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_140
timestamp 1586364061
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use scs8hd_or3_4  _137_
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_24_150
timestamp 1586364061
transform 1 0 14904 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_8  _135_
timestamp 1586364061
transform 1 0 16836 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__127__C
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_167
timestamp 1586364061
transform 1 0 16468 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 18400 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_180
timestamp 1586364061
transform 1 0 17664 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 19412 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 21896 0 -1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_218
timestamp 1586364061
transform 1 0 21160 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_12  FILLER_24_229
timestamp 1586364061
transform 1 0 22172 0 -1 15776
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23644 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_4  FILLER_24_241
timestamp 1586364061
transform 1 0 23276 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_248
timestamp 1586364061
transform 1 0 23920 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_259
timestamp 1586364061
transform 1 0 24932 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_271
timestamp 1586364061
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_11
timestamp 1586364061
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_18
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_22
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_33
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _154_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_40
timestamp 1586364061
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_66
timestamp 1586364061
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 9200 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_84
timestamp 1586364061
transform 1 0 8832 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_97
timestamp 1586364061
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_136
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_inv_8  _136_
timestamp 1586364061
transform 1 0 15272 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _169_
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_163
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_167
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_buf_1  _161_
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_203
timestamp 1586364061
transform 1 0 19780 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 21068 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_215
timestamp 1586364061
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_conb_1  _206_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_236
timestamp 1586364061
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_248
timestamp 1586364061
transform 1 0 23920 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_252
timestamp 1586364061
transform 1 0 24288 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_259
timestamp 1586364061
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_263
timestamp 1586364061
transform 1 0 25300 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_275
timestamp 1586364061
transform 1 0 26404 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_6
timestamp 1586364061
transform 1 0 1656 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_7
timestamp 1586364061
transform 1 0 1748 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use scs8hd_buf_2  _221_
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_17
timestamp 1586364061
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_21
timestamp 1586364061
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3220 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_32
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_30
timestamp 1586364061
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_35
timestamp 1586364061
transform 1 0 4324 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_18
timestamp 1586364061
transform 1 0 2760 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_50
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_52
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_47
timestamp 1586364061
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 314 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 5612 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_58
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_54
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6624 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_69
timestamp 1586364061
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_65
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_63
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 7636 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_107
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 406 592
use scs8hd_decap_8  FILLER_27_97
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 774 592
use scs8hd_decap_4  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_108
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use scs8hd_inv_8  _083_
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_132
timestamp 1586364061
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_131
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_136
timestamp 1586364061
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13524 0 -1 16864
box -38 -48 866 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 866 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_152
timestamp 1586364061
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_buf_1  _162_
timestamp 1586364061
transform 1 0 16836 0 -1 16864
box -38 -48 314 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_26_174
timestamp 1586364061
transform 1 0 17112 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_164
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_27_168
timestamp 1586364061
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_180
timestamp 1586364061
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_218
timestamp 1586364061
transform 1 0 21160 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_230
timestamp 1586364061
transform 1 0 22264 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 23736 0 1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_right_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23552 0 -1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_26_242
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_247
timestamp 1586364061
transform 1 0 23828 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_27_249
timestamp 1586364061
transform 1 0 24012 0 1 16864
box -38 -48 590 592
use scs8hd_inv_1  mux_right_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_258
timestamp 1586364061
transform 1 0 24840 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_270
timestamp 1586364061
transform 1 0 25944 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_274
timestamp 1586364061
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_7
timestamp 1586364061
transform 1 0 1748 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_46
timestamp 1586364061
transform 1 0 5336 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_58
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_64
timestamp 1586364061
transform 1 0 6992 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_76
timestamp 1586364061
transform 1 0 8096 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _205_
timestamp 1586364061
transform 1 0 12328 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_8  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_142
timestamp 1586364061
transform 1 0 14168 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_28_150
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_160
timestamp 1586364061
transform 1 0 15824 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_172
timestamp 1586364061
transform 1 0 16928 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_28_208
timestamp 1586364061
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_259
timestamp 1586364061
transform 1 0 24932 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_271
timestamp 1586364061
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_14
timestamp 1586364061
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 2760 0 1 17952
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3772 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_21
timestamp 1586364061
transform 1 0 3036 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_48
timestamp 1586364061
transform 1 0 5520 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_60
timestamp 1586364061
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_65
timestamp 1586364061
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_69
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_93
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_105
timestamp 1586364061
transform 1 0 10764 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 -1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_30_6
timestamp 1586364061
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use scs8hd_decap_12  FILLER_30_17
timestamp 1586364061
transform 1 0 2668 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_30_29
timestamp 1586364061
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2392 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_6
timestamp 1586364061
transform 1 0 1656 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_10
timestamp 1586364061
transform 1 0 2024 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_17
timestamp 1586364061
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_21
timestamp 1586364061
transform 1 0 3036 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_33
timestamp 1586364061
transform 1 0 4140 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_45
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_31_57
timestamp 1586364061
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_6
timestamp 1586364061
transform 1 0 1656 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_18
timestamp 1586364061
transform 1 0 2760 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_30
timestamp 1586364061
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_6
timestamp 1586364061
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_10
timestamp 1586364061
transform 1 0 2024 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_22
timestamp 1586364061
transform 1 0 3128 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_34
timestamp 1586364061
transform 1 0 4232 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_46
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_3  FILLER_33_58
timestamp 1586364061
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 1932 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_7
timestamp 1586364061
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_11
timestamp 1586364061
transform 1 0 2116 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_23
timestamp 1586364061
transform 1 0 3220 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_35
timestamp 1586364061
transform 1 0 4324 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_47
timestamp 1586364061
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 24564 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 25116 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_253
timestamp 1586364061
transform 1 0 24380 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_259
timestamp 1586364061
transform 1 0 24932 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_263
timestamp 1586364061
transform 1 0 25300 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_275
timestamp 1586364061
transform 1 0 26404 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _220_
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__220__A
timestamp 1586364061
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_7
timestamp 1586364061
transform 1 0 1748 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_11
timestamp 1586364061
transform 1 0 2116 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_23
timestamp 1586364061
transform 1 0 3220 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_35
timestamp 1586364061
transform 1 0 4324 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_47
timestamp 1586364061
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 11978 0 12034 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 12990 0 13046 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 13910 0 13966 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 14922 0 14978 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 15842 0 15898 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 16854 0 16910 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 17774 0 17830 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 10046 0 10102 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal3 s 0 24216 480 24336 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal3 s 0 25304 480 25424 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 26256 480 26376 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal3 s 0 27344 480 27464 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 27520 9664 28000 9784 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 27520 21088 28000 21208 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal3 s 27520 24216 28000 24336 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal3 s 27520 25304 28000 25424 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 27520 26256 28000 26376 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal3 s 27520 27344 28000 27464 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[0]
port 45 nsew default input
rlabel metal2 s 2318 0 2374 480 6 chany_bottom_in[1]
port 46 nsew default input
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_in[2]
port 47 nsew default input
rlabel metal2 s 4250 0 4306 480 6 chany_bottom_in[3]
port 48 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[4]
port 49 nsew default input
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[5]
port 50 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[6]
port 51 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[7]
port 52 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[8]
port 53 nsew default input
rlabel metal2 s 19706 0 19762 480 6 chany_bottom_out[0]
port 54 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[1]
port 55 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[2]
port 56 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[3]
port 57 nsew default tristate
rlabel metal2 s 23570 0 23626 480 6 chany_bottom_out[4]
port 58 nsew default tristate
rlabel metal2 s 24582 0 24638 480 6 chany_bottom_out[5]
port 59 nsew default tristate
rlabel metal2 s 25502 0 25558 480 6 chany_bottom_out[6]
port 60 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[7]
port 61 nsew default tristate
rlabel metal2 s 27434 0 27490 480 6 chany_bottom_out[8]
port 62 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 data_in
port 63 nsew default input
rlabel metal2 s 11058 0 11114 480 6 enable
port 64 nsew default input
rlabel metal3 s 0 17960 480 18080 6 left_bottom_grid_pin_12_
port 65 nsew default input
rlabel metal3 s 0 5584 480 5704 6 left_top_grid_pin_11_
port 66 nsew default input
rlabel metal3 s 0 6536 480 6656 6 left_top_grid_pin_13_
port 67 nsew default input
rlabel metal3 s 0 7624 480 7744 6 left_top_grid_pin_15_
port 68 nsew default input
rlabel metal3 s 0 416 480 536 6 left_top_grid_pin_1_
port 69 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_top_grid_pin_3_
port 70 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_top_grid_pin_5_
port 71 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_top_grid_pin_7_
port 72 nsew default input
rlabel metal3 s 0 4496 480 4616 6 left_top_grid_pin_9_
port 73 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 right_bottom_grid_pin_12_
port 74 nsew default input
rlabel metal3 s 27520 5584 28000 5704 6 right_top_grid_pin_11_
port 75 nsew default input
rlabel metal3 s 27520 6536 28000 6656 6 right_top_grid_pin_13_
port 76 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 right_top_grid_pin_15_
port 77 nsew default input
rlabel metal3 s 27520 416 28000 536 6 right_top_grid_pin_1_
port 78 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_top_grid_pin_3_
port 79 nsew default input
rlabel metal3 s 27520 2456 28000 2576 6 right_top_grid_pin_5_
port 80 nsew default input
rlabel metal3 s 27520 3408 28000 3528 6 right_top_grid_pin_7_
port 81 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 right_top_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< end >>
