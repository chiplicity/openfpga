magic
tech sky130A
magscale 1 2
timestamp 1609105282
<< viali >>
rect 8387 4165 8421 4199
rect 2131 4029 2165 4063
rect 2131 3349 2165 3383
rect 3511 3349 3545 3383
rect 4523 3349 4557 3383
rect 5995 3349 6029 3383
rect 7467 3349 7501 3383
rect 8387 2941 8421 2975
<< metal1 >>
rect 354 11450 10106 11472
rect 354 11398 3496 11450
rect 3548 11398 3560 11450
rect 3612 11398 3624 11450
rect 3676 11398 3688 11450
rect 3740 11398 6760 11450
rect 6812 11398 6824 11450
rect 6876 11398 6888 11450
rect 6940 11398 6952 11450
rect 7004 11398 10106 11450
rect 354 11376 10106 11398
rect 354 10906 10106 10928
rect 354 10854 1864 10906
rect 1916 10854 1928 10906
rect 1980 10854 1992 10906
rect 2044 10854 2056 10906
rect 2108 10854 5128 10906
rect 5180 10854 5192 10906
rect 5244 10854 5256 10906
rect 5308 10854 5320 10906
rect 5372 10854 8392 10906
rect 8444 10854 8456 10906
rect 8508 10854 8520 10906
rect 8572 10854 8584 10906
rect 8636 10854 10106 10906
rect 354 10832 10106 10854
rect 354 10362 10106 10384
rect 354 10310 3496 10362
rect 3548 10310 3560 10362
rect 3612 10310 3624 10362
rect 3676 10310 3688 10362
rect 3740 10310 6760 10362
rect 6812 10310 6824 10362
rect 6876 10310 6888 10362
rect 6940 10310 6952 10362
rect 7004 10310 10106 10362
rect 354 10288 10106 10310
rect 354 9818 10106 9840
rect 354 9766 1864 9818
rect 1916 9766 1928 9818
rect 1980 9766 1992 9818
rect 2044 9766 2056 9818
rect 2108 9766 5128 9818
rect 5180 9766 5192 9818
rect 5244 9766 5256 9818
rect 5308 9766 5320 9818
rect 5372 9766 8392 9818
rect 8444 9766 8456 9818
rect 8508 9766 8520 9818
rect 8572 9766 8584 9818
rect 8636 9766 10106 9818
rect 354 9744 10106 9766
rect 354 9274 10106 9296
rect 354 9222 3496 9274
rect 3548 9222 3560 9274
rect 3612 9222 3624 9274
rect 3676 9222 3688 9274
rect 3740 9222 6760 9274
rect 6812 9222 6824 9274
rect 6876 9222 6888 9274
rect 6940 9222 6952 9274
rect 7004 9222 10106 9274
rect 354 9200 10106 9222
rect 354 8730 10106 8752
rect 354 8678 1864 8730
rect 1916 8678 1928 8730
rect 1980 8678 1992 8730
rect 2044 8678 2056 8730
rect 2108 8678 5128 8730
rect 5180 8678 5192 8730
rect 5244 8678 5256 8730
rect 5308 8678 5320 8730
rect 5372 8678 8392 8730
rect 8444 8678 8456 8730
rect 8508 8678 8520 8730
rect 8572 8678 8584 8730
rect 8636 8678 10106 8730
rect 354 8656 10106 8678
rect 354 8186 10106 8208
rect 354 8134 3496 8186
rect 3548 8134 3560 8186
rect 3612 8134 3624 8186
rect 3676 8134 3688 8186
rect 3740 8134 6760 8186
rect 6812 8134 6824 8186
rect 6876 8134 6888 8186
rect 6940 8134 6952 8186
rect 7004 8134 10106 8186
rect 354 8112 10106 8134
rect 354 7642 10106 7664
rect 354 7590 1864 7642
rect 1916 7590 1928 7642
rect 1980 7590 1992 7642
rect 2044 7590 2056 7642
rect 2108 7590 5128 7642
rect 5180 7590 5192 7642
rect 5244 7590 5256 7642
rect 5308 7590 5320 7642
rect 5372 7590 8392 7642
rect 8444 7590 8456 7642
rect 8508 7590 8520 7642
rect 8572 7590 8584 7642
rect 8636 7590 10106 7642
rect 354 7568 10106 7590
rect 354 7098 10106 7120
rect 354 7046 3496 7098
rect 3548 7046 3560 7098
rect 3612 7046 3624 7098
rect 3676 7046 3688 7098
rect 3740 7046 6760 7098
rect 6812 7046 6824 7098
rect 6876 7046 6888 7098
rect 6940 7046 6952 7098
rect 7004 7046 10106 7098
rect 354 7024 10106 7046
rect 354 6554 10106 6576
rect 354 6502 1864 6554
rect 1916 6502 1928 6554
rect 1980 6502 1992 6554
rect 2044 6502 2056 6554
rect 2108 6502 5128 6554
rect 5180 6502 5192 6554
rect 5244 6502 5256 6554
rect 5308 6502 5320 6554
rect 5372 6502 8392 6554
rect 8444 6502 8456 6554
rect 8508 6502 8520 6554
rect 8572 6502 8584 6554
rect 8636 6502 10106 6554
rect 354 6480 10106 6502
rect 354 6010 10106 6032
rect 354 5958 3496 6010
rect 3548 5958 3560 6010
rect 3612 5958 3624 6010
rect 3676 5958 3688 6010
rect 3740 5958 6760 6010
rect 6812 5958 6824 6010
rect 6876 5958 6888 6010
rect 6940 5958 6952 6010
rect 7004 5958 10106 6010
rect 354 5936 10106 5958
rect 354 5466 10106 5488
rect 354 5414 1864 5466
rect 1916 5414 1928 5466
rect 1980 5414 1992 5466
rect 2044 5414 2056 5466
rect 2108 5414 5128 5466
rect 5180 5414 5192 5466
rect 5244 5414 5256 5466
rect 5308 5414 5320 5466
rect 5372 5414 8392 5466
rect 8444 5414 8456 5466
rect 8508 5414 8520 5466
rect 8572 5414 8584 5466
rect 8636 5414 10106 5466
rect 354 5392 10106 5414
rect 354 4922 10106 4944
rect 354 4870 3496 4922
rect 3548 4870 3560 4922
rect 3612 4870 3624 4922
rect 3676 4870 3688 4922
rect 3740 4870 6760 4922
rect 6812 4870 6824 4922
rect 6876 4870 6888 4922
rect 6940 4870 6952 4922
rect 7004 4870 10106 4922
rect 354 4848 10106 4870
rect 354 4378 10106 4400
rect 354 4326 1864 4378
rect 1916 4326 1928 4378
rect 1980 4326 1992 4378
rect 2044 4326 2056 4378
rect 2108 4326 5128 4378
rect 5180 4326 5192 4378
rect 5244 4326 5256 4378
rect 5308 4326 5320 4378
rect 5372 4326 8392 4378
rect 8444 4326 8456 4378
rect 8508 4326 8520 4378
rect 8572 4326 8584 4378
rect 8636 4326 10106 4378
rect 354 4304 10106 4326
rect 8375 4199 8433 4205
rect 8375 4165 8387 4199
rect 8421 4196 8433 4199
rect 8924 4196 8930 4208
rect 8421 4168 8930 4196
rect 8421 4165 8433 4168
rect 8375 4159 8433 4165
rect 8924 4156 8930 4168
rect 8982 4156 8988 4208
rect 1472 4020 1478 4072
rect 1530 4060 1536 4072
rect 2119 4063 2177 4069
rect 2119 4060 2131 4063
rect 1530 4032 2131 4060
rect 1530 4020 1536 4032
rect 2119 4029 2131 4032
rect 2165 4029 2177 4063
rect 2119 4023 2177 4029
rect 354 3834 10106 3856
rect 354 3782 3496 3834
rect 3548 3782 3560 3834
rect 3612 3782 3624 3834
rect 3676 3782 3688 3834
rect 3740 3782 6760 3834
rect 6812 3782 6824 3834
rect 6876 3782 6888 3834
rect 6940 3782 6952 3834
rect 7004 3782 10106 3834
rect 354 3760 10106 3782
rect 0 3340 6 3392
rect 58 3380 64 3392
rect 2119 3383 2177 3389
rect 2119 3380 2131 3383
rect 58 3352 2131 3380
rect 58 3340 64 3352
rect 2119 3349 2131 3352
rect 2165 3349 2177 3383
rect 2119 3343 2177 3349
rect 2944 3340 2950 3392
rect 3002 3380 3008 3392
rect 3499 3383 3557 3389
rect 3499 3380 3511 3383
rect 3002 3352 3511 3380
rect 3002 3340 3008 3352
rect 3499 3349 3511 3352
rect 3545 3349 3557 3383
rect 3499 3343 3557 3349
rect 4416 3340 4422 3392
rect 4474 3380 4480 3392
rect 4511 3383 4569 3389
rect 4511 3380 4523 3383
rect 4474 3352 4523 3380
rect 4474 3340 4480 3352
rect 4511 3349 4523 3352
rect 4557 3349 4569 3383
rect 5980 3380 5986 3392
rect 5941 3352 5986 3380
rect 4511 3343 4569 3349
rect 5980 3340 5986 3352
rect 6038 3340 6044 3392
rect 7452 3380 7458 3392
rect 7413 3352 7458 3380
rect 7452 3340 7458 3352
rect 7510 3340 7516 3392
rect 354 3290 10106 3312
rect 354 3238 1864 3290
rect 1916 3238 1928 3290
rect 1980 3238 1992 3290
rect 2044 3238 2056 3290
rect 2108 3238 5128 3290
rect 5180 3238 5192 3290
rect 5244 3238 5256 3290
rect 5308 3238 5320 3290
rect 5372 3238 8392 3290
rect 8444 3238 8456 3290
rect 8508 3238 8520 3290
rect 8572 3238 8584 3290
rect 8636 3238 10106 3290
rect 354 3216 10106 3238
rect 8375 2975 8433 2981
rect 8375 2941 8387 2975
rect 8421 2972 8433 2975
rect 10396 2972 10402 2984
rect 8421 2944 10402 2972
rect 8421 2941 8433 2944
rect 8375 2935 8433 2941
rect 10396 2932 10402 2944
rect 10454 2932 10460 2984
rect 354 2746 10106 2768
rect 354 2694 3496 2746
rect 3548 2694 3560 2746
rect 3612 2694 3624 2746
rect 3676 2694 3688 2746
rect 3740 2694 6760 2746
rect 6812 2694 6824 2746
rect 6876 2694 6888 2746
rect 6940 2694 6952 2746
rect 7004 2694 10106 2746
rect 354 2672 10106 2694
rect 354 2202 10106 2224
rect 354 2150 1864 2202
rect 1916 2150 1928 2202
rect 1980 2150 1992 2202
rect 2044 2150 2056 2202
rect 2108 2150 5128 2202
rect 5180 2150 5192 2202
rect 5244 2150 5256 2202
rect 5308 2150 5320 2202
rect 5372 2150 8392 2202
rect 8444 2150 8456 2202
rect 8508 2150 8520 2202
rect 8572 2150 8584 2202
rect 8636 2150 10106 2202
rect 354 2128 10106 2150
<< via1 >>
rect 3496 11398 3548 11450
rect 3560 11398 3612 11450
rect 3624 11398 3676 11450
rect 3688 11398 3740 11450
rect 6760 11398 6812 11450
rect 6824 11398 6876 11450
rect 6888 11398 6940 11450
rect 6952 11398 7004 11450
rect 1864 10854 1916 10906
rect 1928 10854 1980 10906
rect 1992 10854 2044 10906
rect 2056 10854 2108 10906
rect 5128 10854 5180 10906
rect 5192 10854 5244 10906
rect 5256 10854 5308 10906
rect 5320 10854 5372 10906
rect 8392 10854 8444 10906
rect 8456 10854 8508 10906
rect 8520 10854 8572 10906
rect 8584 10854 8636 10906
rect 3496 10310 3548 10362
rect 3560 10310 3612 10362
rect 3624 10310 3676 10362
rect 3688 10310 3740 10362
rect 6760 10310 6812 10362
rect 6824 10310 6876 10362
rect 6888 10310 6940 10362
rect 6952 10310 7004 10362
rect 1864 9766 1916 9818
rect 1928 9766 1980 9818
rect 1992 9766 2044 9818
rect 2056 9766 2108 9818
rect 5128 9766 5180 9818
rect 5192 9766 5244 9818
rect 5256 9766 5308 9818
rect 5320 9766 5372 9818
rect 8392 9766 8444 9818
rect 8456 9766 8508 9818
rect 8520 9766 8572 9818
rect 8584 9766 8636 9818
rect 3496 9222 3548 9274
rect 3560 9222 3612 9274
rect 3624 9222 3676 9274
rect 3688 9222 3740 9274
rect 6760 9222 6812 9274
rect 6824 9222 6876 9274
rect 6888 9222 6940 9274
rect 6952 9222 7004 9274
rect 1864 8678 1916 8730
rect 1928 8678 1980 8730
rect 1992 8678 2044 8730
rect 2056 8678 2108 8730
rect 5128 8678 5180 8730
rect 5192 8678 5244 8730
rect 5256 8678 5308 8730
rect 5320 8678 5372 8730
rect 8392 8678 8444 8730
rect 8456 8678 8508 8730
rect 8520 8678 8572 8730
rect 8584 8678 8636 8730
rect 3496 8134 3548 8186
rect 3560 8134 3612 8186
rect 3624 8134 3676 8186
rect 3688 8134 3740 8186
rect 6760 8134 6812 8186
rect 6824 8134 6876 8186
rect 6888 8134 6940 8186
rect 6952 8134 7004 8186
rect 1864 7590 1916 7642
rect 1928 7590 1980 7642
rect 1992 7590 2044 7642
rect 2056 7590 2108 7642
rect 5128 7590 5180 7642
rect 5192 7590 5244 7642
rect 5256 7590 5308 7642
rect 5320 7590 5372 7642
rect 8392 7590 8444 7642
rect 8456 7590 8508 7642
rect 8520 7590 8572 7642
rect 8584 7590 8636 7642
rect 3496 7046 3548 7098
rect 3560 7046 3612 7098
rect 3624 7046 3676 7098
rect 3688 7046 3740 7098
rect 6760 7046 6812 7098
rect 6824 7046 6876 7098
rect 6888 7046 6940 7098
rect 6952 7046 7004 7098
rect 1864 6502 1916 6554
rect 1928 6502 1980 6554
rect 1992 6502 2044 6554
rect 2056 6502 2108 6554
rect 5128 6502 5180 6554
rect 5192 6502 5244 6554
rect 5256 6502 5308 6554
rect 5320 6502 5372 6554
rect 8392 6502 8444 6554
rect 8456 6502 8508 6554
rect 8520 6502 8572 6554
rect 8584 6502 8636 6554
rect 3496 5958 3548 6010
rect 3560 5958 3612 6010
rect 3624 5958 3676 6010
rect 3688 5958 3740 6010
rect 6760 5958 6812 6010
rect 6824 5958 6876 6010
rect 6888 5958 6940 6010
rect 6952 5958 7004 6010
rect 1864 5414 1916 5466
rect 1928 5414 1980 5466
rect 1992 5414 2044 5466
rect 2056 5414 2108 5466
rect 5128 5414 5180 5466
rect 5192 5414 5244 5466
rect 5256 5414 5308 5466
rect 5320 5414 5372 5466
rect 8392 5414 8444 5466
rect 8456 5414 8508 5466
rect 8520 5414 8572 5466
rect 8584 5414 8636 5466
rect 3496 4870 3548 4922
rect 3560 4870 3612 4922
rect 3624 4870 3676 4922
rect 3688 4870 3740 4922
rect 6760 4870 6812 4922
rect 6824 4870 6876 4922
rect 6888 4870 6940 4922
rect 6952 4870 7004 4922
rect 1864 4326 1916 4378
rect 1928 4326 1980 4378
rect 1992 4326 2044 4378
rect 2056 4326 2108 4378
rect 5128 4326 5180 4378
rect 5192 4326 5244 4378
rect 5256 4326 5308 4378
rect 5320 4326 5372 4378
rect 8392 4326 8444 4378
rect 8456 4326 8508 4378
rect 8520 4326 8572 4378
rect 8584 4326 8636 4378
rect 8930 4156 8982 4208
rect 1478 4020 1530 4072
rect 3496 3782 3548 3834
rect 3560 3782 3612 3834
rect 3624 3782 3676 3834
rect 3688 3782 3740 3834
rect 6760 3782 6812 3834
rect 6824 3782 6876 3834
rect 6888 3782 6940 3834
rect 6952 3782 7004 3834
rect 6 3340 58 3392
rect 2950 3340 3002 3392
rect 4422 3340 4474 3392
rect 5986 3383 6038 3392
rect 5986 3349 5995 3383
rect 5995 3349 6029 3383
rect 6029 3349 6038 3383
rect 5986 3340 6038 3349
rect 7458 3383 7510 3392
rect 7458 3349 7467 3383
rect 7467 3349 7501 3383
rect 7501 3349 7510 3383
rect 7458 3340 7510 3349
rect 1864 3238 1916 3290
rect 1928 3238 1980 3290
rect 1992 3238 2044 3290
rect 2056 3238 2108 3290
rect 5128 3238 5180 3290
rect 5192 3238 5244 3290
rect 5256 3238 5308 3290
rect 5320 3238 5372 3290
rect 8392 3238 8444 3290
rect 8456 3238 8508 3290
rect 8520 3238 8572 3290
rect 8584 3238 8636 3290
rect 10402 2932 10454 2984
rect 3496 2694 3548 2746
rect 3560 2694 3612 2746
rect 3624 2694 3676 2746
rect 3688 2694 3740 2746
rect 6760 2694 6812 2746
rect 6824 2694 6876 2746
rect 6888 2694 6940 2746
rect 6952 2694 7004 2746
rect 1864 2150 1916 2202
rect 1928 2150 1980 2202
rect 1992 2150 2044 2202
rect 2056 2150 2108 2202
rect 5128 2150 5180 2202
rect 5192 2150 5244 2202
rect 5256 2150 5308 2202
rect 5320 2150 5372 2202
rect 8392 2150 8444 2202
rect 8456 2150 8508 2202
rect 8520 2150 8572 2202
rect 8584 2150 8636 2202
<< metal2 >>
rect 3470 11452 3766 11472
rect 3526 11450 3550 11452
rect 3606 11450 3630 11452
rect 3686 11450 3710 11452
rect 3548 11398 3550 11450
rect 3612 11398 3624 11450
rect 3686 11398 3688 11450
rect 3526 11396 3550 11398
rect 3606 11396 3630 11398
rect 3686 11396 3710 11398
rect 3470 11376 3766 11396
rect 6734 11452 7030 11472
rect 6790 11450 6814 11452
rect 6870 11450 6894 11452
rect 6950 11450 6974 11452
rect 6812 11398 6814 11450
rect 6876 11398 6888 11450
rect 6950 11398 6952 11450
rect 6790 11396 6814 11398
rect 6870 11396 6894 11398
rect 6950 11396 6974 11398
rect 6734 11376 7030 11396
rect 1838 10908 2134 10928
rect 1894 10906 1918 10908
rect 1974 10906 1998 10908
rect 2054 10906 2078 10908
rect 1916 10854 1918 10906
rect 1980 10854 1992 10906
rect 2054 10854 2056 10906
rect 1894 10852 1918 10854
rect 1974 10852 1998 10854
rect 2054 10852 2078 10854
rect 1838 10832 2134 10852
rect 5102 10908 5398 10928
rect 5158 10906 5182 10908
rect 5238 10906 5262 10908
rect 5318 10906 5342 10908
rect 5180 10854 5182 10906
rect 5244 10854 5256 10906
rect 5318 10854 5320 10906
rect 5158 10852 5182 10854
rect 5238 10852 5262 10854
rect 5318 10852 5342 10854
rect 5102 10832 5398 10852
rect 8366 10908 8662 10928
rect 8422 10906 8446 10908
rect 8502 10906 8526 10908
rect 8582 10906 8606 10908
rect 8444 10854 8446 10906
rect 8508 10854 8520 10906
rect 8582 10854 8584 10906
rect 8422 10852 8446 10854
rect 8502 10852 8526 10854
rect 8582 10852 8606 10854
rect 8366 10832 8662 10852
rect 3470 10364 3766 10384
rect 3526 10362 3550 10364
rect 3606 10362 3630 10364
rect 3686 10362 3710 10364
rect 3548 10310 3550 10362
rect 3612 10310 3624 10362
rect 3686 10310 3688 10362
rect 3526 10308 3550 10310
rect 3606 10308 3630 10310
rect 3686 10308 3710 10310
rect 3470 10288 3766 10308
rect 6734 10364 7030 10384
rect 6790 10362 6814 10364
rect 6870 10362 6894 10364
rect 6950 10362 6974 10364
rect 6812 10310 6814 10362
rect 6876 10310 6888 10362
rect 6950 10310 6952 10362
rect 6790 10308 6814 10310
rect 6870 10308 6894 10310
rect 6950 10308 6974 10310
rect 6734 10288 7030 10308
rect 1838 9820 2134 9840
rect 1894 9818 1918 9820
rect 1974 9818 1998 9820
rect 2054 9818 2078 9820
rect 1916 9766 1918 9818
rect 1980 9766 1992 9818
rect 2054 9766 2056 9818
rect 1894 9764 1918 9766
rect 1974 9764 1998 9766
rect 2054 9764 2078 9766
rect 1838 9744 2134 9764
rect 5102 9820 5398 9840
rect 5158 9818 5182 9820
rect 5238 9818 5262 9820
rect 5318 9818 5342 9820
rect 5180 9766 5182 9818
rect 5244 9766 5256 9818
rect 5318 9766 5320 9818
rect 5158 9764 5182 9766
rect 5238 9764 5262 9766
rect 5318 9764 5342 9766
rect 5102 9744 5398 9764
rect 8366 9820 8662 9840
rect 8422 9818 8446 9820
rect 8502 9818 8526 9820
rect 8582 9818 8606 9820
rect 8444 9766 8446 9818
rect 8508 9766 8520 9818
rect 8582 9766 8584 9818
rect 8422 9764 8446 9766
rect 8502 9764 8526 9766
rect 8582 9764 8606 9766
rect 8366 9744 8662 9764
rect 3470 9276 3766 9296
rect 3526 9274 3550 9276
rect 3606 9274 3630 9276
rect 3686 9274 3710 9276
rect 3548 9222 3550 9274
rect 3612 9222 3624 9274
rect 3686 9222 3688 9274
rect 3526 9220 3550 9222
rect 3606 9220 3630 9222
rect 3686 9220 3710 9222
rect 3470 9200 3766 9220
rect 6734 9276 7030 9296
rect 6790 9274 6814 9276
rect 6870 9274 6894 9276
rect 6950 9274 6974 9276
rect 6812 9222 6814 9274
rect 6876 9222 6888 9274
rect 6950 9222 6952 9274
rect 6790 9220 6814 9222
rect 6870 9220 6894 9222
rect 6950 9220 6974 9222
rect 6734 9200 7030 9220
rect 1838 8732 2134 8752
rect 1894 8730 1918 8732
rect 1974 8730 1998 8732
rect 2054 8730 2078 8732
rect 1916 8678 1918 8730
rect 1980 8678 1992 8730
rect 2054 8678 2056 8730
rect 1894 8676 1918 8678
rect 1974 8676 1998 8678
rect 2054 8676 2078 8678
rect 1838 8656 2134 8676
rect 5102 8732 5398 8752
rect 5158 8730 5182 8732
rect 5238 8730 5262 8732
rect 5318 8730 5342 8732
rect 5180 8678 5182 8730
rect 5244 8678 5256 8730
rect 5318 8678 5320 8730
rect 5158 8676 5182 8678
rect 5238 8676 5262 8678
rect 5318 8676 5342 8678
rect 5102 8656 5398 8676
rect 8366 8732 8662 8752
rect 8422 8730 8446 8732
rect 8502 8730 8526 8732
rect 8582 8730 8606 8732
rect 8444 8678 8446 8730
rect 8508 8678 8520 8730
rect 8582 8678 8584 8730
rect 8422 8676 8446 8678
rect 8502 8676 8526 8678
rect 8582 8676 8606 8678
rect 8366 8656 8662 8676
rect 3470 8188 3766 8208
rect 3526 8186 3550 8188
rect 3606 8186 3630 8188
rect 3686 8186 3710 8188
rect 3548 8134 3550 8186
rect 3612 8134 3624 8186
rect 3686 8134 3688 8186
rect 3526 8132 3550 8134
rect 3606 8132 3630 8134
rect 3686 8132 3710 8134
rect 3470 8112 3766 8132
rect 6734 8188 7030 8208
rect 6790 8186 6814 8188
rect 6870 8186 6894 8188
rect 6950 8186 6974 8188
rect 6812 8134 6814 8186
rect 6876 8134 6888 8186
rect 6950 8134 6952 8186
rect 6790 8132 6814 8134
rect 6870 8132 6894 8134
rect 6950 8132 6974 8134
rect 6734 8112 7030 8132
rect 1838 7644 2134 7664
rect 1894 7642 1918 7644
rect 1974 7642 1998 7644
rect 2054 7642 2078 7644
rect 1916 7590 1918 7642
rect 1980 7590 1992 7642
rect 2054 7590 2056 7642
rect 1894 7588 1918 7590
rect 1974 7588 1998 7590
rect 2054 7588 2078 7590
rect 1838 7568 2134 7588
rect 5102 7644 5398 7664
rect 5158 7642 5182 7644
rect 5238 7642 5262 7644
rect 5318 7642 5342 7644
rect 5180 7590 5182 7642
rect 5244 7590 5256 7642
rect 5318 7590 5320 7642
rect 5158 7588 5182 7590
rect 5238 7588 5262 7590
rect 5318 7588 5342 7590
rect 5102 7568 5398 7588
rect 8366 7644 8662 7664
rect 8422 7642 8446 7644
rect 8502 7642 8526 7644
rect 8582 7642 8606 7644
rect 8444 7590 8446 7642
rect 8508 7590 8520 7642
rect 8582 7590 8584 7642
rect 8422 7588 8446 7590
rect 8502 7588 8526 7590
rect 8582 7588 8606 7590
rect 8366 7568 8662 7588
rect 3470 7100 3766 7120
rect 3526 7098 3550 7100
rect 3606 7098 3630 7100
rect 3686 7098 3710 7100
rect 3548 7046 3550 7098
rect 3612 7046 3624 7098
rect 3686 7046 3688 7098
rect 3526 7044 3550 7046
rect 3606 7044 3630 7046
rect 3686 7044 3710 7046
rect 3470 7024 3766 7044
rect 6734 7100 7030 7120
rect 6790 7098 6814 7100
rect 6870 7098 6894 7100
rect 6950 7098 6974 7100
rect 6812 7046 6814 7098
rect 6876 7046 6888 7098
rect 6950 7046 6952 7098
rect 6790 7044 6814 7046
rect 6870 7044 6894 7046
rect 6950 7044 6974 7046
rect 6734 7024 7030 7044
rect 1838 6556 2134 6576
rect 1894 6554 1918 6556
rect 1974 6554 1998 6556
rect 2054 6554 2078 6556
rect 1916 6502 1918 6554
rect 1980 6502 1992 6554
rect 2054 6502 2056 6554
rect 1894 6500 1918 6502
rect 1974 6500 1998 6502
rect 2054 6500 2078 6502
rect 1838 6480 2134 6500
rect 5102 6556 5398 6576
rect 5158 6554 5182 6556
rect 5238 6554 5262 6556
rect 5318 6554 5342 6556
rect 5180 6502 5182 6554
rect 5244 6502 5256 6554
rect 5318 6502 5320 6554
rect 5158 6500 5182 6502
rect 5238 6500 5262 6502
rect 5318 6500 5342 6502
rect 5102 6480 5398 6500
rect 8366 6556 8662 6576
rect 8422 6554 8446 6556
rect 8502 6554 8526 6556
rect 8582 6554 8606 6556
rect 8444 6502 8446 6554
rect 8508 6502 8520 6554
rect 8582 6502 8584 6554
rect 8422 6500 8446 6502
rect 8502 6500 8526 6502
rect 8582 6500 8606 6502
rect 8366 6480 8662 6500
rect 3470 6012 3766 6032
rect 3526 6010 3550 6012
rect 3606 6010 3630 6012
rect 3686 6010 3710 6012
rect 3548 5958 3550 6010
rect 3612 5958 3624 6010
rect 3686 5958 3688 6010
rect 3526 5956 3550 5958
rect 3606 5956 3630 5958
rect 3686 5956 3710 5958
rect 3470 5936 3766 5956
rect 6734 6012 7030 6032
rect 6790 6010 6814 6012
rect 6870 6010 6894 6012
rect 6950 6010 6974 6012
rect 6812 5958 6814 6010
rect 6876 5958 6888 6010
rect 6950 5958 6952 6010
rect 6790 5956 6814 5958
rect 6870 5956 6894 5958
rect 6950 5956 6974 5958
rect 6734 5936 7030 5956
rect 1838 5468 2134 5488
rect 1894 5466 1918 5468
rect 1974 5466 1998 5468
rect 2054 5466 2078 5468
rect 1916 5414 1918 5466
rect 1980 5414 1992 5466
rect 2054 5414 2056 5466
rect 1894 5412 1918 5414
rect 1974 5412 1998 5414
rect 2054 5412 2078 5414
rect 1838 5392 2134 5412
rect 5102 5468 5398 5488
rect 5158 5466 5182 5468
rect 5238 5466 5262 5468
rect 5318 5466 5342 5468
rect 5180 5414 5182 5466
rect 5244 5414 5256 5466
rect 5318 5414 5320 5466
rect 5158 5412 5182 5414
rect 5238 5412 5262 5414
rect 5318 5412 5342 5414
rect 5102 5392 5398 5412
rect 8366 5468 8662 5488
rect 8422 5466 8446 5468
rect 8502 5466 8526 5468
rect 8582 5466 8606 5468
rect 8444 5414 8446 5466
rect 8508 5414 8520 5466
rect 8582 5414 8584 5466
rect 8422 5412 8446 5414
rect 8502 5412 8526 5414
rect 8582 5412 8606 5414
rect 8366 5392 8662 5412
rect 3470 4924 3766 4944
rect 3526 4922 3550 4924
rect 3606 4922 3630 4924
rect 3686 4922 3710 4924
rect 3548 4870 3550 4922
rect 3612 4870 3624 4922
rect 3686 4870 3688 4922
rect 3526 4868 3550 4870
rect 3606 4868 3630 4870
rect 3686 4868 3710 4870
rect 3470 4848 3766 4868
rect 6734 4924 7030 4944
rect 6790 4922 6814 4924
rect 6870 4922 6894 4924
rect 6950 4922 6974 4924
rect 6812 4870 6814 4922
rect 6876 4870 6888 4922
rect 6950 4870 6952 4922
rect 6790 4868 6814 4870
rect 6870 4868 6894 4870
rect 6950 4868 6974 4870
rect 6734 4848 7030 4868
rect 1838 4380 2134 4400
rect 1894 4378 1918 4380
rect 1974 4378 1998 4380
rect 2054 4378 2078 4380
rect 1916 4326 1918 4378
rect 1980 4326 1992 4378
rect 2054 4326 2056 4378
rect 1894 4324 1918 4326
rect 1974 4324 1998 4326
rect 2054 4324 2078 4326
rect 1838 4304 2134 4324
rect 5102 4380 5398 4400
rect 5158 4378 5182 4380
rect 5238 4378 5262 4380
rect 5318 4378 5342 4380
rect 5180 4326 5182 4378
rect 5244 4326 5256 4378
rect 5318 4326 5320 4378
rect 5158 4324 5182 4326
rect 5238 4324 5262 4326
rect 5318 4324 5342 4326
rect 5102 4304 5398 4324
rect 8366 4380 8662 4400
rect 8422 4378 8446 4380
rect 8502 4378 8526 4380
rect 8582 4378 8606 4380
rect 8444 4326 8446 4378
rect 8508 4326 8520 4378
rect 8582 4326 8584 4378
rect 8422 4324 8446 4326
rect 8502 4324 8526 4326
rect 8582 4324 8606 4326
rect 8366 4304 8662 4324
rect 8930 4208 8982 4214
rect 8930 4150 8982 4156
rect 1478 4072 1530 4078
rect 1478 4014 1530 4020
rect 6 3392 58 3398
rect 6 3334 58 3340
rect 18 800 46 3334
rect 1490 800 1518 4014
rect 3470 3836 3766 3856
rect 3526 3834 3550 3836
rect 3606 3834 3630 3836
rect 3686 3834 3710 3836
rect 3548 3782 3550 3834
rect 3612 3782 3624 3834
rect 3686 3782 3688 3834
rect 3526 3780 3550 3782
rect 3606 3780 3630 3782
rect 3686 3780 3710 3782
rect 3470 3760 3766 3780
rect 6734 3836 7030 3856
rect 6790 3834 6814 3836
rect 6870 3834 6894 3836
rect 6950 3834 6974 3836
rect 6812 3782 6814 3834
rect 6876 3782 6888 3834
rect 6950 3782 6952 3834
rect 6790 3780 6814 3782
rect 6870 3780 6894 3782
rect 6950 3780 6974 3782
rect 6734 3760 7030 3780
rect 2950 3392 3002 3398
rect 2950 3334 3002 3340
rect 4422 3392 4474 3398
rect 4422 3334 4474 3340
rect 5986 3392 6038 3398
rect 5986 3334 6038 3340
rect 7458 3392 7510 3398
rect 7458 3334 7510 3340
rect 1838 3292 2134 3312
rect 1894 3290 1918 3292
rect 1974 3290 1998 3292
rect 2054 3290 2078 3292
rect 1916 3238 1918 3290
rect 1980 3238 1992 3290
rect 2054 3238 2056 3290
rect 1894 3236 1918 3238
rect 1974 3236 1998 3238
rect 2054 3236 2078 3238
rect 1838 3216 2134 3236
rect 1838 2204 2134 2224
rect 1894 2202 1918 2204
rect 1974 2202 1998 2204
rect 2054 2202 2078 2204
rect 1916 2150 1918 2202
rect 1980 2150 1992 2202
rect 2054 2150 2056 2202
rect 1894 2148 1918 2150
rect 1974 2148 1998 2150
rect 2054 2148 2078 2150
rect 1838 2128 2134 2148
rect 2962 800 2990 3334
rect 3470 2748 3766 2768
rect 3526 2746 3550 2748
rect 3606 2746 3630 2748
rect 3686 2746 3710 2748
rect 3548 2694 3550 2746
rect 3612 2694 3624 2746
rect 3686 2694 3688 2746
rect 3526 2692 3550 2694
rect 3606 2692 3630 2694
rect 3686 2692 3710 2694
rect 3470 2672 3766 2692
rect 4434 800 4462 3334
rect 5102 3292 5398 3312
rect 5158 3290 5182 3292
rect 5238 3290 5262 3292
rect 5318 3290 5342 3292
rect 5180 3238 5182 3290
rect 5244 3238 5256 3290
rect 5318 3238 5320 3290
rect 5158 3236 5182 3238
rect 5238 3236 5262 3238
rect 5318 3236 5342 3238
rect 5102 3216 5398 3236
rect 5102 2204 5398 2224
rect 5158 2202 5182 2204
rect 5238 2202 5262 2204
rect 5318 2202 5342 2204
rect 5180 2150 5182 2202
rect 5244 2150 5256 2202
rect 5318 2150 5320 2202
rect 5158 2148 5182 2150
rect 5238 2148 5262 2150
rect 5318 2148 5342 2150
rect 5102 2128 5398 2148
rect 5998 800 6026 3334
rect 6734 2748 7030 2768
rect 6790 2746 6814 2748
rect 6870 2746 6894 2748
rect 6950 2746 6974 2748
rect 6812 2694 6814 2746
rect 6876 2694 6888 2746
rect 6950 2694 6952 2746
rect 6790 2692 6814 2694
rect 6870 2692 6894 2694
rect 6950 2692 6974 2694
rect 6734 2672 7030 2692
rect 7470 800 7498 3334
rect 8366 3292 8662 3312
rect 8422 3290 8446 3292
rect 8502 3290 8526 3292
rect 8582 3290 8606 3292
rect 8444 3238 8446 3290
rect 8508 3238 8520 3290
rect 8582 3238 8584 3290
rect 8422 3236 8446 3238
rect 8502 3236 8526 3238
rect 8582 3236 8606 3238
rect 8366 3216 8662 3236
rect 8366 2204 8662 2224
rect 8422 2202 8446 2204
rect 8502 2202 8526 2204
rect 8582 2202 8606 2204
rect 8444 2150 8446 2202
rect 8508 2150 8520 2202
rect 8582 2150 8584 2202
rect 8422 2148 8446 2150
rect 8502 2148 8526 2150
rect 8582 2148 8606 2150
rect 8366 2128 8662 2148
rect 8942 800 8970 4150
rect 10402 2984 10454 2990
rect 10402 2926 10454 2932
rect 10414 800 10442 2926
rect 4 0 60 800
rect 1476 0 1532 800
rect 2948 0 3004 800
rect 4420 0 4476 800
rect 5984 0 6040 800
rect 7456 0 7512 800
rect 8928 0 8984 800
rect 10400 0 10456 800
<< via2 >>
rect 3470 11450 3526 11452
rect 3550 11450 3606 11452
rect 3630 11450 3686 11452
rect 3710 11450 3766 11452
rect 3470 11398 3496 11450
rect 3496 11398 3526 11450
rect 3550 11398 3560 11450
rect 3560 11398 3606 11450
rect 3630 11398 3676 11450
rect 3676 11398 3686 11450
rect 3710 11398 3740 11450
rect 3740 11398 3766 11450
rect 3470 11396 3526 11398
rect 3550 11396 3606 11398
rect 3630 11396 3686 11398
rect 3710 11396 3766 11398
rect 6734 11450 6790 11452
rect 6814 11450 6870 11452
rect 6894 11450 6950 11452
rect 6974 11450 7030 11452
rect 6734 11398 6760 11450
rect 6760 11398 6790 11450
rect 6814 11398 6824 11450
rect 6824 11398 6870 11450
rect 6894 11398 6940 11450
rect 6940 11398 6950 11450
rect 6974 11398 7004 11450
rect 7004 11398 7030 11450
rect 6734 11396 6790 11398
rect 6814 11396 6870 11398
rect 6894 11396 6950 11398
rect 6974 11396 7030 11398
rect 1838 10906 1894 10908
rect 1918 10906 1974 10908
rect 1998 10906 2054 10908
rect 2078 10906 2134 10908
rect 1838 10854 1864 10906
rect 1864 10854 1894 10906
rect 1918 10854 1928 10906
rect 1928 10854 1974 10906
rect 1998 10854 2044 10906
rect 2044 10854 2054 10906
rect 2078 10854 2108 10906
rect 2108 10854 2134 10906
rect 1838 10852 1894 10854
rect 1918 10852 1974 10854
rect 1998 10852 2054 10854
rect 2078 10852 2134 10854
rect 5102 10906 5158 10908
rect 5182 10906 5238 10908
rect 5262 10906 5318 10908
rect 5342 10906 5398 10908
rect 5102 10854 5128 10906
rect 5128 10854 5158 10906
rect 5182 10854 5192 10906
rect 5192 10854 5238 10906
rect 5262 10854 5308 10906
rect 5308 10854 5318 10906
rect 5342 10854 5372 10906
rect 5372 10854 5398 10906
rect 5102 10852 5158 10854
rect 5182 10852 5238 10854
rect 5262 10852 5318 10854
rect 5342 10852 5398 10854
rect 8366 10906 8422 10908
rect 8446 10906 8502 10908
rect 8526 10906 8582 10908
rect 8606 10906 8662 10908
rect 8366 10854 8392 10906
rect 8392 10854 8422 10906
rect 8446 10854 8456 10906
rect 8456 10854 8502 10906
rect 8526 10854 8572 10906
rect 8572 10854 8582 10906
rect 8606 10854 8636 10906
rect 8636 10854 8662 10906
rect 8366 10852 8422 10854
rect 8446 10852 8502 10854
rect 8526 10852 8582 10854
rect 8606 10852 8662 10854
rect 3470 10362 3526 10364
rect 3550 10362 3606 10364
rect 3630 10362 3686 10364
rect 3710 10362 3766 10364
rect 3470 10310 3496 10362
rect 3496 10310 3526 10362
rect 3550 10310 3560 10362
rect 3560 10310 3606 10362
rect 3630 10310 3676 10362
rect 3676 10310 3686 10362
rect 3710 10310 3740 10362
rect 3740 10310 3766 10362
rect 3470 10308 3526 10310
rect 3550 10308 3606 10310
rect 3630 10308 3686 10310
rect 3710 10308 3766 10310
rect 6734 10362 6790 10364
rect 6814 10362 6870 10364
rect 6894 10362 6950 10364
rect 6974 10362 7030 10364
rect 6734 10310 6760 10362
rect 6760 10310 6790 10362
rect 6814 10310 6824 10362
rect 6824 10310 6870 10362
rect 6894 10310 6940 10362
rect 6940 10310 6950 10362
rect 6974 10310 7004 10362
rect 7004 10310 7030 10362
rect 6734 10308 6790 10310
rect 6814 10308 6870 10310
rect 6894 10308 6950 10310
rect 6974 10308 7030 10310
rect 1838 9818 1894 9820
rect 1918 9818 1974 9820
rect 1998 9818 2054 9820
rect 2078 9818 2134 9820
rect 1838 9766 1864 9818
rect 1864 9766 1894 9818
rect 1918 9766 1928 9818
rect 1928 9766 1974 9818
rect 1998 9766 2044 9818
rect 2044 9766 2054 9818
rect 2078 9766 2108 9818
rect 2108 9766 2134 9818
rect 1838 9764 1894 9766
rect 1918 9764 1974 9766
rect 1998 9764 2054 9766
rect 2078 9764 2134 9766
rect 5102 9818 5158 9820
rect 5182 9818 5238 9820
rect 5262 9818 5318 9820
rect 5342 9818 5398 9820
rect 5102 9766 5128 9818
rect 5128 9766 5158 9818
rect 5182 9766 5192 9818
rect 5192 9766 5238 9818
rect 5262 9766 5308 9818
rect 5308 9766 5318 9818
rect 5342 9766 5372 9818
rect 5372 9766 5398 9818
rect 5102 9764 5158 9766
rect 5182 9764 5238 9766
rect 5262 9764 5318 9766
rect 5342 9764 5398 9766
rect 8366 9818 8422 9820
rect 8446 9818 8502 9820
rect 8526 9818 8582 9820
rect 8606 9818 8662 9820
rect 8366 9766 8392 9818
rect 8392 9766 8422 9818
rect 8446 9766 8456 9818
rect 8456 9766 8502 9818
rect 8526 9766 8572 9818
rect 8572 9766 8582 9818
rect 8606 9766 8636 9818
rect 8636 9766 8662 9818
rect 8366 9764 8422 9766
rect 8446 9764 8502 9766
rect 8526 9764 8582 9766
rect 8606 9764 8662 9766
rect 3470 9274 3526 9276
rect 3550 9274 3606 9276
rect 3630 9274 3686 9276
rect 3710 9274 3766 9276
rect 3470 9222 3496 9274
rect 3496 9222 3526 9274
rect 3550 9222 3560 9274
rect 3560 9222 3606 9274
rect 3630 9222 3676 9274
rect 3676 9222 3686 9274
rect 3710 9222 3740 9274
rect 3740 9222 3766 9274
rect 3470 9220 3526 9222
rect 3550 9220 3606 9222
rect 3630 9220 3686 9222
rect 3710 9220 3766 9222
rect 6734 9274 6790 9276
rect 6814 9274 6870 9276
rect 6894 9274 6950 9276
rect 6974 9274 7030 9276
rect 6734 9222 6760 9274
rect 6760 9222 6790 9274
rect 6814 9222 6824 9274
rect 6824 9222 6870 9274
rect 6894 9222 6940 9274
rect 6940 9222 6950 9274
rect 6974 9222 7004 9274
rect 7004 9222 7030 9274
rect 6734 9220 6790 9222
rect 6814 9220 6870 9222
rect 6894 9220 6950 9222
rect 6974 9220 7030 9222
rect 1838 8730 1894 8732
rect 1918 8730 1974 8732
rect 1998 8730 2054 8732
rect 2078 8730 2134 8732
rect 1838 8678 1864 8730
rect 1864 8678 1894 8730
rect 1918 8678 1928 8730
rect 1928 8678 1974 8730
rect 1998 8678 2044 8730
rect 2044 8678 2054 8730
rect 2078 8678 2108 8730
rect 2108 8678 2134 8730
rect 1838 8676 1894 8678
rect 1918 8676 1974 8678
rect 1998 8676 2054 8678
rect 2078 8676 2134 8678
rect 5102 8730 5158 8732
rect 5182 8730 5238 8732
rect 5262 8730 5318 8732
rect 5342 8730 5398 8732
rect 5102 8678 5128 8730
rect 5128 8678 5158 8730
rect 5182 8678 5192 8730
rect 5192 8678 5238 8730
rect 5262 8678 5308 8730
rect 5308 8678 5318 8730
rect 5342 8678 5372 8730
rect 5372 8678 5398 8730
rect 5102 8676 5158 8678
rect 5182 8676 5238 8678
rect 5262 8676 5318 8678
rect 5342 8676 5398 8678
rect 8366 8730 8422 8732
rect 8446 8730 8502 8732
rect 8526 8730 8582 8732
rect 8606 8730 8662 8732
rect 8366 8678 8392 8730
rect 8392 8678 8422 8730
rect 8446 8678 8456 8730
rect 8456 8678 8502 8730
rect 8526 8678 8572 8730
rect 8572 8678 8582 8730
rect 8606 8678 8636 8730
rect 8636 8678 8662 8730
rect 8366 8676 8422 8678
rect 8446 8676 8502 8678
rect 8526 8676 8582 8678
rect 8606 8676 8662 8678
rect 3470 8186 3526 8188
rect 3550 8186 3606 8188
rect 3630 8186 3686 8188
rect 3710 8186 3766 8188
rect 3470 8134 3496 8186
rect 3496 8134 3526 8186
rect 3550 8134 3560 8186
rect 3560 8134 3606 8186
rect 3630 8134 3676 8186
rect 3676 8134 3686 8186
rect 3710 8134 3740 8186
rect 3740 8134 3766 8186
rect 3470 8132 3526 8134
rect 3550 8132 3606 8134
rect 3630 8132 3686 8134
rect 3710 8132 3766 8134
rect 6734 8186 6790 8188
rect 6814 8186 6870 8188
rect 6894 8186 6950 8188
rect 6974 8186 7030 8188
rect 6734 8134 6760 8186
rect 6760 8134 6790 8186
rect 6814 8134 6824 8186
rect 6824 8134 6870 8186
rect 6894 8134 6940 8186
rect 6940 8134 6950 8186
rect 6974 8134 7004 8186
rect 7004 8134 7030 8186
rect 6734 8132 6790 8134
rect 6814 8132 6870 8134
rect 6894 8132 6950 8134
rect 6974 8132 7030 8134
rect 1838 7642 1894 7644
rect 1918 7642 1974 7644
rect 1998 7642 2054 7644
rect 2078 7642 2134 7644
rect 1838 7590 1864 7642
rect 1864 7590 1894 7642
rect 1918 7590 1928 7642
rect 1928 7590 1974 7642
rect 1998 7590 2044 7642
rect 2044 7590 2054 7642
rect 2078 7590 2108 7642
rect 2108 7590 2134 7642
rect 1838 7588 1894 7590
rect 1918 7588 1974 7590
rect 1998 7588 2054 7590
rect 2078 7588 2134 7590
rect 5102 7642 5158 7644
rect 5182 7642 5238 7644
rect 5262 7642 5318 7644
rect 5342 7642 5398 7644
rect 5102 7590 5128 7642
rect 5128 7590 5158 7642
rect 5182 7590 5192 7642
rect 5192 7590 5238 7642
rect 5262 7590 5308 7642
rect 5308 7590 5318 7642
rect 5342 7590 5372 7642
rect 5372 7590 5398 7642
rect 5102 7588 5158 7590
rect 5182 7588 5238 7590
rect 5262 7588 5318 7590
rect 5342 7588 5398 7590
rect 8366 7642 8422 7644
rect 8446 7642 8502 7644
rect 8526 7642 8582 7644
rect 8606 7642 8662 7644
rect 8366 7590 8392 7642
rect 8392 7590 8422 7642
rect 8446 7590 8456 7642
rect 8456 7590 8502 7642
rect 8526 7590 8572 7642
rect 8572 7590 8582 7642
rect 8606 7590 8636 7642
rect 8636 7590 8662 7642
rect 8366 7588 8422 7590
rect 8446 7588 8502 7590
rect 8526 7588 8582 7590
rect 8606 7588 8662 7590
rect 3470 7098 3526 7100
rect 3550 7098 3606 7100
rect 3630 7098 3686 7100
rect 3710 7098 3766 7100
rect 3470 7046 3496 7098
rect 3496 7046 3526 7098
rect 3550 7046 3560 7098
rect 3560 7046 3606 7098
rect 3630 7046 3676 7098
rect 3676 7046 3686 7098
rect 3710 7046 3740 7098
rect 3740 7046 3766 7098
rect 3470 7044 3526 7046
rect 3550 7044 3606 7046
rect 3630 7044 3686 7046
rect 3710 7044 3766 7046
rect 6734 7098 6790 7100
rect 6814 7098 6870 7100
rect 6894 7098 6950 7100
rect 6974 7098 7030 7100
rect 6734 7046 6760 7098
rect 6760 7046 6790 7098
rect 6814 7046 6824 7098
rect 6824 7046 6870 7098
rect 6894 7046 6940 7098
rect 6940 7046 6950 7098
rect 6974 7046 7004 7098
rect 7004 7046 7030 7098
rect 6734 7044 6790 7046
rect 6814 7044 6870 7046
rect 6894 7044 6950 7046
rect 6974 7044 7030 7046
rect 1838 6554 1894 6556
rect 1918 6554 1974 6556
rect 1998 6554 2054 6556
rect 2078 6554 2134 6556
rect 1838 6502 1864 6554
rect 1864 6502 1894 6554
rect 1918 6502 1928 6554
rect 1928 6502 1974 6554
rect 1998 6502 2044 6554
rect 2044 6502 2054 6554
rect 2078 6502 2108 6554
rect 2108 6502 2134 6554
rect 1838 6500 1894 6502
rect 1918 6500 1974 6502
rect 1998 6500 2054 6502
rect 2078 6500 2134 6502
rect 5102 6554 5158 6556
rect 5182 6554 5238 6556
rect 5262 6554 5318 6556
rect 5342 6554 5398 6556
rect 5102 6502 5128 6554
rect 5128 6502 5158 6554
rect 5182 6502 5192 6554
rect 5192 6502 5238 6554
rect 5262 6502 5308 6554
rect 5308 6502 5318 6554
rect 5342 6502 5372 6554
rect 5372 6502 5398 6554
rect 5102 6500 5158 6502
rect 5182 6500 5238 6502
rect 5262 6500 5318 6502
rect 5342 6500 5398 6502
rect 8366 6554 8422 6556
rect 8446 6554 8502 6556
rect 8526 6554 8582 6556
rect 8606 6554 8662 6556
rect 8366 6502 8392 6554
rect 8392 6502 8422 6554
rect 8446 6502 8456 6554
rect 8456 6502 8502 6554
rect 8526 6502 8572 6554
rect 8572 6502 8582 6554
rect 8606 6502 8636 6554
rect 8636 6502 8662 6554
rect 8366 6500 8422 6502
rect 8446 6500 8502 6502
rect 8526 6500 8582 6502
rect 8606 6500 8662 6502
rect 3470 6010 3526 6012
rect 3550 6010 3606 6012
rect 3630 6010 3686 6012
rect 3710 6010 3766 6012
rect 3470 5958 3496 6010
rect 3496 5958 3526 6010
rect 3550 5958 3560 6010
rect 3560 5958 3606 6010
rect 3630 5958 3676 6010
rect 3676 5958 3686 6010
rect 3710 5958 3740 6010
rect 3740 5958 3766 6010
rect 3470 5956 3526 5958
rect 3550 5956 3606 5958
rect 3630 5956 3686 5958
rect 3710 5956 3766 5958
rect 6734 6010 6790 6012
rect 6814 6010 6870 6012
rect 6894 6010 6950 6012
rect 6974 6010 7030 6012
rect 6734 5958 6760 6010
rect 6760 5958 6790 6010
rect 6814 5958 6824 6010
rect 6824 5958 6870 6010
rect 6894 5958 6940 6010
rect 6940 5958 6950 6010
rect 6974 5958 7004 6010
rect 7004 5958 7030 6010
rect 6734 5956 6790 5958
rect 6814 5956 6870 5958
rect 6894 5956 6950 5958
rect 6974 5956 7030 5958
rect 1838 5466 1894 5468
rect 1918 5466 1974 5468
rect 1998 5466 2054 5468
rect 2078 5466 2134 5468
rect 1838 5414 1864 5466
rect 1864 5414 1894 5466
rect 1918 5414 1928 5466
rect 1928 5414 1974 5466
rect 1998 5414 2044 5466
rect 2044 5414 2054 5466
rect 2078 5414 2108 5466
rect 2108 5414 2134 5466
rect 1838 5412 1894 5414
rect 1918 5412 1974 5414
rect 1998 5412 2054 5414
rect 2078 5412 2134 5414
rect 5102 5466 5158 5468
rect 5182 5466 5238 5468
rect 5262 5466 5318 5468
rect 5342 5466 5398 5468
rect 5102 5414 5128 5466
rect 5128 5414 5158 5466
rect 5182 5414 5192 5466
rect 5192 5414 5238 5466
rect 5262 5414 5308 5466
rect 5308 5414 5318 5466
rect 5342 5414 5372 5466
rect 5372 5414 5398 5466
rect 5102 5412 5158 5414
rect 5182 5412 5238 5414
rect 5262 5412 5318 5414
rect 5342 5412 5398 5414
rect 8366 5466 8422 5468
rect 8446 5466 8502 5468
rect 8526 5466 8582 5468
rect 8606 5466 8662 5468
rect 8366 5414 8392 5466
rect 8392 5414 8422 5466
rect 8446 5414 8456 5466
rect 8456 5414 8502 5466
rect 8526 5414 8572 5466
rect 8572 5414 8582 5466
rect 8606 5414 8636 5466
rect 8636 5414 8662 5466
rect 8366 5412 8422 5414
rect 8446 5412 8502 5414
rect 8526 5412 8582 5414
rect 8606 5412 8662 5414
rect 3470 4922 3526 4924
rect 3550 4922 3606 4924
rect 3630 4922 3686 4924
rect 3710 4922 3766 4924
rect 3470 4870 3496 4922
rect 3496 4870 3526 4922
rect 3550 4870 3560 4922
rect 3560 4870 3606 4922
rect 3630 4870 3676 4922
rect 3676 4870 3686 4922
rect 3710 4870 3740 4922
rect 3740 4870 3766 4922
rect 3470 4868 3526 4870
rect 3550 4868 3606 4870
rect 3630 4868 3686 4870
rect 3710 4868 3766 4870
rect 6734 4922 6790 4924
rect 6814 4922 6870 4924
rect 6894 4922 6950 4924
rect 6974 4922 7030 4924
rect 6734 4870 6760 4922
rect 6760 4870 6790 4922
rect 6814 4870 6824 4922
rect 6824 4870 6870 4922
rect 6894 4870 6940 4922
rect 6940 4870 6950 4922
rect 6974 4870 7004 4922
rect 7004 4870 7030 4922
rect 6734 4868 6790 4870
rect 6814 4868 6870 4870
rect 6894 4868 6950 4870
rect 6974 4868 7030 4870
rect 1838 4378 1894 4380
rect 1918 4378 1974 4380
rect 1998 4378 2054 4380
rect 2078 4378 2134 4380
rect 1838 4326 1864 4378
rect 1864 4326 1894 4378
rect 1918 4326 1928 4378
rect 1928 4326 1974 4378
rect 1998 4326 2044 4378
rect 2044 4326 2054 4378
rect 2078 4326 2108 4378
rect 2108 4326 2134 4378
rect 1838 4324 1894 4326
rect 1918 4324 1974 4326
rect 1998 4324 2054 4326
rect 2078 4324 2134 4326
rect 5102 4378 5158 4380
rect 5182 4378 5238 4380
rect 5262 4378 5318 4380
rect 5342 4378 5398 4380
rect 5102 4326 5128 4378
rect 5128 4326 5158 4378
rect 5182 4326 5192 4378
rect 5192 4326 5238 4378
rect 5262 4326 5308 4378
rect 5308 4326 5318 4378
rect 5342 4326 5372 4378
rect 5372 4326 5398 4378
rect 5102 4324 5158 4326
rect 5182 4324 5238 4326
rect 5262 4324 5318 4326
rect 5342 4324 5398 4326
rect 8366 4378 8422 4380
rect 8446 4378 8502 4380
rect 8526 4378 8582 4380
rect 8606 4378 8662 4380
rect 8366 4326 8392 4378
rect 8392 4326 8422 4378
rect 8446 4326 8456 4378
rect 8456 4326 8502 4378
rect 8526 4326 8572 4378
rect 8572 4326 8582 4378
rect 8606 4326 8636 4378
rect 8636 4326 8662 4378
rect 8366 4324 8422 4326
rect 8446 4324 8502 4326
rect 8526 4324 8582 4326
rect 8606 4324 8662 4326
rect 3470 3834 3526 3836
rect 3550 3834 3606 3836
rect 3630 3834 3686 3836
rect 3710 3834 3766 3836
rect 3470 3782 3496 3834
rect 3496 3782 3526 3834
rect 3550 3782 3560 3834
rect 3560 3782 3606 3834
rect 3630 3782 3676 3834
rect 3676 3782 3686 3834
rect 3710 3782 3740 3834
rect 3740 3782 3766 3834
rect 3470 3780 3526 3782
rect 3550 3780 3606 3782
rect 3630 3780 3686 3782
rect 3710 3780 3766 3782
rect 6734 3834 6790 3836
rect 6814 3834 6870 3836
rect 6894 3834 6950 3836
rect 6974 3834 7030 3836
rect 6734 3782 6760 3834
rect 6760 3782 6790 3834
rect 6814 3782 6824 3834
rect 6824 3782 6870 3834
rect 6894 3782 6940 3834
rect 6940 3782 6950 3834
rect 6974 3782 7004 3834
rect 7004 3782 7030 3834
rect 6734 3780 6790 3782
rect 6814 3780 6870 3782
rect 6894 3780 6950 3782
rect 6974 3780 7030 3782
rect 1838 3290 1894 3292
rect 1918 3290 1974 3292
rect 1998 3290 2054 3292
rect 2078 3290 2134 3292
rect 1838 3238 1864 3290
rect 1864 3238 1894 3290
rect 1918 3238 1928 3290
rect 1928 3238 1974 3290
rect 1998 3238 2044 3290
rect 2044 3238 2054 3290
rect 2078 3238 2108 3290
rect 2108 3238 2134 3290
rect 1838 3236 1894 3238
rect 1918 3236 1974 3238
rect 1998 3236 2054 3238
rect 2078 3236 2134 3238
rect 1838 2202 1894 2204
rect 1918 2202 1974 2204
rect 1998 2202 2054 2204
rect 2078 2202 2134 2204
rect 1838 2150 1864 2202
rect 1864 2150 1894 2202
rect 1918 2150 1928 2202
rect 1928 2150 1974 2202
rect 1998 2150 2044 2202
rect 2044 2150 2054 2202
rect 2078 2150 2108 2202
rect 2108 2150 2134 2202
rect 1838 2148 1894 2150
rect 1918 2148 1974 2150
rect 1998 2148 2054 2150
rect 2078 2148 2134 2150
rect 3470 2746 3526 2748
rect 3550 2746 3606 2748
rect 3630 2746 3686 2748
rect 3710 2746 3766 2748
rect 3470 2694 3496 2746
rect 3496 2694 3526 2746
rect 3550 2694 3560 2746
rect 3560 2694 3606 2746
rect 3630 2694 3676 2746
rect 3676 2694 3686 2746
rect 3710 2694 3740 2746
rect 3740 2694 3766 2746
rect 3470 2692 3526 2694
rect 3550 2692 3606 2694
rect 3630 2692 3686 2694
rect 3710 2692 3766 2694
rect 5102 3290 5158 3292
rect 5182 3290 5238 3292
rect 5262 3290 5318 3292
rect 5342 3290 5398 3292
rect 5102 3238 5128 3290
rect 5128 3238 5158 3290
rect 5182 3238 5192 3290
rect 5192 3238 5238 3290
rect 5262 3238 5308 3290
rect 5308 3238 5318 3290
rect 5342 3238 5372 3290
rect 5372 3238 5398 3290
rect 5102 3236 5158 3238
rect 5182 3236 5238 3238
rect 5262 3236 5318 3238
rect 5342 3236 5398 3238
rect 5102 2202 5158 2204
rect 5182 2202 5238 2204
rect 5262 2202 5318 2204
rect 5342 2202 5398 2204
rect 5102 2150 5128 2202
rect 5128 2150 5158 2202
rect 5182 2150 5192 2202
rect 5192 2150 5238 2202
rect 5262 2150 5308 2202
rect 5308 2150 5318 2202
rect 5342 2150 5372 2202
rect 5372 2150 5398 2202
rect 5102 2148 5158 2150
rect 5182 2148 5238 2150
rect 5262 2148 5318 2150
rect 5342 2148 5398 2150
rect 6734 2746 6790 2748
rect 6814 2746 6870 2748
rect 6894 2746 6950 2748
rect 6974 2746 7030 2748
rect 6734 2694 6760 2746
rect 6760 2694 6790 2746
rect 6814 2694 6824 2746
rect 6824 2694 6870 2746
rect 6894 2694 6940 2746
rect 6940 2694 6950 2746
rect 6974 2694 7004 2746
rect 7004 2694 7030 2746
rect 6734 2692 6790 2694
rect 6814 2692 6870 2694
rect 6894 2692 6950 2694
rect 6974 2692 7030 2694
rect 8366 3290 8422 3292
rect 8446 3290 8502 3292
rect 8526 3290 8582 3292
rect 8606 3290 8662 3292
rect 8366 3238 8392 3290
rect 8392 3238 8422 3290
rect 8446 3238 8456 3290
rect 8456 3238 8502 3290
rect 8526 3238 8572 3290
rect 8572 3238 8582 3290
rect 8606 3238 8636 3290
rect 8636 3238 8662 3290
rect 8366 3236 8422 3238
rect 8446 3236 8502 3238
rect 8526 3236 8582 3238
rect 8606 3236 8662 3238
rect 8366 2202 8422 2204
rect 8446 2202 8502 2204
rect 8526 2202 8582 2204
rect 8606 2202 8662 2204
rect 8366 2150 8392 2202
rect 8392 2150 8422 2202
rect 8446 2150 8456 2202
rect 8456 2150 8502 2202
rect 8526 2150 8572 2202
rect 8572 2150 8582 2202
rect 8606 2150 8636 2202
rect 8636 2150 8662 2202
rect 8366 2148 8422 2150
rect 8446 2148 8502 2150
rect 8526 2148 8582 2150
rect 8606 2148 8662 2150
<< metal3 >>
rect 3458 11456 3778 11457
rect 3458 11392 3466 11456
rect 3530 11392 3546 11456
rect 3610 11392 3626 11456
rect 3690 11392 3706 11456
rect 3770 11392 3778 11456
rect 3458 11391 3778 11392
rect 6722 11456 7042 11457
rect 6722 11392 6730 11456
rect 6794 11392 6810 11456
rect 6874 11392 6890 11456
rect 6954 11392 6970 11456
rect 7034 11392 7042 11456
rect 6722 11391 7042 11392
rect 1826 10912 2146 10913
rect 1826 10848 1834 10912
rect 1898 10848 1914 10912
rect 1978 10848 1994 10912
rect 2058 10848 2074 10912
rect 2138 10848 2146 10912
rect 1826 10847 2146 10848
rect 5090 10912 5410 10913
rect 5090 10848 5098 10912
rect 5162 10848 5178 10912
rect 5242 10848 5258 10912
rect 5322 10848 5338 10912
rect 5402 10848 5410 10912
rect 5090 10847 5410 10848
rect 8354 10912 8674 10913
rect 8354 10848 8362 10912
rect 8426 10848 8442 10912
rect 8506 10848 8522 10912
rect 8586 10848 8602 10912
rect 8666 10848 8674 10912
rect 8354 10847 8674 10848
rect 3458 10368 3778 10369
rect 3458 10304 3466 10368
rect 3530 10304 3546 10368
rect 3610 10304 3626 10368
rect 3690 10304 3706 10368
rect 3770 10304 3778 10368
rect 3458 10303 3778 10304
rect 6722 10368 7042 10369
rect 6722 10304 6730 10368
rect 6794 10304 6810 10368
rect 6874 10304 6890 10368
rect 6954 10304 6970 10368
rect 7034 10304 7042 10368
rect 6722 10303 7042 10304
rect 1826 9824 2146 9825
rect 1826 9760 1834 9824
rect 1898 9760 1914 9824
rect 1978 9760 1994 9824
rect 2058 9760 2074 9824
rect 2138 9760 2146 9824
rect 1826 9759 2146 9760
rect 5090 9824 5410 9825
rect 5090 9760 5098 9824
rect 5162 9760 5178 9824
rect 5242 9760 5258 9824
rect 5322 9760 5338 9824
rect 5402 9760 5410 9824
rect 5090 9759 5410 9760
rect 8354 9824 8674 9825
rect 8354 9760 8362 9824
rect 8426 9760 8442 9824
rect 8506 9760 8522 9824
rect 8586 9760 8602 9824
rect 8666 9760 8674 9824
rect 8354 9759 8674 9760
rect 3458 9280 3778 9281
rect 3458 9216 3466 9280
rect 3530 9216 3546 9280
rect 3610 9216 3626 9280
rect 3690 9216 3706 9280
rect 3770 9216 3778 9280
rect 3458 9215 3778 9216
rect 6722 9280 7042 9281
rect 6722 9216 6730 9280
rect 6794 9216 6810 9280
rect 6874 9216 6890 9280
rect 6954 9216 6970 9280
rect 7034 9216 7042 9280
rect 6722 9215 7042 9216
rect 1826 8736 2146 8737
rect 1826 8672 1834 8736
rect 1898 8672 1914 8736
rect 1978 8672 1994 8736
rect 2058 8672 2074 8736
rect 2138 8672 2146 8736
rect 1826 8671 2146 8672
rect 5090 8736 5410 8737
rect 5090 8672 5098 8736
rect 5162 8672 5178 8736
rect 5242 8672 5258 8736
rect 5322 8672 5338 8736
rect 5402 8672 5410 8736
rect 5090 8671 5410 8672
rect 8354 8736 8674 8737
rect 8354 8672 8362 8736
rect 8426 8672 8442 8736
rect 8506 8672 8522 8736
rect 8586 8672 8602 8736
rect 8666 8672 8674 8736
rect 8354 8671 8674 8672
rect 3458 8192 3778 8193
rect 3458 8128 3466 8192
rect 3530 8128 3546 8192
rect 3610 8128 3626 8192
rect 3690 8128 3706 8192
rect 3770 8128 3778 8192
rect 3458 8127 3778 8128
rect 6722 8192 7042 8193
rect 6722 8128 6730 8192
rect 6794 8128 6810 8192
rect 6874 8128 6890 8192
rect 6954 8128 6970 8192
rect 7034 8128 7042 8192
rect 6722 8127 7042 8128
rect 1826 7648 2146 7649
rect 1826 7584 1834 7648
rect 1898 7584 1914 7648
rect 1978 7584 1994 7648
rect 2058 7584 2074 7648
rect 2138 7584 2146 7648
rect 1826 7583 2146 7584
rect 5090 7648 5410 7649
rect 5090 7584 5098 7648
rect 5162 7584 5178 7648
rect 5242 7584 5258 7648
rect 5322 7584 5338 7648
rect 5402 7584 5410 7648
rect 5090 7583 5410 7584
rect 8354 7648 8674 7649
rect 8354 7584 8362 7648
rect 8426 7584 8442 7648
rect 8506 7584 8522 7648
rect 8586 7584 8602 7648
rect 8666 7584 8674 7648
rect 8354 7583 8674 7584
rect 3458 7104 3778 7105
rect 3458 7040 3466 7104
rect 3530 7040 3546 7104
rect 3610 7040 3626 7104
rect 3690 7040 3706 7104
rect 3770 7040 3778 7104
rect 3458 7039 3778 7040
rect 6722 7104 7042 7105
rect 6722 7040 6730 7104
rect 6794 7040 6810 7104
rect 6874 7040 6890 7104
rect 6954 7040 6970 7104
rect 7034 7040 7042 7104
rect 6722 7039 7042 7040
rect 1826 6560 2146 6561
rect 1826 6496 1834 6560
rect 1898 6496 1914 6560
rect 1978 6496 1994 6560
rect 2058 6496 2074 6560
rect 2138 6496 2146 6560
rect 1826 6495 2146 6496
rect 5090 6560 5410 6561
rect 5090 6496 5098 6560
rect 5162 6496 5178 6560
rect 5242 6496 5258 6560
rect 5322 6496 5338 6560
rect 5402 6496 5410 6560
rect 5090 6495 5410 6496
rect 8354 6560 8674 6561
rect 8354 6496 8362 6560
rect 8426 6496 8442 6560
rect 8506 6496 8522 6560
rect 8586 6496 8602 6560
rect 8666 6496 8674 6560
rect 8354 6495 8674 6496
rect 3458 6016 3778 6017
rect 3458 5952 3466 6016
rect 3530 5952 3546 6016
rect 3610 5952 3626 6016
rect 3690 5952 3706 6016
rect 3770 5952 3778 6016
rect 3458 5951 3778 5952
rect 6722 6016 7042 6017
rect 6722 5952 6730 6016
rect 6794 5952 6810 6016
rect 6874 5952 6890 6016
rect 6954 5952 6970 6016
rect 7034 5952 7042 6016
rect 6722 5951 7042 5952
rect 1826 5472 2146 5473
rect 1826 5408 1834 5472
rect 1898 5408 1914 5472
rect 1978 5408 1994 5472
rect 2058 5408 2074 5472
rect 2138 5408 2146 5472
rect 1826 5407 2146 5408
rect 5090 5472 5410 5473
rect 5090 5408 5098 5472
rect 5162 5408 5178 5472
rect 5242 5408 5258 5472
rect 5322 5408 5338 5472
rect 5402 5408 5410 5472
rect 5090 5407 5410 5408
rect 8354 5472 8674 5473
rect 8354 5408 8362 5472
rect 8426 5408 8442 5472
rect 8506 5408 8522 5472
rect 8586 5408 8602 5472
rect 8666 5408 8674 5472
rect 8354 5407 8674 5408
rect 3458 4928 3778 4929
rect 3458 4864 3466 4928
rect 3530 4864 3546 4928
rect 3610 4864 3626 4928
rect 3690 4864 3706 4928
rect 3770 4864 3778 4928
rect 3458 4863 3778 4864
rect 6722 4928 7042 4929
rect 6722 4864 6730 4928
rect 6794 4864 6810 4928
rect 6874 4864 6890 4928
rect 6954 4864 6970 4928
rect 7034 4864 7042 4928
rect 6722 4863 7042 4864
rect 1826 4384 2146 4385
rect 1826 4320 1834 4384
rect 1898 4320 1914 4384
rect 1978 4320 1994 4384
rect 2058 4320 2074 4384
rect 2138 4320 2146 4384
rect 1826 4319 2146 4320
rect 5090 4384 5410 4385
rect 5090 4320 5098 4384
rect 5162 4320 5178 4384
rect 5242 4320 5258 4384
rect 5322 4320 5338 4384
rect 5402 4320 5410 4384
rect 5090 4319 5410 4320
rect 8354 4384 8674 4385
rect 8354 4320 8362 4384
rect 8426 4320 8442 4384
rect 8506 4320 8522 4384
rect 8586 4320 8602 4384
rect 8666 4320 8674 4384
rect 8354 4319 8674 4320
rect 3458 3840 3778 3841
rect 3458 3776 3466 3840
rect 3530 3776 3546 3840
rect 3610 3776 3626 3840
rect 3690 3776 3706 3840
rect 3770 3776 3778 3840
rect 3458 3775 3778 3776
rect 6722 3840 7042 3841
rect 6722 3776 6730 3840
rect 6794 3776 6810 3840
rect 6874 3776 6890 3840
rect 6954 3776 6970 3840
rect 7034 3776 7042 3840
rect 6722 3775 7042 3776
rect 1826 3296 2146 3297
rect 1826 3232 1834 3296
rect 1898 3232 1914 3296
rect 1978 3232 1994 3296
rect 2058 3232 2074 3296
rect 2138 3232 2146 3296
rect 1826 3231 2146 3232
rect 5090 3296 5410 3297
rect 5090 3232 5098 3296
rect 5162 3232 5178 3296
rect 5242 3232 5258 3296
rect 5322 3232 5338 3296
rect 5402 3232 5410 3296
rect 5090 3231 5410 3232
rect 8354 3296 8674 3297
rect 8354 3232 8362 3296
rect 8426 3232 8442 3296
rect 8506 3232 8522 3296
rect 8586 3232 8602 3296
rect 8666 3232 8674 3296
rect 8354 3231 8674 3232
rect 3458 2752 3778 2753
rect 3458 2688 3466 2752
rect 3530 2688 3546 2752
rect 3610 2688 3626 2752
rect 3690 2688 3706 2752
rect 3770 2688 3778 2752
rect 3458 2687 3778 2688
rect 6722 2752 7042 2753
rect 6722 2688 6730 2752
rect 6794 2688 6810 2752
rect 6874 2688 6890 2752
rect 6954 2688 6970 2752
rect 7034 2688 7042 2752
rect 6722 2687 7042 2688
rect 1826 2208 2146 2209
rect 1826 2144 1834 2208
rect 1898 2144 1914 2208
rect 1978 2144 1994 2208
rect 2058 2144 2074 2208
rect 2138 2144 2146 2208
rect 1826 2143 2146 2144
rect 5090 2208 5410 2209
rect 5090 2144 5098 2208
rect 5162 2144 5178 2208
rect 5242 2144 5258 2208
rect 5322 2144 5338 2208
rect 5402 2144 5410 2208
rect 5090 2143 5410 2144
rect 8354 2208 8674 2209
rect 8354 2144 8362 2208
rect 8426 2144 8442 2208
rect 8506 2144 8522 2208
rect 8586 2144 8602 2208
rect 8666 2144 8674 2208
rect 8354 2143 8674 2144
<< via3 >>
rect 3466 11452 3530 11456
rect 3466 11396 3470 11452
rect 3470 11396 3526 11452
rect 3526 11396 3530 11452
rect 3466 11392 3530 11396
rect 3546 11452 3610 11456
rect 3546 11396 3550 11452
rect 3550 11396 3606 11452
rect 3606 11396 3610 11452
rect 3546 11392 3610 11396
rect 3626 11452 3690 11456
rect 3626 11396 3630 11452
rect 3630 11396 3686 11452
rect 3686 11396 3690 11452
rect 3626 11392 3690 11396
rect 3706 11452 3770 11456
rect 3706 11396 3710 11452
rect 3710 11396 3766 11452
rect 3766 11396 3770 11452
rect 3706 11392 3770 11396
rect 6730 11452 6794 11456
rect 6730 11396 6734 11452
rect 6734 11396 6790 11452
rect 6790 11396 6794 11452
rect 6730 11392 6794 11396
rect 6810 11452 6874 11456
rect 6810 11396 6814 11452
rect 6814 11396 6870 11452
rect 6870 11396 6874 11452
rect 6810 11392 6874 11396
rect 6890 11452 6954 11456
rect 6890 11396 6894 11452
rect 6894 11396 6950 11452
rect 6950 11396 6954 11452
rect 6890 11392 6954 11396
rect 6970 11452 7034 11456
rect 6970 11396 6974 11452
rect 6974 11396 7030 11452
rect 7030 11396 7034 11452
rect 6970 11392 7034 11396
rect 1834 10908 1898 10912
rect 1834 10852 1838 10908
rect 1838 10852 1894 10908
rect 1894 10852 1898 10908
rect 1834 10848 1898 10852
rect 1914 10908 1978 10912
rect 1914 10852 1918 10908
rect 1918 10852 1974 10908
rect 1974 10852 1978 10908
rect 1914 10848 1978 10852
rect 1994 10908 2058 10912
rect 1994 10852 1998 10908
rect 1998 10852 2054 10908
rect 2054 10852 2058 10908
rect 1994 10848 2058 10852
rect 2074 10908 2138 10912
rect 2074 10852 2078 10908
rect 2078 10852 2134 10908
rect 2134 10852 2138 10908
rect 2074 10848 2138 10852
rect 5098 10908 5162 10912
rect 5098 10852 5102 10908
rect 5102 10852 5158 10908
rect 5158 10852 5162 10908
rect 5098 10848 5162 10852
rect 5178 10908 5242 10912
rect 5178 10852 5182 10908
rect 5182 10852 5238 10908
rect 5238 10852 5242 10908
rect 5178 10848 5242 10852
rect 5258 10908 5322 10912
rect 5258 10852 5262 10908
rect 5262 10852 5318 10908
rect 5318 10852 5322 10908
rect 5258 10848 5322 10852
rect 5338 10908 5402 10912
rect 5338 10852 5342 10908
rect 5342 10852 5398 10908
rect 5398 10852 5402 10908
rect 5338 10848 5402 10852
rect 8362 10908 8426 10912
rect 8362 10852 8366 10908
rect 8366 10852 8422 10908
rect 8422 10852 8426 10908
rect 8362 10848 8426 10852
rect 8442 10908 8506 10912
rect 8442 10852 8446 10908
rect 8446 10852 8502 10908
rect 8502 10852 8506 10908
rect 8442 10848 8506 10852
rect 8522 10908 8586 10912
rect 8522 10852 8526 10908
rect 8526 10852 8582 10908
rect 8582 10852 8586 10908
rect 8522 10848 8586 10852
rect 8602 10908 8666 10912
rect 8602 10852 8606 10908
rect 8606 10852 8662 10908
rect 8662 10852 8666 10908
rect 8602 10848 8666 10852
rect 3466 10364 3530 10368
rect 3466 10308 3470 10364
rect 3470 10308 3526 10364
rect 3526 10308 3530 10364
rect 3466 10304 3530 10308
rect 3546 10364 3610 10368
rect 3546 10308 3550 10364
rect 3550 10308 3606 10364
rect 3606 10308 3610 10364
rect 3546 10304 3610 10308
rect 3626 10364 3690 10368
rect 3626 10308 3630 10364
rect 3630 10308 3686 10364
rect 3686 10308 3690 10364
rect 3626 10304 3690 10308
rect 3706 10364 3770 10368
rect 3706 10308 3710 10364
rect 3710 10308 3766 10364
rect 3766 10308 3770 10364
rect 3706 10304 3770 10308
rect 6730 10364 6794 10368
rect 6730 10308 6734 10364
rect 6734 10308 6790 10364
rect 6790 10308 6794 10364
rect 6730 10304 6794 10308
rect 6810 10364 6874 10368
rect 6810 10308 6814 10364
rect 6814 10308 6870 10364
rect 6870 10308 6874 10364
rect 6810 10304 6874 10308
rect 6890 10364 6954 10368
rect 6890 10308 6894 10364
rect 6894 10308 6950 10364
rect 6950 10308 6954 10364
rect 6890 10304 6954 10308
rect 6970 10364 7034 10368
rect 6970 10308 6974 10364
rect 6974 10308 7030 10364
rect 7030 10308 7034 10364
rect 6970 10304 7034 10308
rect 1834 9820 1898 9824
rect 1834 9764 1838 9820
rect 1838 9764 1894 9820
rect 1894 9764 1898 9820
rect 1834 9760 1898 9764
rect 1914 9820 1978 9824
rect 1914 9764 1918 9820
rect 1918 9764 1974 9820
rect 1974 9764 1978 9820
rect 1914 9760 1978 9764
rect 1994 9820 2058 9824
rect 1994 9764 1998 9820
rect 1998 9764 2054 9820
rect 2054 9764 2058 9820
rect 1994 9760 2058 9764
rect 2074 9820 2138 9824
rect 2074 9764 2078 9820
rect 2078 9764 2134 9820
rect 2134 9764 2138 9820
rect 2074 9760 2138 9764
rect 5098 9820 5162 9824
rect 5098 9764 5102 9820
rect 5102 9764 5158 9820
rect 5158 9764 5162 9820
rect 5098 9760 5162 9764
rect 5178 9820 5242 9824
rect 5178 9764 5182 9820
rect 5182 9764 5238 9820
rect 5238 9764 5242 9820
rect 5178 9760 5242 9764
rect 5258 9820 5322 9824
rect 5258 9764 5262 9820
rect 5262 9764 5318 9820
rect 5318 9764 5322 9820
rect 5258 9760 5322 9764
rect 5338 9820 5402 9824
rect 5338 9764 5342 9820
rect 5342 9764 5398 9820
rect 5398 9764 5402 9820
rect 5338 9760 5402 9764
rect 8362 9820 8426 9824
rect 8362 9764 8366 9820
rect 8366 9764 8422 9820
rect 8422 9764 8426 9820
rect 8362 9760 8426 9764
rect 8442 9820 8506 9824
rect 8442 9764 8446 9820
rect 8446 9764 8502 9820
rect 8502 9764 8506 9820
rect 8442 9760 8506 9764
rect 8522 9820 8586 9824
rect 8522 9764 8526 9820
rect 8526 9764 8582 9820
rect 8582 9764 8586 9820
rect 8522 9760 8586 9764
rect 8602 9820 8666 9824
rect 8602 9764 8606 9820
rect 8606 9764 8662 9820
rect 8662 9764 8666 9820
rect 8602 9760 8666 9764
rect 3466 9276 3530 9280
rect 3466 9220 3470 9276
rect 3470 9220 3526 9276
rect 3526 9220 3530 9276
rect 3466 9216 3530 9220
rect 3546 9276 3610 9280
rect 3546 9220 3550 9276
rect 3550 9220 3606 9276
rect 3606 9220 3610 9276
rect 3546 9216 3610 9220
rect 3626 9276 3690 9280
rect 3626 9220 3630 9276
rect 3630 9220 3686 9276
rect 3686 9220 3690 9276
rect 3626 9216 3690 9220
rect 3706 9276 3770 9280
rect 3706 9220 3710 9276
rect 3710 9220 3766 9276
rect 3766 9220 3770 9276
rect 3706 9216 3770 9220
rect 6730 9276 6794 9280
rect 6730 9220 6734 9276
rect 6734 9220 6790 9276
rect 6790 9220 6794 9276
rect 6730 9216 6794 9220
rect 6810 9276 6874 9280
rect 6810 9220 6814 9276
rect 6814 9220 6870 9276
rect 6870 9220 6874 9276
rect 6810 9216 6874 9220
rect 6890 9276 6954 9280
rect 6890 9220 6894 9276
rect 6894 9220 6950 9276
rect 6950 9220 6954 9276
rect 6890 9216 6954 9220
rect 6970 9276 7034 9280
rect 6970 9220 6974 9276
rect 6974 9220 7030 9276
rect 7030 9220 7034 9276
rect 6970 9216 7034 9220
rect 1834 8732 1898 8736
rect 1834 8676 1838 8732
rect 1838 8676 1894 8732
rect 1894 8676 1898 8732
rect 1834 8672 1898 8676
rect 1914 8732 1978 8736
rect 1914 8676 1918 8732
rect 1918 8676 1974 8732
rect 1974 8676 1978 8732
rect 1914 8672 1978 8676
rect 1994 8732 2058 8736
rect 1994 8676 1998 8732
rect 1998 8676 2054 8732
rect 2054 8676 2058 8732
rect 1994 8672 2058 8676
rect 2074 8732 2138 8736
rect 2074 8676 2078 8732
rect 2078 8676 2134 8732
rect 2134 8676 2138 8732
rect 2074 8672 2138 8676
rect 5098 8732 5162 8736
rect 5098 8676 5102 8732
rect 5102 8676 5158 8732
rect 5158 8676 5162 8732
rect 5098 8672 5162 8676
rect 5178 8732 5242 8736
rect 5178 8676 5182 8732
rect 5182 8676 5238 8732
rect 5238 8676 5242 8732
rect 5178 8672 5242 8676
rect 5258 8732 5322 8736
rect 5258 8676 5262 8732
rect 5262 8676 5318 8732
rect 5318 8676 5322 8732
rect 5258 8672 5322 8676
rect 5338 8732 5402 8736
rect 5338 8676 5342 8732
rect 5342 8676 5398 8732
rect 5398 8676 5402 8732
rect 5338 8672 5402 8676
rect 8362 8732 8426 8736
rect 8362 8676 8366 8732
rect 8366 8676 8422 8732
rect 8422 8676 8426 8732
rect 8362 8672 8426 8676
rect 8442 8732 8506 8736
rect 8442 8676 8446 8732
rect 8446 8676 8502 8732
rect 8502 8676 8506 8732
rect 8442 8672 8506 8676
rect 8522 8732 8586 8736
rect 8522 8676 8526 8732
rect 8526 8676 8582 8732
rect 8582 8676 8586 8732
rect 8522 8672 8586 8676
rect 8602 8732 8666 8736
rect 8602 8676 8606 8732
rect 8606 8676 8662 8732
rect 8662 8676 8666 8732
rect 8602 8672 8666 8676
rect 3466 8188 3530 8192
rect 3466 8132 3470 8188
rect 3470 8132 3526 8188
rect 3526 8132 3530 8188
rect 3466 8128 3530 8132
rect 3546 8188 3610 8192
rect 3546 8132 3550 8188
rect 3550 8132 3606 8188
rect 3606 8132 3610 8188
rect 3546 8128 3610 8132
rect 3626 8188 3690 8192
rect 3626 8132 3630 8188
rect 3630 8132 3686 8188
rect 3686 8132 3690 8188
rect 3626 8128 3690 8132
rect 3706 8188 3770 8192
rect 3706 8132 3710 8188
rect 3710 8132 3766 8188
rect 3766 8132 3770 8188
rect 3706 8128 3770 8132
rect 6730 8188 6794 8192
rect 6730 8132 6734 8188
rect 6734 8132 6790 8188
rect 6790 8132 6794 8188
rect 6730 8128 6794 8132
rect 6810 8188 6874 8192
rect 6810 8132 6814 8188
rect 6814 8132 6870 8188
rect 6870 8132 6874 8188
rect 6810 8128 6874 8132
rect 6890 8188 6954 8192
rect 6890 8132 6894 8188
rect 6894 8132 6950 8188
rect 6950 8132 6954 8188
rect 6890 8128 6954 8132
rect 6970 8188 7034 8192
rect 6970 8132 6974 8188
rect 6974 8132 7030 8188
rect 7030 8132 7034 8188
rect 6970 8128 7034 8132
rect 1834 7644 1898 7648
rect 1834 7588 1838 7644
rect 1838 7588 1894 7644
rect 1894 7588 1898 7644
rect 1834 7584 1898 7588
rect 1914 7644 1978 7648
rect 1914 7588 1918 7644
rect 1918 7588 1974 7644
rect 1974 7588 1978 7644
rect 1914 7584 1978 7588
rect 1994 7644 2058 7648
rect 1994 7588 1998 7644
rect 1998 7588 2054 7644
rect 2054 7588 2058 7644
rect 1994 7584 2058 7588
rect 2074 7644 2138 7648
rect 2074 7588 2078 7644
rect 2078 7588 2134 7644
rect 2134 7588 2138 7644
rect 2074 7584 2138 7588
rect 5098 7644 5162 7648
rect 5098 7588 5102 7644
rect 5102 7588 5158 7644
rect 5158 7588 5162 7644
rect 5098 7584 5162 7588
rect 5178 7644 5242 7648
rect 5178 7588 5182 7644
rect 5182 7588 5238 7644
rect 5238 7588 5242 7644
rect 5178 7584 5242 7588
rect 5258 7644 5322 7648
rect 5258 7588 5262 7644
rect 5262 7588 5318 7644
rect 5318 7588 5322 7644
rect 5258 7584 5322 7588
rect 5338 7644 5402 7648
rect 5338 7588 5342 7644
rect 5342 7588 5398 7644
rect 5398 7588 5402 7644
rect 5338 7584 5402 7588
rect 8362 7644 8426 7648
rect 8362 7588 8366 7644
rect 8366 7588 8422 7644
rect 8422 7588 8426 7644
rect 8362 7584 8426 7588
rect 8442 7644 8506 7648
rect 8442 7588 8446 7644
rect 8446 7588 8502 7644
rect 8502 7588 8506 7644
rect 8442 7584 8506 7588
rect 8522 7644 8586 7648
rect 8522 7588 8526 7644
rect 8526 7588 8582 7644
rect 8582 7588 8586 7644
rect 8522 7584 8586 7588
rect 8602 7644 8666 7648
rect 8602 7588 8606 7644
rect 8606 7588 8662 7644
rect 8662 7588 8666 7644
rect 8602 7584 8666 7588
rect 3466 7100 3530 7104
rect 3466 7044 3470 7100
rect 3470 7044 3526 7100
rect 3526 7044 3530 7100
rect 3466 7040 3530 7044
rect 3546 7100 3610 7104
rect 3546 7044 3550 7100
rect 3550 7044 3606 7100
rect 3606 7044 3610 7100
rect 3546 7040 3610 7044
rect 3626 7100 3690 7104
rect 3626 7044 3630 7100
rect 3630 7044 3686 7100
rect 3686 7044 3690 7100
rect 3626 7040 3690 7044
rect 3706 7100 3770 7104
rect 3706 7044 3710 7100
rect 3710 7044 3766 7100
rect 3766 7044 3770 7100
rect 3706 7040 3770 7044
rect 6730 7100 6794 7104
rect 6730 7044 6734 7100
rect 6734 7044 6790 7100
rect 6790 7044 6794 7100
rect 6730 7040 6794 7044
rect 6810 7100 6874 7104
rect 6810 7044 6814 7100
rect 6814 7044 6870 7100
rect 6870 7044 6874 7100
rect 6810 7040 6874 7044
rect 6890 7100 6954 7104
rect 6890 7044 6894 7100
rect 6894 7044 6950 7100
rect 6950 7044 6954 7100
rect 6890 7040 6954 7044
rect 6970 7100 7034 7104
rect 6970 7044 6974 7100
rect 6974 7044 7030 7100
rect 7030 7044 7034 7100
rect 6970 7040 7034 7044
rect 1834 6556 1898 6560
rect 1834 6500 1838 6556
rect 1838 6500 1894 6556
rect 1894 6500 1898 6556
rect 1834 6496 1898 6500
rect 1914 6556 1978 6560
rect 1914 6500 1918 6556
rect 1918 6500 1974 6556
rect 1974 6500 1978 6556
rect 1914 6496 1978 6500
rect 1994 6556 2058 6560
rect 1994 6500 1998 6556
rect 1998 6500 2054 6556
rect 2054 6500 2058 6556
rect 1994 6496 2058 6500
rect 2074 6556 2138 6560
rect 2074 6500 2078 6556
rect 2078 6500 2134 6556
rect 2134 6500 2138 6556
rect 2074 6496 2138 6500
rect 5098 6556 5162 6560
rect 5098 6500 5102 6556
rect 5102 6500 5158 6556
rect 5158 6500 5162 6556
rect 5098 6496 5162 6500
rect 5178 6556 5242 6560
rect 5178 6500 5182 6556
rect 5182 6500 5238 6556
rect 5238 6500 5242 6556
rect 5178 6496 5242 6500
rect 5258 6556 5322 6560
rect 5258 6500 5262 6556
rect 5262 6500 5318 6556
rect 5318 6500 5322 6556
rect 5258 6496 5322 6500
rect 5338 6556 5402 6560
rect 5338 6500 5342 6556
rect 5342 6500 5398 6556
rect 5398 6500 5402 6556
rect 5338 6496 5402 6500
rect 8362 6556 8426 6560
rect 8362 6500 8366 6556
rect 8366 6500 8422 6556
rect 8422 6500 8426 6556
rect 8362 6496 8426 6500
rect 8442 6556 8506 6560
rect 8442 6500 8446 6556
rect 8446 6500 8502 6556
rect 8502 6500 8506 6556
rect 8442 6496 8506 6500
rect 8522 6556 8586 6560
rect 8522 6500 8526 6556
rect 8526 6500 8582 6556
rect 8582 6500 8586 6556
rect 8522 6496 8586 6500
rect 8602 6556 8666 6560
rect 8602 6500 8606 6556
rect 8606 6500 8662 6556
rect 8662 6500 8666 6556
rect 8602 6496 8666 6500
rect 3466 6012 3530 6016
rect 3466 5956 3470 6012
rect 3470 5956 3526 6012
rect 3526 5956 3530 6012
rect 3466 5952 3530 5956
rect 3546 6012 3610 6016
rect 3546 5956 3550 6012
rect 3550 5956 3606 6012
rect 3606 5956 3610 6012
rect 3546 5952 3610 5956
rect 3626 6012 3690 6016
rect 3626 5956 3630 6012
rect 3630 5956 3686 6012
rect 3686 5956 3690 6012
rect 3626 5952 3690 5956
rect 3706 6012 3770 6016
rect 3706 5956 3710 6012
rect 3710 5956 3766 6012
rect 3766 5956 3770 6012
rect 3706 5952 3770 5956
rect 6730 6012 6794 6016
rect 6730 5956 6734 6012
rect 6734 5956 6790 6012
rect 6790 5956 6794 6012
rect 6730 5952 6794 5956
rect 6810 6012 6874 6016
rect 6810 5956 6814 6012
rect 6814 5956 6870 6012
rect 6870 5956 6874 6012
rect 6810 5952 6874 5956
rect 6890 6012 6954 6016
rect 6890 5956 6894 6012
rect 6894 5956 6950 6012
rect 6950 5956 6954 6012
rect 6890 5952 6954 5956
rect 6970 6012 7034 6016
rect 6970 5956 6974 6012
rect 6974 5956 7030 6012
rect 7030 5956 7034 6012
rect 6970 5952 7034 5956
rect 1834 5468 1898 5472
rect 1834 5412 1838 5468
rect 1838 5412 1894 5468
rect 1894 5412 1898 5468
rect 1834 5408 1898 5412
rect 1914 5468 1978 5472
rect 1914 5412 1918 5468
rect 1918 5412 1974 5468
rect 1974 5412 1978 5468
rect 1914 5408 1978 5412
rect 1994 5468 2058 5472
rect 1994 5412 1998 5468
rect 1998 5412 2054 5468
rect 2054 5412 2058 5468
rect 1994 5408 2058 5412
rect 2074 5468 2138 5472
rect 2074 5412 2078 5468
rect 2078 5412 2134 5468
rect 2134 5412 2138 5468
rect 2074 5408 2138 5412
rect 5098 5468 5162 5472
rect 5098 5412 5102 5468
rect 5102 5412 5158 5468
rect 5158 5412 5162 5468
rect 5098 5408 5162 5412
rect 5178 5468 5242 5472
rect 5178 5412 5182 5468
rect 5182 5412 5238 5468
rect 5238 5412 5242 5468
rect 5178 5408 5242 5412
rect 5258 5468 5322 5472
rect 5258 5412 5262 5468
rect 5262 5412 5318 5468
rect 5318 5412 5322 5468
rect 5258 5408 5322 5412
rect 5338 5468 5402 5472
rect 5338 5412 5342 5468
rect 5342 5412 5398 5468
rect 5398 5412 5402 5468
rect 5338 5408 5402 5412
rect 8362 5468 8426 5472
rect 8362 5412 8366 5468
rect 8366 5412 8422 5468
rect 8422 5412 8426 5468
rect 8362 5408 8426 5412
rect 8442 5468 8506 5472
rect 8442 5412 8446 5468
rect 8446 5412 8502 5468
rect 8502 5412 8506 5468
rect 8442 5408 8506 5412
rect 8522 5468 8586 5472
rect 8522 5412 8526 5468
rect 8526 5412 8582 5468
rect 8582 5412 8586 5468
rect 8522 5408 8586 5412
rect 8602 5468 8666 5472
rect 8602 5412 8606 5468
rect 8606 5412 8662 5468
rect 8662 5412 8666 5468
rect 8602 5408 8666 5412
rect 3466 4924 3530 4928
rect 3466 4868 3470 4924
rect 3470 4868 3526 4924
rect 3526 4868 3530 4924
rect 3466 4864 3530 4868
rect 3546 4924 3610 4928
rect 3546 4868 3550 4924
rect 3550 4868 3606 4924
rect 3606 4868 3610 4924
rect 3546 4864 3610 4868
rect 3626 4924 3690 4928
rect 3626 4868 3630 4924
rect 3630 4868 3686 4924
rect 3686 4868 3690 4924
rect 3626 4864 3690 4868
rect 3706 4924 3770 4928
rect 3706 4868 3710 4924
rect 3710 4868 3766 4924
rect 3766 4868 3770 4924
rect 3706 4864 3770 4868
rect 6730 4924 6794 4928
rect 6730 4868 6734 4924
rect 6734 4868 6790 4924
rect 6790 4868 6794 4924
rect 6730 4864 6794 4868
rect 6810 4924 6874 4928
rect 6810 4868 6814 4924
rect 6814 4868 6870 4924
rect 6870 4868 6874 4924
rect 6810 4864 6874 4868
rect 6890 4924 6954 4928
rect 6890 4868 6894 4924
rect 6894 4868 6950 4924
rect 6950 4868 6954 4924
rect 6890 4864 6954 4868
rect 6970 4924 7034 4928
rect 6970 4868 6974 4924
rect 6974 4868 7030 4924
rect 7030 4868 7034 4924
rect 6970 4864 7034 4868
rect 1834 4380 1898 4384
rect 1834 4324 1838 4380
rect 1838 4324 1894 4380
rect 1894 4324 1898 4380
rect 1834 4320 1898 4324
rect 1914 4380 1978 4384
rect 1914 4324 1918 4380
rect 1918 4324 1974 4380
rect 1974 4324 1978 4380
rect 1914 4320 1978 4324
rect 1994 4380 2058 4384
rect 1994 4324 1998 4380
rect 1998 4324 2054 4380
rect 2054 4324 2058 4380
rect 1994 4320 2058 4324
rect 2074 4380 2138 4384
rect 2074 4324 2078 4380
rect 2078 4324 2134 4380
rect 2134 4324 2138 4380
rect 2074 4320 2138 4324
rect 5098 4380 5162 4384
rect 5098 4324 5102 4380
rect 5102 4324 5158 4380
rect 5158 4324 5162 4380
rect 5098 4320 5162 4324
rect 5178 4380 5242 4384
rect 5178 4324 5182 4380
rect 5182 4324 5238 4380
rect 5238 4324 5242 4380
rect 5178 4320 5242 4324
rect 5258 4380 5322 4384
rect 5258 4324 5262 4380
rect 5262 4324 5318 4380
rect 5318 4324 5322 4380
rect 5258 4320 5322 4324
rect 5338 4380 5402 4384
rect 5338 4324 5342 4380
rect 5342 4324 5398 4380
rect 5398 4324 5402 4380
rect 5338 4320 5402 4324
rect 8362 4380 8426 4384
rect 8362 4324 8366 4380
rect 8366 4324 8422 4380
rect 8422 4324 8426 4380
rect 8362 4320 8426 4324
rect 8442 4380 8506 4384
rect 8442 4324 8446 4380
rect 8446 4324 8502 4380
rect 8502 4324 8506 4380
rect 8442 4320 8506 4324
rect 8522 4380 8586 4384
rect 8522 4324 8526 4380
rect 8526 4324 8582 4380
rect 8582 4324 8586 4380
rect 8522 4320 8586 4324
rect 8602 4380 8666 4384
rect 8602 4324 8606 4380
rect 8606 4324 8662 4380
rect 8662 4324 8666 4380
rect 8602 4320 8666 4324
rect 3466 3836 3530 3840
rect 3466 3780 3470 3836
rect 3470 3780 3526 3836
rect 3526 3780 3530 3836
rect 3466 3776 3530 3780
rect 3546 3836 3610 3840
rect 3546 3780 3550 3836
rect 3550 3780 3606 3836
rect 3606 3780 3610 3836
rect 3546 3776 3610 3780
rect 3626 3836 3690 3840
rect 3626 3780 3630 3836
rect 3630 3780 3686 3836
rect 3686 3780 3690 3836
rect 3626 3776 3690 3780
rect 3706 3836 3770 3840
rect 3706 3780 3710 3836
rect 3710 3780 3766 3836
rect 3766 3780 3770 3836
rect 3706 3776 3770 3780
rect 6730 3836 6794 3840
rect 6730 3780 6734 3836
rect 6734 3780 6790 3836
rect 6790 3780 6794 3836
rect 6730 3776 6794 3780
rect 6810 3836 6874 3840
rect 6810 3780 6814 3836
rect 6814 3780 6870 3836
rect 6870 3780 6874 3836
rect 6810 3776 6874 3780
rect 6890 3836 6954 3840
rect 6890 3780 6894 3836
rect 6894 3780 6950 3836
rect 6950 3780 6954 3836
rect 6890 3776 6954 3780
rect 6970 3836 7034 3840
rect 6970 3780 6974 3836
rect 6974 3780 7030 3836
rect 7030 3780 7034 3836
rect 6970 3776 7034 3780
rect 1834 3292 1898 3296
rect 1834 3236 1838 3292
rect 1838 3236 1894 3292
rect 1894 3236 1898 3292
rect 1834 3232 1898 3236
rect 1914 3292 1978 3296
rect 1914 3236 1918 3292
rect 1918 3236 1974 3292
rect 1974 3236 1978 3292
rect 1914 3232 1978 3236
rect 1994 3292 2058 3296
rect 1994 3236 1998 3292
rect 1998 3236 2054 3292
rect 2054 3236 2058 3292
rect 1994 3232 2058 3236
rect 2074 3292 2138 3296
rect 2074 3236 2078 3292
rect 2078 3236 2134 3292
rect 2134 3236 2138 3292
rect 2074 3232 2138 3236
rect 5098 3292 5162 3296
rect 5098 3236 5102 3292
rect 5102 3236 5158 3292
rect 5158 3236 5162 3292
rect 5098 3232 5162 3236
rect 5178 3292 5242 3296
rect 5178 3236 5182 3292
rect 5182 3236 5238 3292
rect 5238 3236 5242 3292
rect 5178 3232 5242 3236
rect 5258 3292 5322 3296
rect 5258 3236 5262 3292
rect 5262 3236 5318 3292
rect 5318 3236 5322 3292
rect 5258 3232 5322 3236
rect 5338 3292 5402 3296
rect 5338 3236 5342 3292
rect 5342 3236 5398 3292
rect 5398 3236 5402 3292
rect 5338 3232 5402 3236
rect 8362 3292 8426 3296
rect 8362 3236 8366 3292
rect 8366 3236 8422 3292
rect 8422 3236 8426 3292
rect 8362 3232 8426 3236
rect 8442 3292 8506 3296
rect 8442 3236 8446 3292
rect 8446 3236 8502 3292
rect 8502 3236 8506 3292
rect 8442 3232 8506 3236
rect 8522 3292 8586 3296
rect 8522 3236 8526 3292
rect 8526 3236 8582 3292
rect 8582 3236 8586 3292
rect 8522 3232 8586 3236
rect 8602 3292 8666 3296
rect 8602 3236 8606 3292
rect 8606 3236 8662 3292
rect 8662 3236 8666 3292
rect 8602 3232 8666 3236
rect 3466 2748 3530 2752
rect 3466 2692 3470 2748
rect 3470 2692 3526 2748
rect 3526 2692 3530 2748
rect 3466 2688 3530 2692
rect 3546 2748 3610 2752
rect 3546 2692 3550 2748
rect 3550 2692 3606 2748
rect 3606 2692 3610 2748
rect 3546 2688 3610 2692
rect 3626 2748 3690 2752
rect 3626 2692 3630 2748
rect 3630 2692 3686 2748
rect 3686 2692 3690 2748
rect 3626 2688 3690 2692
rect 3706 2748 3770 2752
rect 3706 2692 3710 2748
rect 3710 2692 3766 2748
rect 3766 2692 3770 2748
rect 3706 2688 3770 2692
rect 6730 2748 6794 2752
rect 6730 2692 6734 2748
rect 6734 2692 6790 2748
rect 6790 2692 6794 2748
rect 6730 2688 6794 2692
rect 6810 2748 6874 2752
rect 6810 2692 6814 2748
rect 6814 2692 6870 2748
rect 6870 2692 6874 2748
rect 6810 2688 6874 2692
rect 6890 2748 6954 2752
rect 6890 2692 6894 2748
rect 6894 2692 6950 2748
rect 6950 2692 6954 2748
rect 6890 2688 6954 2692
rect 6970 2748 7034 2752
rect 6970 2692 6974 2748
rect 6974 2692 7030 2748
rect 7030 2692 7034 2748
rect 6970 2688 7034 2692
rect 1834 2204 1898 2208
rect 1834 2148 1838 2204
rect 1838 2148 1894 2204
rect 1894 2148 1898 2204
rect 1834 2144 1898 2148
rect 1914 2204 1978 2208
rect 1914 2148 1918 2204
rect 1918 2148 1974 2204
rect 1974 2148 1978 2204
rect 1914 2144 1978 2148
rect 1994 2204 2058 2208
rect 1994 2148 1998 2204
rect 1998 2148 2054 2204
rect 2054 2148 2058 2204
rect 1994 2144 2058 2148
rect 2074 2204 2138 2208
rect 2074 2148 2078 2204
rect 2078 2148 2134 2204
rect 2134 2148 2138 2204
rect 2074 2144 2138 2148
rect 5098 2204 5162 2208
rect 5098 2148 5102 2204
rect 5102 2148 5158 2204
rect 5158 2148 5162 2204
rect 5098 2144 5162 2148
rect 5178 2204 5242 2208
rect 5178 2148 5182 2204
rect 5182 2148 5238 2204
rect 5238 2148 5242 2204
rect 5178 2144 5242 2148
rect 5258 2204 5322 2208
rect 5258 2148 5262 2204
rect 5262 2148 5318 2204
rect 5318 2148 5322 2204
rect 5258 2144 5322 2148
rect 5338 2204 5402 2208
rect 5338 2148 5342 2204
rect 5342 2148 5398 2204
rect 5398 2148 5402 2204
rect 5338 2144 5402 2148
rect 8362 2204 8426 2208
rect 8362 2148 8366 2204
rect 8366 2148 8422 2204
rect 8422 2148 8426 2204
rect 8362 2144 8426 2148
rect 8442 2204 8506 2208
rect 8442 2148 8446 2204
rect 8446 2148 8502 2204
rect 8502 2148 8506 2204
rect 8442 2144 8506 2148
rect 8522 2204 8586 2208
rect 8522 2148 8526 2204
rect 8526 2148 8582 2204
rect 8582 2148 8586 2204
rect 8522 2144 8586 2148
rect 8602 2204 8666 2208
rect 8602 2148 8606 2204
rect 8606 2148 8662 2204
rect 8662 2148 8666 2204
rect 8602 2144 8666 2148
<< metal4 >>
rect 1826 10912 2146 11472
rect 1826 10848 1834 10912
rect 1898 10848 1914 10912
rect 1978 10848 1994 10912
rect 2058 10848 2074 10912
rect 2138 10848 2146 10912
rect 1826 9824 2146 10848
rect 1826 9760 1834 9824
rect 1898 9760 1914 9824
rect 1978 9760 1994 9824
rect 2058 9760 2074 9824
rect 2138 9760 2146 9824
rect 1826 8736 2146 9760
rect 1826 8672 1834 8736
rect 1898 8672 1914 8736
rect 1978 8672 1994 8736
rect 2058 8672 2074 8736
rect 2138 8672 2146 8736
rect 1826 7648 2146 8672
rect 1826 7584 1834 7648
rect 1898 7584 1914 7648
rect 1978 7584 1994 7648
rect 2058 7584 2074 7648
rect 2138 7584 2146 7648
rect 1826 6560 2146 7584
rect 1826 6496 1834 6560
rect 1898 6496 1914 6560
rect 1978 6496 1994 6560
rect 2058 6496 2074 6560
rect 2138 6496 2146 6560
rect 1826 5472 2146 6496
rect 1826 5408 1834 5472
rect 1898 5408 1914 5472
rect 1978 5408 1994 5472
rect 2058 5408 2074 5472
rect 2138 5408 2146 5472
rect 1826 4384 2146 5408
rect 1826 4320 1834 4384
rect 1898 4320 1914 4384
rect 1978 4320 1994 4384
rect 2058 4320 2074 4384
rect 2138 4320 2146 4384
rect 1826 3296 2146 4320
rect 1826 3232 1834 3296
rect 1898 3232 1914 3296
rect 1978 3232 1994 3296
rect 2058 3232 2074 3296
rect 2138 3232 2146 3296
rect 1826 2208 2146 3232
rect 1826 2144 1834 2208
rect 1898 2144 1914 2208
rect 1978 2144 1994 2208
rect 2058 2144 2074 2208
rect 2138 2144 2146 2208
rect 1826 2128 2146 2144
rect 3458 11456 3778 11472
rect 3458 11392 3466 11456
rect 3530 11392 3546 11456
rect 3610 11392 3626 11456
rect 3690 11392 3706 11456
rect 3770 11392 3778 11456
rect 3458 10368 3778 11392
rect 3458 10304 3466 10368
rect 3530 10304 3546 10368
rect 3610 10304 3626 10368
rect 3690 10304 3706 10368
rect 3770 10304 3778 10368
rect 3458 9280 3778 10304
rect 3458 9216 3466 9280
rect 3530 9216 3546 9280
rect 3610 9216 3626 9280
rect 3690 9216 3706 9280
rect 3770 9216 3778 9280
rect 3458 8192 3778 9216
rect 3458 8128 3466 8192
rect 3530 8128 3546 8192
rect 3610 8128 3626 8192
rect 3690 8128 3706 8192
rect 3770 8128 3778 8192
rect 3458 7104 3778 8128
rect 3458 7040 3466 7104
rect 3530 7040 3546 7104
rect 3610 7040 3626 7104
rect 3690 7040 3706 7104
rect 3770 7040 3778 7104
rect 3458 6016 3778 7040
rect 3458 5952 3466 6016
rect 3530 5952 3546 6016
rect 3610 5952 3626 6016
rect 3690 5952 3706 6016
rect 3770 5952 3778 6016
rect 3458 4928 3778 5952
rect 3458 4864 3466 4928
rect 3530 4864 3546 4928
rect 3610 4864 3626 4928
rect 3690 4864 3706 4928
rect 3770 4864 3778 4928
rect 3458 3840 3778 4864
rect 3458 3776 3466 3840
rect 3530 3776 3546 3840
rect 3610 3776 3626 3840
rect 3690 3776 3706 3840
rect 3770 3776 3778 3840
rect 3458 2752 3778 3776
rect 3458 2688 3466 2752
rect 3530 2688 3546 2752
rect 3610 2688 3626 2752
rect 3690 2688 3706 2752
rect 3770 2688 3778 2752
rect 3458 2128 3778 2688
rect 5090 10912 5410 11472
rect 5090 10848 5098 10912
rect 5162 10848 5178 10912
rect 5242 10848 5258 10912
rect 5322 10848 5338 10912
rect 5402 10848 5410 10912
rect 5090 9824 5410 10848
rect 5090 9760 5098 9824
rect 5162 9760 5178 9824
rect 5242 9760 5258 9824
rect 5322 9760 5338 9824
rect 5402 9760 5410 9824
rect 5090 8736 5410 9760
rect 5090 8672 5098 8736
rect 5162 8672 5178 8736
rect 5242 8672 5258 8736
rect 5322 8672 5338 8736
rect 5402 8672 5410 8736
rect 5090 7648 5410 8672
rect 5090 7584 5098 7648
rect 5162 7584 5178 7648
rect 5242 7584 5258 7648
rect 5322 7584 5338 7648
rect 5402 7584 5410 7648
rect 5090 6560 5410 7584
rect 5090 6496 5098 6560
rect 5162 6496 5178 6560
rect 5242 6496 5258 6560
rect 5322 6496 5338 6560
rect 5402 6496 5410 6560
rect 5090 5472 5410 6496
rect 5090 5408 5098 5472
rect 5162 5408 5178 5472
rect 5242 5408 5258 5472
rect 5322 5408 5338 5472
rect 5402 5408 5410 5472
rect 5090 4384 5410 5408
rect 5090 4320 5098 4384
rect 5162 4320 5178 4384
rect 5242 4320 5258 4384
rect 5322 4320 5338 4384
rect 5402 4320 5410 4384
rect 5090 3296 5410 4320
rect 5090 3232 5098 3296
rect 5162 3232 5178 3296
rect 5242 3232 5258 3296
rect 5322 3232 5338 3296
rect 5402 3232 5410 3296
rect 5090 2208 5410 3232
rect 5090 2144 5098 2208
rect 5162 2144 5178 2208
rect 5242 2144 5258 2208
rect 5322 2144 5338 2208
rect 5402 2144 5410 2208
rect 5090 2128 5410 2144
rect 6722 11456 7042 11472
rect 6722 11392 6730 11456
rect 6794 11392 6810 11456
rect 6874 11392 6890 11456
rect 6954 11392 6970 11456
rect 7034 11392 7042 11456
rect 6722 10368 7042 11392
rect 6722 10304 6730 10368
rect 6794 10304 6810 10368
rect 6874 10304 6890 10368
rect 6954 10304 6970 10368
rect 7034 10304 7042 10368
rect 6722 9280 7042 10304
rect 6722 9216 6730 9280
rect 6794 9216 6810 9280
rect 6874 9216 6890 9280
rect 6954 9216 6970 9280
rect 7034 9216 7042 9280
rect 6722 8192 7042 9216
rect 6722 8128 6730 8192
rect 6794 8128 6810 8192
rect 6874 8128 6890 8192
rect 6954 8128 6970 8192
rect 7034 8128 7042 8192
rect 6722 7104 7042 8128
rect 6722 7040 6730 7104
rect 6794 7040 6810 7104
rect 6874 7040 6890 7104
rect 6954 7040 6970 7104
rect 7034 7040 7042 7104
rect 6722 6016 7042 7040
rect 6722 5952 6730 6016
rect 6794 5952 6810 6016
rect 6874 5952 6890 6016
rect 6954 5952 6970 6016
rect 7034 5952 7042 6016
rect 6722 4928 7042 5952
rect 6722 4864 6730 4928
rect 6794 4864 6810 4928
rect 6874 4864 6890 4928
rect 6954 4864 6970 4928
rect 7034 4864 7042 4928
rect 6722 3840 7042 4864
rect 6722 3776 6730 3840
rect 6794 3776 6810 3840
rect 6874 3776 6890 3840
rect 6954 3776 6970 3840
rect 7034 3776 7042 3840
rect 6722 2752 7042 3776
rect 6722 2688 6730 2752
rect 6794 2688 6810 2752
rect 6874 2688 6890 2752
rect 6954 2688 6970 2752
rect 7034 2688 7042 2752
rect 6722 2128 7042 2688
rect 8354 10912 8674 11472
rect 8354 10848 8362 10912
rect 8426 10848 8442 10912
rect 8506 10848 8522 10912
rect 8586 10848 8602 10912
rect 8666 10848 8674 10912
rect 8354 9824 8674 10848
rect 8354 9760 8362 9824
rect 8426 9760 8442 9824
rect 8506 9760 8522 9824
rect 8586 9760 8602 9824
rect 8666 9760 8674 9824
rect 8354 8736 8674 9760
rect 8354 8672 8362 8736
rect 8426 8672 8442 8736
rect 8506 8672 8522 8736
rect 8586 8672 8602 8736
rect 8666 8672 8674 8736
rect 8354 7648 8674 8672
rect 8354 7584 8362 7648
rect 8426 7584 8442 7648
rect 8506 7584 8522 7648
rect 8586 7584 8602 7648
rect 8666 7584 8674 7648
rect 8354 6560 8674 7584
rect 8354 6496 8362 6560
rect 8426 6496 8442 6560
rect 8506 6496 8522 6560
rect 8586 6496 8602 6560
rect 8666 6496 8674 6560
rect 8354 5472 8674 6496
rect 8354 5408 8362 5472
rect 8426 5408 8442 5472
rect 8506 5408 8522 5472
rect 8586 5408 8602 5472
rect 8666 5408 8674 5472
rect 8354 4384 8674 5408
rect 8354 4320 8362 4384
rect 8426 4320 8442 4384
rect 8506 4320 8522 4384
rect 8586 4320 8602 4384
rect 8666 4320 8674 4384
rect 8354 3296 8674 4320
rect 8354 3232 8362 3296
rect 8426 3232 8442 3296
rect 8506 3232 8522 3296
rect 8586 3232 8602 3296
rect 8666 3232 8674 3296
rect 8354 2208 8674 3232
rect 8354 2144 8362 2208
rect 8426 2144 8442 2208
rect 8506 2144 8522 2208
rect 8586 2144 8602 2208
rect 8666 2144 8674 2208
rect 8354 2128 8674 2144
use sky130_fd_sc_hd__decap_12  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 630 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1608910539
transform 1 0 630 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 354 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 354 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1608910539
transform 1 0 1734 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1608910539
transform 1 0 1734 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1608910539
transform 1 0 2838 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1608910539
transform 1 0 3298 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2838 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3206 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5046 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1608910539
transform 1 0 3942 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1608910539
transform 1 0 4402 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1608910539
transform 1 0 6058 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5782 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1608910539
transform 1 0 6150 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 5506 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1608910539
transform 1 0 5966 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1608910539
transform 1 0 6058 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1608910539
transform 1 0 7162 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1608910539
transform 1 0 7254 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_88
timestamp 1608910539
transform 1 0 8450 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_82
timestamp 1608910539
transform 1 0 7898 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1608910539
transform 1 0 8358 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  conb_1\[7\] tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 8174 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_100
timestamp 1608910539
transform 1 0 9554 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_102 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9738 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_94
timestamp 1608910539
transform 1 0 9002 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1608910539
transform 1 0 8910 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 10106 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 10106 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1608910539
transform 1 0 630 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 354 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1608910539
transform 1 0 2194 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_15
timestamp 1608910539
transform 1 0 1734 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  conb_1\[0\]
timestamp 1608910539
transform 1 0 1918 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_35
timestamp 1608910539
transform 1 0 3574 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 1608910539
transform 1 0 2930 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1608910539
transform 1 0 3206 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  conb_1\[2\]
timestamp 1608910539
transform 1 0 3298 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_46
timestamp 1608910539
transform 1 0 4586 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  conb_1\[3\]
timestamp 1608910539
transform 1 0 4310 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1608910539
transform 1 0 6058 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp 1608910539
transform 1 0 5690 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  conb_1\[4\]
timestamp 1608910539
transform 1 0 5782 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1608910539
transform 1 0 7162 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  conb_1\[5\]
timestamp 1608910539
transform 1 0 7254 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_78
timestamp 1608910539
transform 1 0 7530 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1608910539
transform 1 0 9646 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1608910539
transform 1 0 8910 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1608910539
transform 1 0 8634 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1608910539
transform 1 0 8818 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 10106 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1608910539
transform 1 0 630 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 354 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_20
timestamp 1608910539
transform 1 0 2194 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 1608910539
transform 1 0 1734 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  conb_1\[1\]
timestamp 1608910539
transform 1 0 1918 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1608910539
transform 1 0 3298 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1608910539
transform 1 0 4402 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1608910539
transform 1 0 6058 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 5874 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_56
timestamp 1608910539
transform 1 0 5506 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1608910539
transform 1 0 5966 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_74
timestamp 1608910539
transform 1 0 7162 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_88
timestamp 1608910539
transform 1 0 8450 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_82
timestamp 1608910539
transform 1 0 7898 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  conb_1\[6\]
timestamp 1608910539
transform 1 0 8174 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_100
timestamp 1608910539
transform 1 0 9554 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 10106 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1608910539
transform 1 0 630 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 354 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1608910539
transform 1 0 1734 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1608910539
transform 1 0 3298 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1608910539
transform 1 0 2838 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1608910539
transform 1 0 3206 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1608910539
transform 1 0 4402 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1608910539
transform 1 0 5506 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1608910539
transform 1 0 6610 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1608910539
transform 1 0 7714 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1608910539
transform 1 0 9646 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1608910539
transform 1 0 8910 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1608910539
transform 1 0 8818 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 10106 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1608910539
transform 1 0 630 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 354 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1608910539
transform 1 0 1734 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1608910539
transform 1 0 2838 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1608910539
transform 1 0 5046 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1608910539
transform 1 0 3942 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1608910539
transform 1 0 6058 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1608910539
transform 1 0 5782 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1608910539
transform 1 0 5966 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1608910539
transform 1 0 7162 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1608910539
transform 1 0 8266 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_102
timestamp 1608910539
transform 1 0 9738 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1608910539
transform 1 0 9370 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 10106 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1608910539
transform 1 0 630 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1608910539
transform 1 0 630 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 354 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 354 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1608910539
transform 1 0 1734 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1608910539
transform 1 0 1734 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1608910539
transform 1 0 2838 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1608910539
transform 1 0 3298 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1608910539
transform 1 0 2838 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1608910539
transform 1 0 3206 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1608910539
transform 1 0 5046 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1608910539
transform 1 0 3942 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1608910539
transform 1 0 4402 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1608910539
transform 1 0 6058 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1608910539
transform 1 0 5782 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1608910539
transform 1 0 5506 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1608910539
transform 1 0 5966 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1608910539
transform 1 0 7162 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1608910539
transform 1 0 6610 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1608910539
transform 1 0 8266 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1608910539
transform 1 0 7714 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1608910539
transform 1 0 9738 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1608910539
transform 1 0 9370 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_101
timestamp 1608910539
transform 1 0 9646 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1608910539
transform 1 0 8910 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1608910539
transform 1 0 8818 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 10106 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 10106 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1608910539
transform 1 0 630 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 354 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1608910539
transform 1 0 1734 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1608910539
transform 1 0 3298 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1608910539
transform 1 0 2838 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608910539
transform 1 0 3206 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1608910539
transform 1 0 4402 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1608910539
transform 1 0 5506 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1608910539
transform 1 0 6610 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1608910539
transform 1 0 7714 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1608910539
transform 1 0 9646 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1608910539
transform 1 0 8910 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608910539
transform 1 0 8818 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 10106 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1608910539
transform 1 0 630 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 354 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1608910539
transform 1 0 1734 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1608910539
transform 1 0 2838 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1608910539
transform 1 0 5046 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1608910539
transform 1 0 3942 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1608910539
transform 1 0 6058 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1608910539
transform 1 0 5782 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608910539
transform 1 0 5966 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1608910539
transform 1 0 7162 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1608910539
transform 1 0 8266 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1608910539
transform 1 0 9738 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1608910539
transform 1 0 9370 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 10106 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1608910539
transform 1 0 630 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 354 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1608910539
transform 1 0 1734 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1608910539
transform 1 0 3298 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1608910539
transform 1 0 2838 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608910539
transform 1 0 3206 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1608910539
transform 1 0 4402 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1608910539
transform 1 0 5506 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1608910539
transform 1 0 6610 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1608910539
transform 1 0 7714 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1608910539
transform 1 0 9646 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1608910539
transform 1 0 8910 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608910539
transform 1 0 8818 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 10106 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1608910539
transform 1 0 630 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 354 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1608910539
transform 1 0 1734 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1608910539
transform 1 0 2838 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1608910539
transform 1 0 5046 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1608910539
transform 1 0 3942 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1608910539
transform 1 0 6058 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1608910539
transform 1 0 5782 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608910539
transform 1 0 5966 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1608910539
transform 1 0 7162 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1608910539
transform 1 0 8266 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_102
timestamp 1608910539
transform 1 0 9738 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_98
timestamp 1608910539
transform 1 0 9370 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 10106 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1608910539
transform 1 0 630 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 354 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1608910539
transform 1 0 1734 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1608910539
transform 1 0 3298 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1608910539
transform 1 0 2838 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608910539
transform 1 0 3206 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1608910539
transform 1 0 4402 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1608910539
transform 1 0 5506 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1608910539
transform 1 0 6610 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1608910539
transform 1 0 7714 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1608910539
transform 1 0 9646 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1608910539
transform 1 0 8910 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608910539
transform 1 0 8818 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 10106 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1608910539
transform 1 0 630 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1608910539
transform 1 0 630 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 354 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 354 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1608910539
transform 1 0 1734 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1608910539
transform 1 0 1734 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1608910539
transform 1 0 3298 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1608910539
transform 1 0 2838 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1608910539
transform 1 0 2838 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608910539
transform 1 0 3206 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1608910539
transform 1 0 4402 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1608910539
transform 1 0 5046 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1608910539
transform 1 0 3942 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1608910539
transform 1 0 5506 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1608910539
transform 1 0 6058 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1608910539
transform 1 0 5782 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608910539
transform 1 0 5966 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1608910539
transform 1 0 6610 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1608910539
transform 1 0 7162 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1608910539
transform 1 0 7714 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1608910539
transform 1 0 8266 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_101
timestamp 1608910539
transform 1 0 9646 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_93
timestamp 1608910539
transform 1 0 8910 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_102
timestamp 1608910539
transform 1 0 9738 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_98
timestamp 1608910539
transform 1 0 9370 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 8818 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 10106 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 10106 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1608910539
transform 1 0 630 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 354 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1608910539
transform 1 0 1734 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1608910539
transform 1 0 2838 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1608910539
transform 1 0 5046 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1608910539
transform 1 0 3942 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1608910539
transform 1 0 6058 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1608910539
transform 1 0 5782 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 5966 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1608910539
transform 1 0 7162 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1608910539
transform 1 0 8266 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1608910539
transform 1 0 9738 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_98
timestamp 1608910539
transform 1 0 9370 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 10106 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1608910539
transform 1 0 630 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 354 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1608910539
transform 1 0 1734 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1608910539
transform 1 0 3298 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1608910539
transform 1 0 2838 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 3206 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1608910539
transform 1 0 4402 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_63
timestamp 1608910539
transform 1 0 6150 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_56
timestamp 1608910539
transform 1 0 5506 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 6058 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_75
timestamp 1608910539
transform 1 0 7254 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_87
timestamp 1608910539
transform 1 0 8358 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_102
timestamp 1608910539
transform 1 0 9738 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_94
timestamp 1608910539
transform 1 0 9002 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 8910 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 10106 0 -1 11424
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4 0 60 800 6 x[0]
port 0 nsew signal tristate
rlabel metal2 s 1476 0 1532 800 6 x[1]
port 1 nsew signal tristate
rlabel metal2 s 2948 0 3004 800 6 x[2]
port 2 nsew signal tristate
rlabel metal2 s 4420 0 4476 800 6 x[3]
port 3 nsew signal tristate
rlabel metal2 s 5984 0 6040 800 6 x[4]
port 4 nsew signal tristate
rlabel metal2 s 7456 0 7512 800 6 x[5]
port 5 nsew signal tristate
rlabel metal2 s 8928 0 8984 800 6 x[6]
port 6 nsew signal tristate
rlabel metal2 s 10400 0 10456 800 6 x[7]
port 7 nsew signal tristate
rlabel metal4 s 8354 2128 8674 11472 6 VPWR
port 8 nsew power bidirectional
rlabel metal4 s 5090 2128 5410 11472 6 VPWR
port 9 nsew power bidirectional
rlabel metal4 s 1826 2128 2146 11472 6 VPWR
port 10 nsew power bidirectional
rlabel metal4 s 6722 2128 7042 11472 6 VGND
port 11 nsew ground bidirectional
rlabel metal4 s 3458 2128 3778 11472 6 VGND
port 12 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 10460 11472
<< end >>
