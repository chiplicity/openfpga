magic
tech EFS8A
magscale 1 2
timestamp 1602042237
<< locali >>
rect 16589 18207 16623 18377
rect 8493 17697 8654 17731
rect 8493 17527 8527 17697
rect 6779 14909 6906 14943
rect 2605 8993 2766 9027
rect 15243 8993 15370 9027
rect 2605 8823 2639 8993
rect 4479 7905 4514 7939
rect 14105 6817 14266 6851
rect 14105 6715 14139 6817
rect 11483 5049 11621 5083
<< viali >>
rect 14197 18377 14231 18411
rect 16589 18377 16623 18411
rect 16865 18377 16899 18411
rect 8769 18309 8803 18343
rect 7481 18241 7515 18275
rect 4604 18173 4638 18207
rect 4997 18173 5031 18207
rect 5800 18173 5834 18207
rect 6996 18173 7030 18207
rect 8284 18173 8318 18207
rect 9816 18173 9850 18207
rect 10241 18173 10275 18207
rect 13712 18173 13746 18207
rect 16380 18173 16414 18207
rect 16589 18173 16623 18207
rect 6193 18105 6227 18139
rect 4675 18037 4709 18071
rect 5871 18037 5905 18071
rect 7067 18037 7101 18071
rect 8355 18037 8389 18071
rect 9919 18037 9953 18071
rect 13783 18037 13817 18071
rect 16451 18037 16485 18071
rect 5641 17765 5675 17799
rect 1476 17697 1510 17731
rect 4144 17697 4178 17731
rect 10584 17697 10618 17731
rect 12332 17697 12366 17731
rect 13691 17697 13725 17731
rect 5917 17629 5951 17663
rect 7481 17629 7515 17663
rect 13783 17629 13817 17663
rect 15393 17629 15427 17663
rect 15945 17561 15979 17595
rect 1547 17493 1581 17527
rect 4215 17493 4249 17527
rect 8493 17493 8527 17527
rect 8723 17493 8757 17527
rect 10655 17493 10689 17527
rect 12403 17493 12437 17527
rect 1593 17289 1627 17323
rect 3985 17289 4019 17323
rect 5549 17289 5583 17323
rect 5825 17289 5859 17323
rect 9321 17289 9355 17323
rect 11345 17289 11379 17323
rect 12633 17289 12667 17323
rect 13001 17289 13035 17323
rect 14197 17289 14231 17323
rect 15761 17289 15795 17323
rect 1869 17153 1903 17187
rect 3617 17153 3651 17187
rect 4169 17153 4203 17187
rect 4813 17153 4847 17187
rect 8585 17153 8619 17187
rect 10149 17153 10183 17187
rect 10333 17153 10367 17187
rect 10609 17153 10643 17187
rect 13277 17153 13311 17187
rect 16037 17153 16071 17187
rect 16313 17153 16347 17187
rect 5641 17085 5675 17119
rect 6193 17085 6227 17119
rect 9137 17085 9171 17119
rect 9689 17085 9723 17119
rect 15000 17085 15034 17119
rect 2513 17017 2547 17051
rect 7389 17017 7423 17051
rect 8033 17017 8067 17051
rect 13921 17017 13955 17051
rect 15485 17017 15519 17051
rect 7113 16949 7147 16983
rect 15071 16949 15105 16983
rect 1869 16745 1903 16779
rect 16313 16745 16347 16779
rect 2513 16677 2547 16711
rect 4905 16677 4939 16711
rect 6009 16677 6043 16711
rect 8125 16677 8159 16711
rect 9781 16677 9815 16711
rect 10425 16677 10459 16711
rect 13737 16677 13771 16711
rect 1476 16609 1510 16643
rect 4261 16541 4295 16575
rect 6285 16541 6319 16575
rect 8401 16541 8435 16575
rect 14013 16541 14047 16575
rect 15393 16541 15427 16575
rect 16037 16541 16071 16575
rect 3065 16473 3099 16507
rect 1547 16405 1581 16439
rect 2237 16405 2271 16439
rect 6193 16201 6227 16235
rect 7665 16201 7699 16235
rect 8769 16201 8803 16235
rect 9505 16201 9539 16235
rect 13737 16201 13771 16235
rect 15025 16201 15059 16235
rect 2513 16065 2547 16099
rect 3065 16065 3099 16099
rect 4905 16065 4939 16099
rect 7849 16065 7883 16099
rect 8125 16065 8159 16099
rect 9689 16065 9723 16099
rect 9965 16065 9999 16099
rect 15485 16065 15519 16099
rect 15669 16065 15703 16099
rect 15945 16065 15979 16099
rect 2145 15929 2179 15963
rect 4261 15929 4295 15963
rect 1593 15861 1627 15895
rect 3617 15861 3651 15895
rect 4077 15861 4111 15895
rect 5733 15861 5767 15895
rect 9873 15657 9907 15691
rect 2237 15589 2271 15623
rect 2881 15589 2915 15623
rect 8125 15589 8159 15623
rect 15577 15589 15611 15623
rect 4997 15453 5031 15487
rect 6101 15453 6135 15487
rect 6745 15453 6779 15487
rect 15853 15453 15887 15487
rect 8677 15385 8711 15419
rect 2651 15113 2685 15147
rect 6101 15113 6135 15147
rect 6561 15113 6595 15147
rect 6975 15113 7009 15147
rect 7757 15113 7791 15147
rect 15393 15113 15427 15147
rect 7297 15045 7331 15079
rect 2145 14977 2179 15011
rect 8677 14977 8711 15011
rect 16313 14977 16347 15011
rect 1409 14909 1443 14943
rect 2580 14909 2614 14943
rect 3592 14909 3626 14943
rect 5708 14909 5742 14943
rect 6745 14909 6779 14943
rect 14841 14909 14875 14943
rect 14968 14909 15002 14943
rect 2973 14841 3007 14875
rect 4077 14841 4111 14875
rect 8125 14841 8159 14875
rect 8309 14841 8343 14875
rect 13921 14841 13955 14875
rect 15761 14841 15795 14875
rect 16037 14841 16071 14875
rect 1593 14773 1627 14807
rect 3663 14773 3697 14807
rect 5779 14773 5813 14807
rect 15071 14773 15105 14807
rect 7941 14569 7975 14603
rect 2421 14501 2455 14535
rect 4261 14501 4295 14535
rect 16037 14501 16071 14535
rect 5733 14433 5767 14467
rect 9724 14433 9758 14467
rect 2697 14365 2731 14399
rect 4537 14365 4571 14399
rect 16313 14365 16347 14399
rect 1685 14229 1719 14263
rect 5917 14229 5951 14263
rect 9827 14229 9861 14263
rect 2789 14025 2823 14059
rect 4813 14025 4847 14059
rect 5825 14025 5859 14059
rect 9321 14025 9355 14059
rect 9689 14025 9723 14059
rect 16037 14025 16071 14059
rect 16497 14025 16531 14059
rect 2329 13957 2363 13991
rect 1777 13889 1811 13923
rect 4537 13889 4571 13923
rect 5365 13889 5399 13923
rect 8677 13821 8711 13855
rect 16313 13821 16347 13855
rect 16865 13821 16899 13855
rect 3709 13753 3743 13787
rect 3893 13753 3927 13787
rect 8861 13685 8895 13719
rect 14657 13685 14691 13719
rect 1777 13481 1811 13515
rect 2053 13413 2087 13447
rect 15393 13413 15427 13447
rect 16037 13413 16071 13447
rect 4144 13345 4178 13379
rect 2329 13277 2363 13311
rect 4215 13141 4249 13175
rect 1547 12937 1581 12971
rect 2053 12937 2087 12971
rect 2329 12937 2363 12971
rect 3249 12937 3283 12971
rect 4169 12937 4203 12971
rect 15761 12937 15795 12971
rect 16129 12937 16163 12971
rect 3525 12869 3559 12903
rect 16497 12869 16531 12903
rect 4445 12801 4479 12835
rect 1476 12733 1510 12767
rect 3341 12733 3375 12767
rect 15352 12733 15386 12767
rect 15439 12733 15473 12767
rect 16313 12733 16347 12767
rect 16865 12733 16899 12767
rect 1685 12189 1719 12223
rect 2053 12189 2087 12223
rect 1547 11849 1581 11883
rect 2237 11849 2271 11883
rect 1476 11645 1510 11679
rect 1869 11645 1903 11679
rect 4144 11169 4178 11203
rect 16037 11101 16071 11135
rect 16313 11101 16347 11135
rect 4215 10965 4249 10999
rect 4629 10761 4663 10795
rect 16589 10761 16623 10795
rect 3433 10625 3467 10659
rect 3617 10625 3651 10659
rect 3893 10625 3927 10659
rect 15945 10625 15979 10659
rect 1869 10489 1903 10523
rect 2513 10489 2547 10523
rect 15669 10489 15703 10523
rect 1593 10421 1627 10455
rect 14565 10421 14599 10455
rect 15393 10421 15427 10455
rect 16451 10217 16485 10251
rect 1476 10081 1510 10115
rect 15368 10081 15402 10115
rect 16380 10081 16414 10115
rect 2513 10013 2547 10047
rect 2789 10013 2823 10047
rect 1547 9877 1581 9911
rect 1869 9877 1903 9911
rect 15439 9877 15473 9911
rect 1593 9673 1627 9707
rect 2053 9673 2087 9707
rect 7389 9673 7423 9707
rect 15393 9673 15427 9707
rect 16129 9673 16163 9707
rect 16497 9605 16531 9639
rect 2513 9537 2547 9571
rect 3801 9537 3835 9571
rect 1409 9469 1443 9503
rect 6904 9469 6938 9503
rect 16313 9469 16347 9503
rect 2973 9401 3007 9435
rect 3157 9401 3191 9435
rect 6975 9333 7009 9367
rect 16957 9333 16991 9367
rect 1593 9129 1627 9163
rect 2835 9129 2869 9163
rect 16497 9129 16531 9163
rect 6377 9061 6411 9095
rect 15209 8993 15243 9027
rect 15439 8993 15473 9027
rect 16313 8993 16347 9027
rect 6653 8925 6687 8959
rect 2605 8789 2639 8823
rect 6377 8585 6411 8619
rect 15301 8585 15335 8619
rect 16865 8585 16899 8619
rect 5917 8449 5951 8483
rect 16221 8449 16255 8483
rect 5273 8313 5307 8347
rect 14841 8313 14875 8347
rect 15669 8313 15703 8347
rect 15945 8313 15979 8347
rect 2789 8245 2823 8279
rect 4997 8245 5031 8279
rect 4583 8041 4617 8075
rect 6377 7973 6411 8007
rect 4445 7905 4479 7939
rect 14264 7905 14298 7939
rect 7021 7837 7055 7871
rect 16037 7837 16071 7871
rect 16405 7837 16439 7871
rect 14335 7701 14369 7735
rect 4445 7497 4479 7531
rect 6377 7497 6411 7531
rect 14473 7497 14507 7531
rect 14841 7497 14875 7531
rect 15485 7497 15519 7531
rect 16313 7361 16347 7395
rect 16957 7361 16991 7395
rect 13972 7293 14006 7327
rect 14984 7293 15018 7327
rect 14059 7225 14093 7259
rect 15071 7225 15105 7259
rect 15761 7225 15795 7259
rect 16037 7225 16071 7259
rect 6837 7157 6871 7191
rect 6377 6885 6411 6919
rect 7021 6885 7055 6919
rect 7884 6817 7918 6851
rect 12700 6817 12734 6851
rect 15945 6749 15979 6783
rect 16313 6749 16347 6783
rect 14105 6681 14139 6715
rect 7987 6613 8021 6647
rect 12771 6613 12805 6647
rect 14335 6613 14369 6647
rect 6377 6409 6411 6443
rect 7481 6409 7515 6443
rect 7849 6409 7883 6443
rect 15807 6409 15841 6443
rect 16497 6409 16531 6443
rect 15209 6341 15243 6375
rect 13185 6273 13219 6307
rect 6837 6205 6871 6239
rect 12700 6205 12734 6239
rect 13712 6205 13746 6239
rect 14724 6205 14758 6239
rect 15736 6205 15770 6239
rect 14565 6137 14599 6171
rect 7021 6069 7055 6103
rect 12771 6069 12805 6103
rect 13461 6069 13495 6103
rect 13783 6069 13817 6103
rect 14197 6069 14231 6103
rect 14795 6069 14829 6103
rect 16221 6069 16255 6103
rect 15393 5797 15427 5831
rect 12541 5661 12575 5695
rect 14105 5661 14139 5695
rect 15669 5661 15703 5695
rect 15761 5321 15795 5355
rect 15393 5253 15427 5287
rect 11897 5185 11931 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 9940 5117 9974 5151
rect 11412 5117 11446 5151
rect 11621 5049 11655 5083
rect 13461 5049 13495 5083
rect 13645 5049 13679 5083
rect 14289 5049 14323 5083
rect 10011 4981 10045 5015
rect 10425 4981 10459 5015
rect 12541 4981 12575 5015
rect 10103 4777 10137 4811
rect 12357 4777 12391 4811
rect 13737 4709 13771 4743
rect 14381 4709 14415 4743
rect 10032 4641 10066 4675
rect 11044 4641 11078 4675
rect 12173 4641 12207 4675
rect 15577 4573 15611 4607
rect 15853 4573 15887 4607
rect 11115 4437 11149 4471
rect 1869 4233 1903 4267
rect 12173 4233 12207 4267
rect 12633 4233 12667 4267
rect 13921 4233 13955 4267
rect 16037 4233 16071 4267
rect 14841 4165 14875 4199
rect 10149 4097 10183 4131
rect 12909 4097 12943 4131
rect 15117 4097 15151 4131
rect 15761 4097 15795 4131
rect 1476 4029 1510 4063
rect 5400 4029 5434 4063
rect 5825 4029 5859 4063
rect 9264 4029 9298 4063
rect 9689 4029 9723 4063
rect 11412 4029 11446 4063
rect 13553 3961 13587 3995
rect 1547 3893 1581 3927
rect 5503 3893 5537 3927
rect 7021 3893 7055 3927
rect 9367 3893 9401 3927
rect 10333 3893 10367 3927
rect 11069 3893 11103 3927
rect 11483 3893 11517 3927
rect 11897 3893 11931 3927
rect 2145 3621 2179 3655
rect 6285 3621 6319 3655
rect 10149 3621 10183 3655
rect 15393 3621 15427 3655
rect 7757 3553 7791 3587
rect 13829 3553 13863 3587
rect 2789 3485 2823 3519
rect 4169 3485 4203 3519
rect 4813 3485 4847 3519
rect 6929 3485 6963 3519
rect 10793 3485 10827 3519
rect 11713 3485 11747 3519
rect 12357 3485 12391 3519
rect 15669 3485 15703 3519
rect 7941 3349 7975 3383
rect 14013 3349 14047 3383
rect 2145 3145 2179 3179
rect 6285 3145 6319 3179
rect 10241 3145 10275 3179
rect 12173 3145 12207 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 15485 3145 15519 3179
rect 3985 3077 4019 3111
rect 9873 3077 9907 3111
rect 11437 3077 11471 3111
rect 11805 3077 11839 3111
rect 2329 3009 2363 3043
rect 4353 3009 4387 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 9137 3009 9171 3043
rect 9321 3009 9355 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 12817 3009 12851 3043
rect 14473 3009 14507 3043
rect 14749 3009 14783 3043
rect 15853 3009 15887 3043
rect 16037 3009 16071 3043
rect 4940 2941 4974 2975
rect 5365 2941 5399 2975
rect 3433 2873 3467 2907
rect 5043 2873 5077 2907
rect 8033 2873 8067 2907
rect 12541 2873 12575 2907
rect 16681 2873 16715 2907
rect 3157 2805 3191 2839
rect 8309 2805 8343 2839
rect 2007 2601 2041 2635
rect 3525 2601 3559 2635
rect 3801 2601 3835 2635
rect 5963 2601 5997 2635
rect 7113 2601 7147 2635
rect 10517 2601 10551 2635
rect 12449 2601 12483 2635
rect 15761 2601 15795 2635
rect 4169 2533 4203 2567
rect 4813 2533 4847 2567
rect 7389 2533 7423 2567
rect 8033 2533 8067 2567
rect 10977 2533 11011 2567
rect 13001 2533 13035 2567
rect 13645 2533 13679 2567
rect 16037 2533 16071 2567
rect 1936 2465 1970 2499
rect 2881 2465 2915 2499
rect 5892 2465 5926 2499
rect 10333 2465 10367 2499
rect 11437 2465 11471 2499
rect 11989 2465 12023 2499
rect 6377 2397 6411 2431
rect 16313 2397 16347 2431
rect 3065 2329 3099 2363
rect 11621 2329 11655 2363
rect 2421 2261 2455 2295
<< metal1 >>
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 13170 20584 13176 20596
rect 12492 20556 13176 20584
rect 12492 20544 12498 20556
rect 13170 20544 13176 20556
rect 13228 20544 13234 20596
rect 1104 18522 17756 18544
rect 1104 18470 4135 18522
rect 4187 18470 4199 18522
rect 4251 18470 4263 18522
rect 4315 18470 4327 18522
rect 4379 18470 10441 18522
rect 10493 18470 10505 18522
rect 10557 18470 10569 18522
rect 10621 18470 10633 18522
rect 10685 18470 16748 18522
rect 16800 18470 16812 18522
rect 16864 18470 16876 18522
rect 16928 18470 16940 18522
rect 16992 18470 17756 18522
rect 1104 18448 17756 18470
rect 14182 18408 14188 18420
rect 14143 18380 14188 18408
rect 14182 18368 14188 18380
rect 14240 18368 14246 18420
rect 16577 18411 16635 18417
rect 16577 18377 16589 18411
rect 16623 18408 16635 18411
rect 16853 18411 16911 18417
rect 16853 18408 16865 18411
rect 16623 18380 16865 18408
rect 16623 18377 16635 18380
rect 16577 18371 16635 18377
rect 16853 18377 16865 18380
rect 16899 18408 16911 18411
rect 18230 18408 18236 18420
rect 16899 18380 18236 18408
rect 16899 18377 16911 18380
rect 16853 18371 16911 18377
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 8757 18343 8815 18349
rect 8757 18309 8769 18343
rect 8803 18340 8815 18343
rect 18414 18340 18420 18352
rect 8803 18312 18420 18340
rect 8803 18309 8815 18312
rect 8757 18303 8815 18309
rect 7466 18272 7472 18284
rect 6999 18244 7472 18272
rect 4592 18207 4650 18213
rect 4592 18173 4604 18207
rect 4638 18204 4650 18207
rect 4890 18204 4896 18216
rect 4638 18176 4896 18204
rect 4638 18173 4650 18176
rect 4592 18167 4650 18173
rect 4890 18164 4896 18176
rect 4948 18204 4954 18216
rect 6999 18213 7027 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 4985 18207 5043 18213
rect 4985 18204 4997 18207
rect 4948 18176 4997 18204
rect 4948 18164 4954 18176
rect 4985 18173 4997 18176
rect 5031 18173 5043 18207
rect 4985 18167 5043 18173
rect 5788 18207 5846 18213
rect 5788 18173 5800 18207
rect 5834 18204 5846 18207
rect 6984 18207 7042 18213
rect 5834 18176 6224 18204
rect 5834 18173 5846 18176
rect 5788 18167 5846 18173
rect 6196 18145 6224 18176
rect 6984 18173 6996 18207
rect 7030 18173 7042 18207
rect 6984 18167 7042 18173
rect 8272 18207 8330 18213
rect 8272 18173 8284 18207
rect 8318 18204 8330 18207
rect 8772 18204 8800 18303
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 17034 18272 17040 18284
rect 8318 18176 8800 18204
rect 8864 18244 17040 18272
rect 8318 18173 8330 18176
rect 8272 18167 8330 18173
rect 6181 18139 6239 18145
rect 6181 18105 6193 18139
rect 6227 18136 6239 18139
rect 8864 18136 8892 18244
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 9398 18164 9404 18216
rect 9456 18204 9462 18216
rect 9804 18207 9862 18213
rect 9804 18204 9816 18207
rect 9456 18176 9816 18204
rect 9456 18164 9462 18176
rect 9804 18173 9816 18176
rect 9850 18204 9862 18207
rect 10229 18207 10287 18213
rect 10229 18204 10241 18207
rect 9850 18176 10241 18204
rect 9850 18173 9862 18176
rect 9804 18167 9862 18173
rect 10229 18173 10241 18176
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 13700 18207 13758 18213
rect 13700 18173 13712 18207
rect 13746 18204 13758 18207
rect 14182 18204 14188 18216
rect 13746 18176 14188 18204
rect 13746 18173 13758 18176
rect 13700 18167 13758 18173
rect 14182 18164 14188 18176
rect 14240 18164 14246 18216
rect 16368 18207 16426 18213
rect 16368 18173 16380 18207
rect 16414 18204 16426 18207
rect 16577 18207 16635 18213
rect 16577 18204 16589 18207
rect 16414 18176 16589 18204
rect 16414 18173 16426 18176
rect 16368 18167 16426 18173
rect 16577 18173 16589 18176
rect 16623 18173 16635 18207
rect 16577 18167 16635 18173
rect 6227 18108 8892 18136
rect 6227 18105 6239 18108
rect 6181 18099 6239 18105
rect 8938 18096 8944 18148
rect 8996 18136 9002 18148
rect 18506 18136 18512 18148
rect 8996 18108 18512 18136
rect 8996 18096 9002 18108
rect 18506 18096 18512 18108
rect 18564 18096 18570 18148
rect 4663 18071 4721 18077
rect 4663 18037 4675 18071
rect 4709 18068 4721 18071
rect 5534 18068 5540 18080
rect 4709 18040 5540 18068
rect 4709 18037 4721 18040
rect 4663 18031 4721 18037
rect 5534 18028 5540 18040
rect 5592 18028 5598 18080
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 5859 18071 5917 18077
rect 5859 18068 5871 18071
rect 5684 18040 5871 18068
rect 5684 18028 5690 18040
rect 5859 18037 5871 18040
rect 5905 18037 5917 18071
rect 5859 18031 5917 18037
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 7055 18071 7113 18077
rect 7055 18068 7067 18071
rect 6328 18040 7067 18068
rect 6328 18028 6334 18040
rect 7055 18037 7067 18040
rect 7101 18037 7113 18071
rect 7055 18031 7113 18037
rect 8110 18028 8116 18080
rect 8168 18068 8174 18080
rect 8343 18071 8401 18077
rect 8343 18068 8355 18071
rect 8168 18040 8355 18068
rect 8168 18028 8174 18040
rect 8343 18037 8355 18040
rect 8389 18037 8401 18071
rect 8343 18031 8401 18037
rect 9766 18028 9772 18080
rect 9824 18068 9830 18080
rect 9907 18071 9965 18077
rect 9907 18068 9919 18071
rect 9824 18040 9919 18068
rect 9824 18028 9830 18040
rect 9907 18037 9919 18040
rect 9953 18037 9965 18071
rect 9907 18031 9965 18037
rect 13771 18071 13829 18077
rect 13771 18037 13783 18071
rect 13817 18068 13829 18071
rect 13906 18068 13912 18080
rect 13817 18040 13912 18068
rect 13817 18037 13829 18040
rect 13771 18031 13829 18037
rect 13906 18028 13912 18040
rect 13964 18028 13970 18080
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16439 18071 16497 18077
rect 16439 18068 16451 18071
rect 16080 18040 16451 18068
rect 16080 18028 16086 18040
rect 16439 18037 16451 18040
rect 16485 18037 16497 18071
rect 16439 18031 16497 18037
rect 1104 17978 17756 18000
rect 1104 17926 7288 17978
rect 7340 17926 7352 17978
rect 7404 17926 7416 17978
rect 7468 17926 7480 17978
rect 7532 17926 13595 17978
rect 13647 17926 13659 17978
rect 13711 17926 13723 17978
rect 13775 17926 13787 17978
rect 13839 17926 17756 17978
rect 1104 17904 17756 17926
rect 1210 17756 1216 17808
rect 1268 17796 1274 17808
rect 5626 17796 5632 17808
rect 1268 17768 1507 17796
rect 5587 17768 5632 17796
rect 1268 17756 1274 17768
rect 1479 17737 1507 17768
rect 5626 17756 5632 17768
rect 5684 17756 5690 17808
rect 8386 17756 8392 17808
rect 8444 17796 8450 17808
rect 8444 17768 12756 17796
rect 8444 17756 8450 17768
rect 1464 17731 1522 17737
rect 1464 17697 1476 17731
rect 1510 17697 1522 17731
rect 1464 17691 1522 17697
rect 4132 17731 4190 17737
rect 4132 17697 4144 17731
rect 4178 17728 4190 17731
rect 4430 17728 4436 17740
rect 4178 17700 4436 17728
rect 4178 17697 4190 17700
rect 4132 17691 4190 17697
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 10572 17731 10630 17737
rect 10572 17697 10584 17731
rect 10618 17728 10630 17731
rect 11882 17728 11888 17740
rect 10618 17700 11888 17728
rect 10618 17697 10630 17700
rect 10572 17691 10630 17697
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12320 17731 12378 17737
rect 12320 17697 12332 17731
rect 12366 17728 12378 17731
rect 12618 17728 12624 17740
rect 12366 17700 12624 17728
rect 12366 17697 12378 17700
rect 12320 17691 12378 17697
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 12728 17728 12756 17768
rect 13679 17731 13737 17737
rect 13679 17728 13691 17731
rect 12728 17700 13691 17728
rect 13679 17697 13691 17700
rect 13725 17728 13737 17731
rect 14182 17728 14188 17740
rect 13725 17700 14188 17728
rect 13725 17697 13737 17700
rect 13679 17691 13737 17697
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 5905 17663 5963 17669
rect 5905 17660 5917 17663
rect 4856 17632 5917 17660
rect 4856 17620 4862 17632
rect 5905 17629 5917 17632
rect 5951 17629 5963 17663
rect 5905 17623 5963 17629
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17660 7527 17663
rect 7650 17660 7656 17672
rect 7515 17632 7656 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 13771 17663 13829 17669
rect 13771 17629 13783 17663
rect 13817 17660 13829 17663
rect 15381 17663 15439 17669
rect 15381 17660 15393 17663
rect 13817 17632 15393 17660
rect 13817 17629 13829 17632
rect 13771 17623 13829 17629
rect 15381 17629 15393 17632
rect 15427 17660 15439 17663
rect 15746 17660 15752 17672
rect 15427 17632 15752 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 15654 17552 15660 17604
rect 15712 17592 15718 17604
rect 15933 17595 15991 17601
rect 15933 17592 15945 17595
rect 15712 17564 15945 17592
rect 15712 17552 15718 17564
rect 15933 17561 15945 17564
rect 15979 17561 15991 17595
rect 15933 17555 15991 17561
rect 1535 17527 1593 17533
rect 1535 17493 1547 17527
rect 1581 17524 1593 17527
rect 1854 17524 1860 17536
rect 1581 17496 1860 17524
rect 1581 17493 1593 17496
rect 1535 17487 1593 17493
rect 1854 17484 1860 17496
rect 1912 17484 1918 17536
rect 3970 17484 3976 17536
rect 4028 17524 4034 17536
rect 4203 17527 4261 17533
rect 4203 17524 4215 17527
rect 4028 17496 4215 17524
rect 4028 17484 4034 17496
rect 4203 17493 4215 17496
rect 4249 17493 4261 17527
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 4203 17487 4261 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8711 17527 8769 17533
rect 8711 17493 8723 17527
rect 8757 17524 8769 17527
rect 9122 17524 9128 17536
rect 8757 17496 9128 17524
rect 8757 17493 8769 17496
rect 8711 17487 8769 17493
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 10643 17527 10701 17533
rect 10643 17524 10655 17527
rect 10376 17496 10655 17524
rect 10376 17484 10382 17496
rect 10643 17493 10655 17496
rect 10689 17493 10701 17527
rect 10643 17487 10701 17493
rect 12391 17527 12449 17533
rect 12391 17493 12403 17527
rect 12437 17524 12449 17527
rect 12986 17524 12992 17536
rect 12437 17496 12992 17524
rect 12437 17493 12449 17496
rect 12391 17487 12449 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 1104 17434 17756 17456
rect 1104 17382 4135 17434
rect 4187 17382 4199 17434
rect 4251 17382 4263 17434
rect 4315 17382 4327 17434
rect 4379 17382 10441 17434
rect 10493 17382 10505 17434
rect 10557 17382 10569 17434
rect 10621 17382 10633 17434
rect 10685 17382 16748 17434
rect 16800 17382 16812 17434
rect 16864 17382 16876 17434
rect 16928 17382 16940 17434
rect 16992 17382 17756 17434
rect 1104 17360 17756 17382
rect 1210 17280 1216 17332
rect 1268 17320 1274 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1268 17292 1593 17320
rect 1268 17280 1274 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 1581 17283 1639 17289
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4430 17320 4436 17332
rect 4019 17292 4436 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 5537 17323 5595 17329
rect 5537 17289 5549 17323
rect 5583 17320 5595 17323
rect 5626 17320 5632 17332
rect 5583 17292 5632 17320
rect 5583 17289 5595 17292
rect 5537 17283 5595 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5810 17320 5816 17332
rect 5771 17292 5816 17320
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 9309 17323 9367 17329
rect 9309 17289 9321 17323
rect 9355 17320 9367 17323
rect 10226 17320 10232 17332
rect 9355 17292 10232 17320
rect 9355 17289 9367 17292
rect 9309 17283 9367 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11882 17320 11888 17332
rect 11379 17292 11888 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 12618 17320 12624 17332
rect 12579 17292 12624 17320
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 12986 17320 12992 17332
rect 12947 17292 12992 17320
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 14182 17320 14188 17332
rect 14143 17292 14188 17320
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 15746 17320 15752 17332
rect 15707 17292 15752 17320
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 1854 17184 1860 17196
rect 1815 17156 1860 17184
rect 1854 17144 1860 17156
rect 1912 17144 1918 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 3970 17184 3976 17196
rect 3651 17156 3976 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 3970 17144 3976 17156
rect 4028 17184 4034 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 4028 17156 4169 17184
rect 4028 17144 4034 17156
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 4798 17184 4804 17196
rect 4759 17156 4804 17184
rect 4157 17147 4215 17153
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8478 17184 8484 17196
rect 8076 17156 8484 17184
rect 8076 17144 8082 17156
rect 8478 17144 8484 17156
rect 8536 17184 8542 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 8536 17156 8585 17184
rect 8536 17144 8542 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10318 17184 10324 17196
rect 10183 17156 10324 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 10594 17184 10600 17196
rect 10555 17156 10600 17184
rect 10594 17144 10600 17156
rect 10652 17144 10658 17196
rect 13004 17184 13032 17280
rect 13265 17187 13323 17193
rect 13265 17184 13277 17187
rect 13004 17156 13277 17184
rect 13265 17153 13277 17156
rect 13311 17153 13323 17187
rect 16022 17184 16028 17196
rect 15983 17156 16028 17184
rect 13265 17147 13323 17153
rect 16022 17144 16028 17156
rect 16080 17144 16086 17196
rect 16114 17144 16120 17196
rect 16172 17184 16178 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 16172 17156 16313 17184
rect 16172 17144 16178 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5592 17088 5641 17116
rect 5592 17076 5598 17088
rect 5629 17085 5641 17088
rect 5675 17116 5687 17119
rect 6181 17119 6239 17125
rect 6181 17116 6193 17119
rect 5675 17088 6193 17116
rect 5675 17085 5687 17088
rect 5629 17079 5687 17085
rect 6181 17085 6193 17088
rect 6227 17085 6239 17119
rect 9122 17116 9128 17128
rect 9083 17088 9128 17116
rect 6181 17079 6239 17085
rect 9122 17076 9128 17088
rect 9180 17116 9186 17128
rect 9677 17119 9735 17125
rect 9677 17116 9689 17119
rect 9180 17088 9689 17116
rect 9180 17076 9186 17088
rect 9677 17085 9689 17088
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 14988 17119 15046 17125
rect 14988 17085 15000 17119
rect 15034 17085 15046 17119
rect 14988 17079 15046 17085
rect 2498 17048 2504 17060
rect 2459 17020 2504 17048
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 7377 17051 7435 17057
rect 7377 17048 7389 17051
rect 7116 17020 7389 17048
rect 7116 16992 7144 17020
rect 7377 17017 7389 17020
rect 7423 17017 7435 17051
rect 7377 17011 7435 17017
rect 8021 17051 8079 17057
rect 8021 17017 8033 17051
rect 8067 17048 8079 17051
rect 8386 17048 8392 17060
rect 8067 17020 8392 17048
rect 8067 17017 8079 17020
rect 8021 17011 8079 17017
rect 8386 17008 8392 17020
rect 8444 17008 8450 17060
rect 13909 17051 13967 17057
rect 13909 17017 13921 17051
rect 13955 17048 13967 17051
rect 13998 17048 14004 17060
rect 13955 17020 14004 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 15003 17048 15031 17079
rect 15470 17048 15476 17060
rect 15003 17020 15476 17048
rect 15470 17008 15476 17020
rect 15528 17008 15534 17060
rect 7098 16980 7104 16992
rect 7059 16952 7104 16980
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 15059 16983 15117 16989
rect 15059 16949 15071 16983
rect 15105 16980 15117 16983
rect 15286 16980 15292 16992
rect 15105 16952 15292 16980
rect 15105 16949 15117 16952
rect 15059 16943 15117 16949
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 1104 16890 17756 16912
rect 1104 16838 7288 16890
rect 7340 16838 7352 16890
rect 7404 16838 7416 16890
rect 7468 16838 7480 16890
rect 7532 16838 13595 16890
rect 13647 16838 13659 16890
rect 13711 16838 13723 16890
rect 13775 16838 13787 16890
rect 13839 16838 17756 16890
rect 1104 16816 17756 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16301 16779 16359 16785
rect 16301 16776 16313 16779
rect 16080 16748 16313 16776
rect 16080 16736 16086 16748
rect 16301 16745 16313 16748
rect 16347 16745 16359 16779
rect 16301 16739 16359 16745
rect 2498 16708 2504 16720
rect 2459 16680 2504 16708
rect 2498 16668 2504 16680
rect 2556 16668 2562 16720
rect 4890 16708 4896 16720
rect 4851 16680 4896 16708
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 5997 16711 6055 16717
rect 5997 16677 6009 16711
rect 6043 16708 6055 16711
rect 6270 16708 6276 16720
rect 6043 16680 6276 16708
rect 6043 16677 6055 16680
rect 5997 16671 6055 16677
rect 6270 16668 6276 16680
rect 6328 16668 6334 16720
rect 8110 16708 8116 16720
rect 8071 16680 8116 16708
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 9766 16708 9772 16720
rect 9727 16680 9772 16708
rect 9766 16668 9772 16680
rect 9824 16668 9830 16720
rect 9858 16668 9864 16720
rect 9916 16708 9922 16720
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 9916 16680 10425 16708
rect 9916 16668 9922 16680
rect 10413 16677 10425 16680
rect 10459 16708 10471 16711
rect 10594 16708 10600 16720
rect 10459 16680 10600 16708
rect 10459 16677 10471 16680
rect 10413 16671 10471 16677
rect 10594 16668 10600 16680
rect 10652 16668 10658 16720
rect 13725 16711 13783 16717
rect 13725 16677 13737 16711
rect 13771 16708 13783 16711
rect 13906 16708 13912 16720
rect 13771 16680 13912 16708
rect 13771 16677 13783 16680
rect 13725 16671 13783 16677
rect 13906 16668 13912 16680
rect 13964 16668 13970 16720
rect 1464 16643 1522 16649
rect 1464 16609 1476 16643
rect 1510 16640 1522 16643
rect 1578 16640 1584 16652
rect 1510 16612 1584 16640
rect 1510 16609 1522 16612
rect 1464 16603 1522 16609
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 4430 16572 4436 16584
rect 4295 16544 4436 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 8386 16572 8392 16584
rect 8347 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 13998 16572 14004 16584
rect 13959 16544 14004 16572
rect 13998 16532 14004 16544
rect 14056 16572 14062 16584
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 14056 16544 15393 16572
rect 14056 16532 14062 16544
rect 15381 16541 15393 16544
rect 15427 16541 15439 16575
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 15381 16535 15439 16541
rect 16022 16532 16028 16544
rect 16080 16532 16086 16584
rect 3053 16507 3111 16513
rect 3053 16473 3065 16507
rect 3099 16504 3111 16507
rect 8018 16504 8024 16516
rect 3099 16476 8024 16504
rect 3099 16473 3111 16476
rect 3053 16467 3111 16473
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 1535 16439 1593 16445
rect 1535 16405 1547 16439
rect 1581 16436 1593 16439
rect 2038 16436 2044 16448
rect 1581 16408 2044 16436
rect 1581 16405 1593 16408
rect 1535 16399 1593 16405
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 2130 16396 2136 16448
rect 2188 16436 2194 16448
rect 2225 16439 2283 16445
rect 2225 16436 2237 16439
rect 2188 16408 2237 16436
rect 2188 16396 2194 16408
rect 2225 16405 2237 16408
rect 2271 16405 2283 16439
rect 2225 16399 2283 16405
rect 1104 16346 17756 16368
rect 1104 16294 4135 16346
rect 4187 16294 4199 16346
rect 4251 16294 4263 16346
rect 4315 16294 4327 16346
rect 4379 16294 10441 16346
rect 10493 16294 10505 16346
rect 10557 16294 10569 16346
rect 10621 16294 10633 16346
rect 10685 16294 16748 16346
rect 16800 16294 16812 16346
rect 16864 16294 16876 16346
rect 16928 16294 16940 16346
rect 16992 16294 17756 16346
rect 1104 16272 17756 16294
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 7650 16232 7656 16244
rect 7611 16204 7656 16232
rect 7650 16192 7656 16204
rect 7708 16232 7714 16244
rect 7708 16204 7880 16232
rect 7708 16192 7714 16204
rect 2498 16096 2504 16108
rect 2459 16068 2504 16096
rect 2498 16056 2504 16068
rect 2556 16096 2562 16108
rect 3053 16099 3111 16105
rect 3053 16096 3065 16099
rect 2556 16068 3065 16096
rect 2556 16056 2562 16068
rect 3053 16065 3065 16068
rect 3099 16065 3111 16099
rect 3053 16059 3111 16065
rect 3602 16056 3608 16108
rect 3660 16096 3666 16108
rect 4246 16096 4252 16108
rect 3660 16068 4252 16096
rect 3660 16056 3666 16068
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 4890 16096 4896 16108
rect 4851 16068 4896 16096
rect 4890 16056 4896 16068
rect 4948 16056 4954 16108
rect 7852 16105 7880 16204
rect 8110 16192 8116 16244
rect 8168 16232 8174 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8168 16204 8769 16232
rect 8168 16192 8174 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 9766 16232 9772 16244
rect 9539 16204 9772 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 13725 16235 13783 16241
rect 13725 16201 13737 16235
rect 13771 16232 13783 16235
rect 13906 16232 13912 16244
rect 13771 16204 13912 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 13998 16192 14004 16244
rect 14056 16232 14062 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14056 16204 15025 16232
rect 14056 16192 14062 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16065 7895 16099
rect 7837 16059 7895 16065
rect 8018 16056 8024 16108
rect 8076 16096 8082 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 8076 16068 8125 16096
rect 8076 16056 8082 16068
rect 8113 16065 8125 16068
rect 8159 16065 8171 16099
rect 8113 16059 8171 16065
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9858 16096 9864 16108
rect 9723 16068 9864 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 9950 16056 9956 16108
rect 10008 16096 10014 16108
rect 15473 16099 15531 16105
rect 10008 16068 10053 16096
rect 10008 16056 10014 16068
rect 15473 16065 15485 16099
rect 15519 16096 15531 16099
rect 15654 16096 15660 16108
rect 15519 16068 15660 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15654 16056 15660 16068
rect 15712 16056 15718 16108
rect 15930 16096 15936 16108
rect 15891 16068 15936 16096
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 2130 15960 2136 15972
rect 2091 15932 2136 15960
rect 2130 15920 2136 15932
rect 2188 15920 2194 15972
rect 4246 15960 4252 15972
rect 4159 15932 4252 15960
rect 4246 15920 4252 15932
rect 4304 15960 4310 15972
rect 6270 15960 6276 15972
rect 4304 15932 6276 15960
rect 4304 15920 4310 15932
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 3602 15892 3608 15904
rect 3563 15864 3608 15892
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 4065 15895 4123 15901
rect 4065 15861 4077 15895
rect 4111 15892 4123 15895
rect 4430 15892 4436 15904
rect 4111 15864 4436 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 4430 15852 4436 15864
rect 4488 15892 4494 15904
rect 5721 15895 5779 15901
rect 5721 15892 5733 15895
rect 4488 15864 5733 15892
rect 4488 15852 4494 15864
rect 5721 15861 5733 15864
rect 5767 15861 5779 15895
rect 5721 15855 5779 15861
rect 1104 15802 17756 15824
rect 1104 15750 7288 15802
rect 7340 15750 7352 15802
rect 7404 15750 7416 15802
rect 7468 15750 7480 15802
rect 7532 15750 13595 15802
rect 13647 15750 13659 15802
rect 13711 15750 13723 15802
rect 13775 15750 13787 15802
rect 13839 15750 17756 15802
rect 1104 15728 17756 15750
rect 9858 15688 9864 15700
rect 9819 15660 9864 15688
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 2038 15580 2044 15632
rect 2096 15620 2102 15632
rect 2225 15623 2283 15629
rect 2225 15620 2237 15623
rect 2096 15592 2237 15620
rect 2096 15580 2102 15592
rect 2225 15589 2237 15592
rect 2271 15589 2283 15623
rect 2225 15583 2283 15589
rect 2869 15623 2927 15629
rect 2869 15589 2881 15623
rect 2915 15620 2927 15623
rect 3602 15620 3608 15632
rect 2915 15592 3608 15620
rect 2915 15589 2927 15592
rect 2869 15583 2927 15589
rect 3602 15580 3608 15592
rect 3660 15580 3666 15632
rect 8113 15623 8171 15629
rect 8113 15589 8125 15623
rect 8159 15620 8171 15623
rect 8386 15620 8392 15632
rect 8159 15592 8392 15620
rect 8159 15589 8171 15592
rect 8113 15583 8171 15589
rect 8386 15580 8392 15592
rect 8444 15580 8450 15632
rect 15286 15580 15292 15632
rect 15344 15620 15350 15632
rect 15565 15623 15623 15629
rect 15565 15620 15577 15623
rect 15344 15592 15577 15620
rect 15344 15580 15350 15592
rect 15565 15589 15577 15592
rect 15611 15589 15623 15623
rect 15565 15583 15623 15589
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 6086 15484 6092 15496
rect 5031 15456 6092 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 6546 15444 6552 15496
rect 6604 15484 6610 15496
rect 6733 15487 6791 15493
rect 6733 15484 6745 15487
rect 6604 15456 6745 15484
rect 6604 15444 6610 15456
rect 6733 15453 6745 15456
rect 6779 15484 6791 15487
rect 9950 15484 9956 15496
rect 6779 15456 9956 15484
rect 6779 15453 6791 15456
rect 6733 15447 6791 15453
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15712 15456 15853 15484
rect 15712 15444 15718 15456
rect 15841 15453 15853 15456
rect 15887 15453 15899 15487
rect 15841 15447 15899 15453
rect 8662 15416 8668 15428
rect 8623 15388 8668 15416
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 1104 15258 17756 15280
rect 1104 15206 4135 15258
rect 4187 15206 4199 15258
rect 4251 15206 4263 15258
rect 4315 15206 4327 15258
rect 4379 15206 10441 15258
rect 10493 15206 10505 15258
rect 10557 15206 10569 15258
rect 10621 15206 10633 15258
rect 10685 15206 16748 15258
rect 16800 15206 16812 15258
rect 16864 15206 16876 15258
rect 16928 15206 16940 15258
rect 16992 15206 17756 15258
rect 1104 15184 17756 15206
rect 2130 15104 2136 15156
rect 2188 15144 2194 15156
rect 2639 15147 2697 15153
rect 2639 15144 2651 15147
rect 2188 15116 2651 15144
rect 2188 15104 2194 15116
rect 2639 15113 2651 15116
rect 2685 15113 2697 15147
rect 6086 15144 6092 15156
rect 6047 15116 6092 15144
rect 2639 15107 2697 15113
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 6546 15144 6552 15156
rect 6507 15116 6552 15144
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6963 15147 7021 15153
rect 6963 15113 6975 15147
rect 7009 15144 7021 15147
rect 7098 15144 7104 15156
rect 7009 15116 7104 15144
rect 7009 15113 7021 15116
rect 6963 15107 7021 15113
rect 7098 15104 7104 15116
rect 7156 15104 7162 15156
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 8386 15144 8392 15156
rect 7791 15116 8392 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 15381 15147 15439 15153
rect 15381 15144 15393 15147
rect 15344 15116 15393 15144
rect 15344 15104 15350 15116
rect 15381 15113 15393 15116
rect 15427 15113 15439 15147
rect 15381 15107 15439 15113
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7285 15079 7343 15085
rect 7285 15076 7297 15079
rect 6880 15048 7297 15076
rect 6880 15036 6886 15048
rect 7285 15045 7297 15048
rect 7331 15045 7343 15079
rect 7285 15039 7343 15045
rect 2038 14968 2044 15020
rect 2096 15008 2102 15020
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 2096 14980 2145 15008
rect 2096 14968 2102 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1670 14940 1676 14952
rect 1443 14912 1676 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 1670 14900 1676 14912
rect 1728 14900 1734 14952
rect 2568 14943 2626 14949
rect 2568 14909 2580 14943
rect 2614 14909 2626 14943
rect 2568 14903 2626 14909
rect 3580 14943 3638 14949
rect 3580 14909 3592 14943
rect 3626 14940 3638 14943
rect 5696 14943 5754 14949
rect 3626 14912 4108 14940
rect 3626 14909 3638 14912
rect 3580 14903 3638 14909
rect 1486 14832 1492 14884
rect 1544 14872 1550 14884
rect 2583 14872 2611 14903
rect 4080 14881 4108 14912
rect 5696 14909 5708 14943
rect 5742 14940 5754 14943
rect 6546 14940 6552 14952
rect 5742 14912 6552 14940
rect 5742 14909 5754 14912
rect 5696 14903 5754 14909
rect 6546 14900 6552 14912
rect 6604 14900 6610 14952
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14940 6791 14943
rect 6840 14940 6868 15036
rect 8662 15008 8668 15020
rect 8623 14980 8668 15008
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 16298 15008 16304 15020
rect 14971 14980 16304 15008
rect 14971 14949 14999 14980
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 6779 14912 6868 14940
rect 14829 14943 14887 14949
rect 6779 14909 6791 14912
rect 6733 14903 6791 14909
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 14956 14943 15014 14949
rect 14956 14940 14968 14943
rect 14875 14912 14968 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 14956 14909 14968 14912
rect 15002 14909 15014 14943
rect 14956 14903 15014 14909
rect 2961 14875 3019 14881
rect 2961 14872 2973 14875
rect 1544 14844 2973 14872
rect 1544 14832 1550 14844
rect 2961 14841 2973 14844
rect 3007 14841 3019 14875
rect 2961 14835 3019 14841
rect 4065 14875 4123 14881
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4111 14844 6040 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 106 14764 112 14816
rect 164 14804 170 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 164 14776 1593 14804
rect 164 14764 170 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3651 14807 3709 14813
rect 3651 14804 3663 14807
rect 3108 14776 3663 14804
rect 3108 14764 3114 14776
rect 3651 14773 3663 14776
rect 3697 14773 3709 14807
rect 3651 14767 3709 14773
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 5767 14807 5825 14813
rect 5767 14804 5779 14807
rect 5684 14776 5779 14804
rect 5684 14764 5690 14776
rect 5767 14773 5779 14776
rect 5813 14773 5825 14807
rect 6012 14804 6040 14844
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8113 14875 8171 14881
rect 8113 14872 8125 14875
rect 7984 14844 8125 14872
rect 7984 14832 7990 14844
rect 8113 14841 8125 14844
rect 8159 14872 8171 14875
rect 8297 14875 8355 14881
rect 8297 14872 8309 14875
rect 8159 14844 8309 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 8297 14841 8309 14844
rect 8343 14841 8355 14875
rect 8297 14835 8355 14841
rect 13909 14875 13967 14881
rect 13909 14841 13921 14875
rect 13955 14872 13967 14875
rect 15749 14875 15807 14881
rect 15749 14872 15761 14875
rect 13955 14844 15761 14872
rect 13955 14841 13967 14844
rect 13909 14835 13967 14841
rect 15749 14841 15761 14844
rect 15795 14872 15807 14875
rect 16025 14875 16083 14881
rect 16025 14872 16037 14875
rect 15795 14844 16037 14872
rect 15795 14841 15807 14844
rect 15749 14835 15807 14841
rect 16025 14841 16037 14844
rect 16071 14841 16083 14875
rect 16025 14835 16083 14841
rect 8938 14804 8944 14816
rect 6012 14776 8944 14804
rect 5767 14767 5825 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 15059 14807 15117 14813
rect 15059 14773 15071 14807
rect 15105 14804 15117 14807
rect 16206 14804 16212 14816
rect 15105 14776 16212 14804
rect 15105 14773 15117 14776
rect 15059 14767 15117 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 1104 14714 17756 14736
rect 1104 14662 7288 14714
rect 7340 14662 7352 14714
rect 7404 14662 7416 14714
rect 7468 14662 7480 14714
rect 7532 14662 13595 14714
rect 13647 14662 13659 14714
rect 13711 14662 13723 14714
rect 13775 14662 13787 14714
rect 13839 14662 17756 14714
rect 1104 14640 17756 14662
rect 4798 14600 4804 14612
rect 4264 14572 4804 14600
rect 2409 14535 2467 14541
rect 2409 14501 2421 14535
rect 2455 14532 2467 14535
rect 3050 14532 3056 14544
rect 2455 14504 3056 14532
rect 2455 14501 2467 14504
rect 2409 14495 2467 14501
rect 3050 14492 3056 14504
rect 3108 14492 3114 14544
rect 4264 14541 4292 14572
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 4249 14535 4307 14541
rect 4249 14501 4261 14535
rect 4295 14501 4307 14535
rect 4249 14495 4307 14501
rect 16025 14535 16083 14541
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 16114 14532 16120 14544
rect 16071 14504 16120 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 5684 14436 5733 14464
rect 5684 14424 5690 14436
rect 5721 14433 5733 14436
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9674 14464 9680 14476
rect 9732 14473 9738 14476
rect 9732 14467 9770 14473
rect 8720 14436 9680 14464
rect 8720 14424 8726 14436
rect 9674 14424 9680 14436
rect 9758 14433 9770 14467
rect 9732 14427 9770 14433
rect 9732 14424 9738 14427
rect 2682 14396 2688 14408
rect 2643 14368 2688 14396
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 4522 14396 4528 14408
rect 4483 14368 4528 14396
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 16298 14396 16304 14408
rect 16259 14368 16304 14396
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 1670 14260 1676 14272
rect 1631 14232 1676 14260
rect 1670 14220 1676 14232
rect 1728 14220 1734 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5905 14263 5963 14269
rect 5905 14260 5917 14263
rect 5132 14232 5917 14260
rect 5132 14220 5138 14232
rect 5905 14229 5917 14232
rect 5951 14229 5963 14263
rect 5905 14223 5963 14229
rect 9306 14220 9312 14272
rect 9364 14260 9370 14272
rect 9815 14263 9873 14269
rect 9815 14260 9827 14263
rect 9364 14232 9827 14260
rect 9364 14220 9370 14232
rect 9815 14229 9827 14232
rect 9861 14229 9873 14263
rect 9815 14223 9873 14229
rect 1104 14170 17756 14192
rect 1104 14118 4135 14170
rect 4187 14118 4199 14170
rect 4251 14118 4263 14170
rect 4315 14118 4327 14170
rect 4379 14118 10441 14170
rect 10493 14118 10505 14170
rect 10557 14118 10569 14170
rect 10621 14118 10633 14170
rect 10685 14118 16748 14170
rect 16800 14118 16812 14170
rect 16864 14118 16876 14170
rect 16928 14118 16940 14170
rect 16992 14118 17756 14170
rect 1104 14096 17756 14118
rect 2777 14059 2835 14065
rect 2777 14025 2789 14059
rect 2823 14056 2835 14059
rect 3050 14056 3056 14068
rect 2823 14028 3056 14056
rect 2823 14025 2835 14028
rect 2777 14019 2835 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 4798 14056 4804 14068
rect 4759 14028 4804 14056
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5813 14059 5871 14065
rect 5813 14056 5825 14059
rect 5684 14028 5825 14056
rect 5684 14016 5690 14028
rect 5813 14025 5825 14028
rect 5859 14025 5871 14059
rect 9306 14056 9312 14068
rect 9267 14028 9312 14056
rect 5813 14019 5871 14025
rect 9306 14016 9312 14028
rect 9364 14016 9370 14068
rect 9674 14056 9680 14068
rect 9635 14028 9680 14056
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 16025 14059 16083 14065
rect 16025 14025 16037 14059
rect 16071 14056 16083 14059
rect 16114 14056 16120 14068
rect 16071 14028 16120 14056
rect 16071 14025 16083 14028
rect 16025 14019 16083 14025
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16482 14056 16488 14068
rect 16443 14028 16488 14056
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 2314 13988 2320 14000
rect 2275 13960 2320 13988
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 2976 13960 4660 13988
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 1946 13920 1952 13932
rect 1811 13892 1952 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 1946 13880 1952 13892
rect 2004 13920 2010 13932
rect 2976 13920 3004 13960
rect 4522 13920 4528 13932
rect 2004 13892 3004 13920
rect 4483 13892 4528 13920
rect 2004 13880 2010 13892
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4632 13920 4660 13960
rect 5353 13923 5411 13929
rect 5353 13920 5365 13923
rect 4632 13892 5365 13920
rect 5353 13889 5365 13892
rect 5399 13889 5411 13923
rect 5353 13883 5411 13889
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13852 8723 13855
rect 9306 13852 9312 13864
rect 8711 13824 9312 13852
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16301 13855 16359 13861
rect 16301 13852 16313 13855
rect 16264 13824 16313 13852
rect 16264 13812 16270 13824
rect 16301 13821 16313 13824
rect 16347 13852 16359 13855
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16347 13824 16865 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 3697 13787 3755 13793
rect 3697 13753 3709 13787
rect 3743 13784 3755 13787
rect 3878 13784 3884 13796
rect 3743 13756 3884 13784
rect 3743 13753 3755 13756
rect 3697 13747 3755 13753
rect 3878 13744 3884 13756
rect 3936 13744 3942 13796
rect 8849 13719 8907 13725
rect 8849 13685 8861 13719
rect 8895 13716 8907 13719
rect 9030 13716 9036 13728
rect 8895 13688 9036 13716
rect 8895 13685 8907 13688
rect 8849 13679 8907 13685
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 14642 13716 14648 13728
rect 14603 13688 14648 13716
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 1104 13626 17756 13648
rect 1104 13574 7288 13626
rect 7340 13574 7352 13626
rect 7404 13574 7416 13626
rect 7468 13574 7480 13626
rect 7532 13574 13595 13626
rect 13647 13574 13659 13626
rect 13711 13574 13723 13626
rect 13775 13574 13787 13626
rect 13839 13574 17756 13626
rect 1104 13552 17756 13574
rect 1765 13515 1823 13521
rect 1765 13481 1777 13515
rect 1811 13512 1823 13515
rect 1946 13512 1952 13524
rect 1811 13484 1952 13512
rect 1811 13481 1823 13484
rect 1765 13475 1823 13481
rect 1946 13472 1952 13484
rect 2004 13472 2010 13524
rect 2038 13444 2044 13456
rect 1951 13416 2044 13444
rect 2038 13404 2044 13416
rect 2096 13444 2102 13456
rect 2682 13444 2688 13456
rect 2096 13416 2688 13444
rect 2096 13404 2102 13416
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 15381 13447 15439 13453
rect 15381 13444 15393 13447
rect 14700 13416 15393 13444
rect 14700 13404 14706 13416
rect 15381 13413 15393 13416
rect 15427 13444 15439 13447
rect 15746 13444 15752 13456
rect 15427 13416 15752 13444
rect 15427 13413 15439 13416
rect 15381 13407 15439 13413
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 16022 13444 16028 13456
rect 15983 13416 16028 13444
rect 16022 13404 16028 13416
rect 16080 13404 16086 13456
rect 4132 13379 4190 13385
rect 4132 13345 4144 13379
rect 4178 13376 4190 13379
rect 4522 13376 4528 13388
rect 4178 13348 4528 13376
rect 4178 13345 4190 13348
rect 4132 13339 4190 13345
rect 4522 13336 4528 13348
rect 4580 13336 4586 13388
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 3234 13132 3240 13184
rect 3292 13172 3298 13184
rect 4203 13175 4261 13181
rect 4203 13172 4215 13175
rect 3292 13144 4215 13172
rect 3292 13132 3298 13144
rect 4203 13141 4215 13144
rect 4249 13141 4261 13175
rect 4203 13135 4261 13141
rect 1104 13082 17756 13104
rect 1104 13030 4135 13082
rect 4187 13030 4199 13082
rect 4251 13030 4263 13082
rect 4315 13030 4327 13082
rect 4379 13030 10441 13082
rect 10493 13030 10505 13082
rect 10557 13030 10569 13082
rect 10621 13030 10633 13082
rect 10685 13030 16748 13082
rect 16800 13030 16812 13082
rect 16864 13030 16876 13082
rect 16928 13030 16940 13082
rect 16992 13030 17756 13082
rect 1104 13008 17756 13030
rect 1535 12971 1593 12977
rect 1535 12937 1547 12971
rect 1581 12968 1593 12971
rect 1670 12968 1676 12980
rect 1581 12940 1676 12968
rect 1581 12937 1593 12940
rect 1535 12931 1593 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 3234 12968 3240 12980
rect 3195 12940 3240 12968
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4522 12968 4528 12980
rect 4203 12940 4528 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4522 12928 4528 12940
rect 4580 12928 4586 12980
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16022 12928 16028 12980
rect 16080 12968 16086 12980
rect 16117 12971 16175 12977
rect 16117 12968 16129 12971
rect 16080 12940 16129 12968
rect 16080 12928 16086 12940
rect 16117 12937 16129 12940
rect 16163 12937 16175 12971
rect 16117 12931 16175 12937
rect 106 12860 112 12912
rect 164 12900 170 12912
rect 3513 12903 3571 12909
rect 3513 12900 3525 12903
rect 164 12872 3525 12900
rect 164 12860 170 12872
rect 3513 12869 3525 12872
rect 3559 12869 3571 12903
rect 3513 12863 3571 12869
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 3936 12804 4445 12832
rect 3936 12792 3942 12804
rect 4433 12801 4445 12804
rect 4479 12801 4491 12835
rect 16040 12832 16068 12928
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12900 16543 12903
rect 17126 12900 17132 12912
rect 16531 12872 17132 12900
rect 16531 12869 16543 12872
rect 16485 12863 16543 12869
rect 17126 12860 17132 12872
rect 17184 12860 17190 12912
rect 4433 12795 4491 12801
rect 15371 12804 16068 12832
rect 1464 12767 1522 12773
rect 1464 12733 1476 12767
rect 1510 12764 1522 12767
rect 2314 12764 2320 12776
rect 1510 12736 2320 12764
rect 1510 12733 1522 12736
rect 1464 12727 1522 12733
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 15371 12773 15399 12804
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 3292 12736 3341 12764
rect 3292 12724 3298 12736
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 15340 12767 15399 12773
rect 15340 12733 15352 12767
rect 15386 12736 15399 12767
rect 15427 12767 15485 12773
rect 15386 12733 15398 12736
rect 15340 12727 15398 12733
rect 15427 12733 15439 12767
rect 15473 12764 15485 12767
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 15473 12736 16313 12764
rect 15473 12733 15485 12736
rect 15427 12727 15485 12733
rect 16301 12733 16313 12736
rect 16347 12764 16359 12767
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 16347 12736 16865 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 16853 12733 16865 12736
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 1104 12538 17756 12560
rect 1104 12486 7288 12538
rect 7340 12486 7352 12538
rect 7404 12486 7416 12538
rect 7468 12486 7480 12538
rect 7532 12486 13595 12538
rect 13647 12486 13659 12538
rect 13711 12486 13723 12538
rect 13775 12486 13787 12538
rect 13839 12486 17756 12538
rect 1104 12464 17756 12486
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 1104 11994 17756 12016
rect 1104 11942 4135 11994
rect 4187 11942 4199 11994
rect 4251 11942 4263 11994
rect 4315 11942 4327 11994
rect 4379 11942 10441 11994
rect 10493 11942 10505 11994
rect 10557 11942 10569 11994
rect 10621 11942 10633 11994
rect 10685 11942 16748 11994
rect 16800 11942 16812 11994
rect 16864 11942 16876 11994
rect 16928 11942 16940 11994
rect 16992 11942 17756 11994
rect 1104 11920 17756 11942
rect 1535 11883 1593 11889
rect 1535 11849 1547 11883
rect 1581 11880 1593 11883
rect 1670 11880 1676 11892
rect 1581 11852 1676 11880
rect 1581 11849 1593 11852
rect 1535 11843 1593 11849
rect 1670 11840 1676 11852
rect 1728 11880 1734 11892
rect 2225 11883 2283 11889
rect 2225 11880 2237 11883
rect 1728 11852 2237 11880
rect 1728 11840 1734 11852
rect 2225 11849 2237 11852
rect 2271 11849 2283 11883
rect 2225 11843 2283 11849
rect 1464 11679 1522 11685
rect 1464 11645 1476 11679
rect 1510 11676 1522 11679
rect 1670 11676 1676 11688
rect 1510 11648 1676 11676
rect 1510 11645 1522 11648
rect 1464 11639 1522 11645
rect 1670 11636 1676 11648
rect 1728 11676 1734 11688
rect 1857 11679 1915 11685
rect 1857 11676 1869 11679
rect 1728 11648 1869 11676
rect 1728 11636 1734 11648
rect 1857 11645 1869 11648
rect 1903 11645 1915 11679
rect 1857 11639 1915 11645
rect 1104 11450 17756 11472
rect 1104 11398 7288 11450
rect 7340 11398 7352 11450
rect 7404 11398 7416 11450
rect 7468 11398 7480 11450
rect 7532 11398 13595 11450
rect 13647 11398 13659 11450
rect 13711 11398 13723 11450
rect 13775 11398 13787 11450
rect 13839 11398 17756 11450
rect 1104 11376 17756 11398
rect 4132 11203 4190 11209
rect 4132 11169 4144 11203
rect 4178 11200 4190 11203
rect 4614 11200 4620 11212
rect 4178 11172 4620 11200
rect 4178 11169 4190 11172
rect 4132 11163 4190 11169
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 16022 11132 16028 11144
rect 15983 11104 16028 11132
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 16114 11092 16120 11144
rect 16172 11132 16178 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 16172 11104 16313 11132
rect 16172 11092 16178 11104
rect 16301 11101 16313 11104
rect 16347 11101 16359 11135
rect 16301 11095 16359 11101
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 4203 10999 4261 11005
rect 4203 10996 4215 10999
rect 3660 10968 4215 10996
rect 3660 10956 3666 10968
rect 4203 10965 4215 10968
rect 4249 10965 4261 10999
rect 4203 10959 4261 10965
rect 1104 10906 17756 10928
rect 1104 10854 4135 10906
rect 4187 10854 4199 10906
rect 4251 10854 4263 10906
rect 4315 10854 4327 10906
rect 4379 10854 10441 10906
rect 10493 10854 10505 10906
rect 10557 10854 10569 10906
rect 10621 10854 10633 10906
rect 10685 10854 16748 10906
rect 16800 10854 16812 10906
rect 16864 10854 16876 10906
rect 16928 10854 16940 10906
rect 16992 10854 17756 10906
rect 1104 10832 17756 10854
rect 4614 10792 4620 10804
rect 4575 10764 4620 10792
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16577 10795 16635 10801
rect 16577 10792 16589 10795
rect 16080 10764 16589 10792
rect 16080 10752 16086 10764
rect 16577 10761 16589 10764
rect 16623 10761 16635 10795
rect 16577 10755 16635 10761
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 3602 10656 3608 10668
rect 3467 10628 3608 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3881 10659 3939 10665
rect 3881 10656 3893 10659
rect 3844 10628 3893 10656
rect 3844 10616 3850 10628
rect 3881 10625 3893 10628
rect 3927 10625 3939 10659
rect 15930 10656 15936 10668
rect 15891 10628 15936 10656
rect 3881 10619 3939 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 106 10548 112 10600
rect 164 10588 170 10600
rect 1578 10588 1584 10600
rect 164 10560 1584 10588
rect 164 10548 170 10560
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10489 1915 10523
rect 1857 10483 1915 10489
rect 2501 10523 2559 10529
rect 2501 10489 2513 10523
rect 2547 10520 2559 10523
rect 2774 10520 2780 10532
rect 2547 10492 2780 10520
rect 2547 10489 2559 10492
rect 2501 10483 2559 10489
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10452 1642 10464
rect 1872 10452 1900 10483
rect 2774 10480 2780 10492
rect 2832 10480 2838 10532
rect 15657 10523 15715 10529
rect 15657 10489 15669 10523
rect 15703 10489 15715 10523
rect 15657 10483 15715 10489
rect 1636 10424 1900 10452
rect 14553 10455 14611 10461
rect 1636 10412 1642 10424
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 15381 10455 15439 10461
rect 15381 10452 15393 10455
rect 14599 10424 15393 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 15381 10421 15393 10424
rect 15427 10452 15439 10455
rect 15672 10452 15700 10483
rect 15427 10424 15700 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 1104 10362 17756 10384
rect 1104 10310 7288 10362
rect 7340 10310 7352 10362
rect 7404 10310 7416 10362
rect 7468 10310 7480 10362
rect 7532 10310 13595 10362
rect 13647 10310 13659 10362
rect 13711 10310 13723 10362
rect 13775 10310 13787 10362
rect 13839 10310 17756 10362
rect 1104 10288 17756 10310
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 16439 10251 16497 10257
rect 16439 10248 16451 10251
rect 16080 10220 16451 10248
rect 16080 10208 16086 10220
rect 16439 10217 16451 10220
rect 16485 10217 16497 10251
rect 16439 10211 16497 10217
rect 1464 10115 1522 10121
rect 1464 10081 1476 10115
rect 1510 10112 1522 10115
rect 2038 10112 2044 10124
rect 1510 10084 2044 10112
rect 1510 10081 1522 10084
rect 1464 10075 1522 10081
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 15378 10121 15384 10124
rect 15356 10115 15384 10121
rect 15356 10112 15368 10115
rect 15291 10084 15368 10112
rect 15356 10081 15368 10084
rect 15436 10112 15442 10124
rect 15930 10112 15936 10124
rect 15436 10084 15936 10112
rect 15356 10075 15384 10081
rect 15378 10072 15384 10075
rect 15436 10072 15442 10084
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 16368 10115 16426 10121
rect 16368 10081 16380 10115
rect 16414 10112 16426 10115
rect 17034 10112 17040 10124
rect 16414 10084 17040 10112
rect 16414 10081 16426 10084
rect 16368 10075 16426 10081
rect 17034 10072 17040 10084
rect 17092 10072 17098 10124
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2774 10044 2780 10056
rect 2735 10016 2780 10044
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 1486 9908 1492 9920
rect 1445 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9917 1550 9920
rect 1544 9911 1593 9917
rect 1544 9877 1547 9911
rect 1581 9908 1593 9911
rect 1857 9911 1915 9917
rect 1857 9908 1869 9911
rect 1581 9880 1869 9908
rect 1581 9877 1593 9880
rect 1544 9871 1593 9877
rect 1857 9877 1869 9880
rect 1903 9877 1915 9911
rect 1857 9871 1915 9877
rect 15427 9911 15485 9917
rect 15427 9877 15439 9911
rect 15473 9908 15485 9911
rect 16114 9908 16120 9920
rect 15473 9880 16120 9908
rect 15473 9877 15485 9880
rect 15427 9871 15485 9877
rect 1544 9868 1550 9871
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 1104 9818 17756 9840
rect 1104 9766 4135 9818
rect 4187 9766 4199 9818
rect 4251 9766 4263 9818
rect 4315 9766 4327 9818
rect 4379 9766 10441 9818
rect 10493 9766 10505 9818
rect 10557 9766 10569 9818
rect 10621 9766 10633 9818
rect 10685 9766 16748 9818
rect 16800 9766 16812 9818
rect 16864 9766 16876 9818
rect 16928 9766 16940 9818
rect 16992 9766 17756 9818
rect 1104 9744 17756 9766
rect 1302 9664 1308 9716
rect 1360 9704 1366 9716
rect 1581 9707 1639 9713
rect 1581 9704 1593 9707
rect 1360 9676 1593 9704
rect 1360 9664 1366 9676
rect 1581 9673 1593 9676
rect 1627 9673 1639 9707
rect 2038 9704 2044 9716
rect 1951 9676 2044 9704
rect 1581 9667 1639 9673
rect 2038 9664 2044 9676
rect 2096 9704 2102 9716
rect 2774 9704 2780 9716
rect 2096 9676 2780 9704
rect 2096 9664 2102 9676
rect 2774 9664 2780 9676
rect 2832 9664 2838 9716
rect 7377 9707 7435 9713
rect 7377 9673 7389 9707
rect 7423 9704 7435 9707
rect 12434 9704 12440 9716
rect 7423 9676 12440 9704
rect 7423 9673 7435 9676
rect 7377 9667 7435 9673
rect 2498 9568 2504 9580
rect 2411 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9568 2562 9580
rect 3786 9568 3792 9580
rect 2556 9540 3792 9568
rect 2556 9528 2562 9540
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1486 9500 1492 9512
rect 1443 9472 1492 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 6892 9503 6950 9509
rect 6892 9469 6904 9503
rect 6938 9500 6950 9503
rect 7392 9500 7420 9667
rect 12434 9664 12440 9676
rect 12492 9664 12498 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 16114 9704 16120 9716
rect 16075 9676 16120 9704
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 16485 9639 16543 9645
rect 16485 9605 16497 9639
rect 16531 9636 16543 9639
rect 18414 9636 18420 9648
rect 16531 9608 18420 9636
rect 16531 9605 16543 9608
rect 16485 9599 16543 9605
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 6938 9472 7420 9500
rect 6938 9469 6950 9472
rect 6892 9463 6950 9469
rect 16114 9460 16120 9512
rect 16172 9500 16178 9512
rect 16301 9503 16359 9509
rect 16301 9500 16313 9503
rect 16172 9472 16313 9500
rect 16172 9460 16178 9472
rect 16301 9469 16313 9472
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 2958 9432 2964 9444
rect 2871 9404 2964 9432
rect 2958 9392 2964 9404
rect 3016 9432 3022 9444
rect 3145 9435 3203 9441
rect 3145 9432 3157 9435
rect 3016 9404 3157 9432
rect 3016 9392 3022 9404
rect 3145 9401 3157 9404
rect 3191 9401 3203 9435
rect 3145 9395 3203 9401
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6963 9367 7021 9373
rect 6963 9364 6975 9367
rect 6420 9336 6975 9364
rect 6420 9324 6426 9336
rect 6963 9333 6975 9336
rect 7009 9333 7021 9367
rect 6963 9327 7021 9333
rect 16945 9367 17003 9373
rect 16945 9333 16957 9367
rect 16991 9364 17003 9367
rect 17034 9364 17040 9376
rect 16991 9336 17040 9364
rect 16991 9333 17003 9336
rect 16945 9327 17003 9333
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 1104 9274 17756 9296
rect 1104 9222 7288 9274
rect 7340 9222 7352 9274
rect 7404 9222 7416 9274
rect 7468 9222 7480 9274
rect 7532 9222 13595 9274
rect 13647 9222 13659 9274
rect 13711 9222 13723 9274
rect 13775 9222 13787 9274
rect 13839 9222 17756 9274
rect 1104 9200 17756 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 2823 9163 2881 9169
rect 2823 9129 2835 9163
rect 2869 9160 2881 9163
rect 2958 9160 2964 9172
rect 2869 9132 2964 9160
rect 2869 9129 2881 9132
rect 2823 9123 2881 9129
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 16482 9160 16488 9172
rect 16443 9132 16488 9160
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 6362 9092 6368 9104
rect 6323 9064 6368 9092
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 15194 9024 15200 9036
rect 15155 8996 15200 9024
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 15427 9027 15485 9033
rect 15427 8993 15439 9027
rect 15473 9024 15485 9027
rect 16298 9024 16304 9036
rect 15473 8996 16304 9024
rect 15473 8993 15485 8996
rect 15427 8987 15485 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 5960 8928 6653 8956
rect 5960 8916 5966 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6641 8919 6699 8925
rect 2590 8820 2596 8832
rect 2551 8792 2596 8820
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 1104 8730 17756 8752
rect 1104 8678 4135 8730
rect 4187 8678 4199 8730
rect 4251 8678 4263 8730
rect 4315 8678 4327 8730
rect 4379 8678 10441 8730
rect 10493 8678 10505 8730
rect 10557 8678 10569 8730
rect 10621 8678 10633 8730
rect 10685 8678 16748 8730
rect 16800 8678 16812 8730
rect 16864 8678 16876 8730
rect 16928 8678 16940 8730
rect 16992 8678 17756 8730
rect 1104 8656 17756 8678
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15289 8619 15347 8625
rect 15289 8616 15301 8619
rect 15252 8588 15301 8616
rect 15252 8576 15258 8588
rect 15289 8585 15301 8588
rect 15335 8585 15347 8619
rect 15289 8579 15347 8585
rect 5902 8480 5908 8492
rect 5863 8452 5908 8480
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 15304 8480 15332 8579
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16853 8619 16911 8625
rect 16853 8616 16865 8619
rect 16356 8588 16865 8616
rect 16356 8576 16362 8588
rect 16853 8585 16865 8588
rect 16899 8585 16911 8619
rect 16853 8579 16911 8585
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 15304 8452 16221 8480
rect 16209 8449 16221 8452
rect 16255 8480 16267 8483
rect 16390 8480 16396 8492
rect 16255 8452 16396 8480
rect 16255 8449 16267 8452
rect 16209 8443 16267 8449
rect 16390 8440 16396 8452
rect 16448 8440 16454 8492
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 5000 8316 5273 8344
rect 5000 8288 5028 8316
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 14829 8347 14887 8353
rect 14829 8313 14841 8347
rect 14875 8344 14887 8347
rect 15657 8347 15715 8353
rect 15657 8344 15669 8347
rect 14875 8316 15669 8344
rect 14875 8313 14887 8316
rect 14829 8307 14887 8313
rect 15657 8313 15669 8316
rect 15703 8344 15715 8347
rect 15933 8347 15991 8353
rect 15933 8344 15945 8347
rect 15703 8316 15945 8344
rect 15703 8313 15715 8316
rect 15657 8307 15715 8313
rect 15933 8313 15945 8316
rect 15979 8313 15991 8347
rect 15933 8307 15991 8313
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 2777 8279 2835 8285
rect 2777 8276 2789 8279
rect 2648 8248 2789 8276
rect 2648 8236 2654 8248
rect 2777 8245 2789 8248
rect 2823 8276 2835 8279
rect 3234 8276 3240 8288
rect 2823 8248 3240 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 4982 8276 4988 8288
rect 4943 8248 4988 8276
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 1104 8186 17756 8208
rect 1104 8134 7288 8186
rect 7340 8134 7352 8186
rect 7404 8134 7416 8186
rect 7468 8134 7480 8186
rect 7532 8134 13595 8186
rect 13647 8134 13659 8186
rect 13711 8134 13723 8186
rect 13775 8134 13787 8186
rect 13839 8134 17756 8186
rect 1104 8112 17756 8134
rect 4571 8075 4629 8081
rect 4571 8041 4583 8075
rect 4617 8072 4629 8075
rect 4982 8072 4988 8084
rect 4617 8044 4988 8072
rect 4617 8041 4629 8044
rect 4571 8035 4629 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 6362 8004 6368 8016
rect 5960 7976 6368 8004
rect 5960 7964 5966 7976
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 4430 7936 4436 7948
rect 4391 7908 4436 7936
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 14252 7939 14310 7945
rect 14252 7905 14264 7939
rect 14298 7936 14310 7939
rect 14826 7936 14832 7948
rect 14298 7908 14832 7936
rect 14298 7905 14310 7908
rect 14252 7899 14310 7905
rect 14826 7896 14832 7908
rect 14884 7896 14890 7948
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16298 7868 16304 7880
rect 16071 7840 16304 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16448 7840 16493 7868
rect 16448 7828 16454 7840
rect 14323 7735 14381 7741
rect 14323 7701 14335 7735
rect 14369 7732 14381 7735
rect 15378 7732 15384 7744
rect 14369 7704 15384 7732
rect 14369 7701 14381 7704
rect 14323 7695 14381 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 1104 7642 17756 7664
rect 1104 7590 4135 7642
rect 4187 7590 4199 7642
rect 4251 7590 4263 7642
rect 4315 7590 4327 7642
rect 4379 7590 10441 7642
rect 10493 7590 10505 7642
rect 10557 7590 10569 7642
rect 10621 7590 10633 7642
rect 10685 7590 16748 7642
rect 16800 7590 16812 7642
rect 16864 7590 16876 7642
rect 16928 7590 16940 7642
rect 16992 7590 17756 7642
rect 1104 7568 17756 7590
rect 4430 7528 4436 7540
rect 4391 7500 4436 7528
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 6362 7528 6368 7540
rect 6323 7500 6368 7528
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 14458 7528 14464 7540
rect 14419 7500 14464 7528
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 14826 7528 14832 7540
rect 14787 7500 14832 7528
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 16298 7392 16304 7404
rect 16259 7364 16304 7392
rect 16298 7352 16304 7364
rect 16356 7392 16362 7404
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16356 7364 16957 7392
rect 16356 7352 16362 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 13960 7327 14018 7333
rect 13960 7293 13972 7327
rect 14006 7324 14018 7327
rect 14458 7324 14464 7336
rect 14006 7296 14464 7324
rect 14006 7293 14018 7296
rect 13960 7287 14018 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14972 7327 15030 7333
rect 14972 7293 14984 7327
rect 15018 7324 15030 7327
rect 15470 7324 15476 7336
rect 15018 7296 15476 7324
rect 15018 7293 15030 7296
rect 14972 7287 15030 7293
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 14047 7259 14105 7265
rect 14047 7225 14059 7259
rect 14093 7256 14105 7259
rect 14826 7256 14832 7268
rect 14093 7228 14832 7256
rect 14093 7225 14105 7228
rect 14047 7219 14105 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 15059 7259 15117 7265
rect 15059 7225 15071 7259
rect 15105 7256 15117 7259
rect 15749 7259 15807 7265
rect 15749 7256 15761 7259
rect 15105 7228 15761 7256
rect 15105 7225 15117 7228
rect 15059 7219 15117 7225
rect 15749 7225 15761 7228
rect 15795 7256 15807 7259
rect 16025 7259 16083 7265
rect 16025 7256 16037 7259
rect 15795 7228 16037 7256
rect 15795 7225 15807 7228
rect 15749 7219 15807 7225
rect 16025 7225 16037 7228
rect 16071 7225 16083 7259
rect 16025 7219 16083 7225
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 1104 7098 17756 7120
rect 1104 7046 7288 7098
rect 7340 7046 7352 7098
rect 7404 7046 7416 7098
rect 7468 7046 7480 7098
rect 7532 7046 13595 7098
rect 13647 7046 13659 7098
rect 13711 7046 13723 7098
rect 13775 7046 13787 7098
rect 13839 7046 17756 7098
rect 1104 7024 17756 7046
rect 6362 6916 6368 6928
rect 6275 6888 6368 6916
rect 6362 6876 6368 6888
rect 6420 6916 6426 6928
rect 6822 6916 6828 6928
rect 6420 6888 6828 6916
rect 6420 6876 6426 6888
rect 6822 6876 6828 6888
rect 6880 6876 6886 6928
rect 7006 6916 7012 6928
rect 6967 6888 7012 6916
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7024 6848 7052 6876
rect 7834 6848 7840 6860
rect 7892 6857 7898 6860
rect 7892 6851 7930 6857
rect 7024 6820 7840 6848
rect 7834 6808 7840 6820
rect 7918 6817 7930 6851
rect 7892 6811 7930 6817
rect 12688 6851 12746 6857
rect 12688 6817 12700 6851
rect 12734 6848 12746 6851
rect 13446 6848 13452 6860
rect 12734 6820 13452 6848
rect 12734 6817 12746 6820
rect 12688 6811 12746 6817
rect 7892 6808 7898 6811
rect 13446 6808 13452 6820
rect 13504 6808 13510 6860
rect 15930 6780 15936 6792
rect 15891 6752 15936 6780
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 14093 6715 14151 6721
rect 14093 6681 14105 6715
rect 14139 6712 14151 6715
rect 14458 6712 14464 6724
rect 14139 6684 14464 6712
rect 14139 6681 14151 6684
rect 14093 6675 14151 6681
rect 14458 6672 14464 6684
rect 14516 6672 14522 6724
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7975 6647 8033 6653
rect 7975 6644 7987 6647
rect 7524 6616 7987 6644
rect 7524 6604 7530 6616
rect 7975 6613 7987 6616
rect 8021 6613 8033 6647
rect 7975 6607 8033 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 12759 6647 12817 6653
rect 12759 6644 12771 6647
rect 11020 6616 12771 6644
rect 11020 6604 11026 6616
rect 12759 6613 12771 6616
rect 12805 6613 12817 6647
rect 12759 6607 12817 6613
rect 14323 6647 14381 6653
rect 14323 6613 14335 6647
rect 14369 6644 14381 6647
rect 15286 6644 15292 6656
rect 14369 6616 15292 6644
rect 14369 6613 14381 6616
rect 14323 6607 14381 6613
rect 15286 6604 15292 6616
rect 15344 6604 15350 6656
rect 1104 6554 17756 6576
rect 1104 6502 4135 6554
rect 4187 6502 4199 6554
rect 4251 6502 4263 6554
rect 4315 6502 4327 6554
rect 4379 6502 10441 6554
rect 10493 6502 10505 6554
rect 10557 6502 10569 6554
rect 10621 6502 10633 6554
rect 10685 6502 16748 6554
rect 16800 6502 16812 6554
rect 16864 6502 16876 6554
rect 16928 6502 16940 6554
rect 16992 6502 17756 6554
rect 1104 6480 17756 6502
rect 6362 6440 6368 6452
rect 6323 6412 6368 6440
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 7466 6440 7472 6452
rect 7427 6412 7472 6440
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 7834 6440 7840 6452
rect 7795 6412 7840 6440
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 15795 6443 15853 6449
rect 15795 6409 15807 6443
rect 15841 6440 15853 6443
rect 15930 6440 15936 6452
rect 15841 6412 15936 6440
rect 15841 6409 15853 6412
rect 15795 6403 15853 6409
rect 15930 6400 15936 6412
rect 15988 6440 15994 6452
rect 16485 6443 16543 6449
rect 16485 6440 16497 6443
rect 15988 6412 16497 6440
rect 15988 6400 15994 6412
rect 16485 6409 16497 6412
rect 16531 6409 16543 6443
rect 16485 6403 16543 6409
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 17126 6372 17132 6384
rect 15243 6344 17132 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6304 13231 6307
rect 14550 6304 14556 6316
rect 13219 6276 14556 6304
rect 13219 6273 13231 6276
rect 13173 6267 13231 6273
rect 6825 6239 6883 6245
rect 6825 6205 6837 6239
rect 6871 6236 6883 6239
rect 7466 6236 7472 6248
rect 6871 6208 7472 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 12688 6239 12746 6245
rect 12688 6205 12700 6239
rect 12734 6236 12746 6239
rect 13188 6236 13216 6267
rect 14550 6264 14556 6276
rect 14608 6264 14614 6316
rect 12734 6208 13216 6236
rect 13700 6239 13758 6245
rect 12734 6205 12746 6208
rect 12688 6199 12746 6205
rect 13700 6205 13712 6239
rect 13746 6236 13758 6239
rect 14712 6239 14770 6245
rect 13746 6208 14228 6236
rect 13746 6205 13758 6208
rect 13700 6199 13758 6205
rect 14200 6112 14228 6208
rect 14712 6205 14724 6239
rect 14758 6236 14770 6239
rect 15212 6236 15240 6335
rect 17126 6332 17132 6344
rect 17184 6332 17190 6384
rect 17218 6304 17224 6316
rect 14758 6208 15240 6236
rect 15304 6276 17224 6304
rect 14758 6205 14770 6208
rect 14712 6199 14770 6205
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 14553 6171 14611 6177
rect 14553 6168 14565 6171
rect 14516 6140 14565 6168
rect 14516 6128 14522 6140
rect 14553 6137 14565 6140
rect 14599 6168 14611 6171
rect 15304 6168 15332 6276
rect 17218 6264 17224 6276
rect 17276 6264 17282 6316
rect 15724 6239 15782 6245
rect 15724 6205 15736 6239
rect 15770 6236 15782 6239
rect 15770 6208 16252 6236
rect 15770 6205 15782 6208
rect 15724 6199 15782 6205
rect 14599 6140 15332 6168
rect 14599 6137 14611 6140
rect 14553 6131 14611 6137
rect 16224 6112 16252 6208
rect 7009 6103 7067 6109
rect 7009 6069 7021 6103
rect 7055 6100 7067 6103
rect 7098 6100 7104 6112
rect 7055 6072 7104 6100
rect 7055 6069 7067 6072
rect 7009 6063 7067 6069
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 12759 6103 12817 6109
rect 12759 6069 12771 6103
rect 12805 6100 12817 6103
rect 12986 6100 12992 6112
rect 12805 6072 12992 6100
rect 12805 6069 12817 6072
rect 12759 6063 12817 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13446 6100 13452 6112
rect 13407 6072 13452 6100
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13771 6103 13829 6109
rect 13771 6069 13783 6103
rect 13817 6100 13829 6103
rect 13906 6100 13912 6112
rect 13817 6072 13912 6100
rect 13817 6069 13829 6072
rect 13771 6063 13829 6069
rect 13906 6060 13912 6072
rect 13964 6060 13970 6112
rect 14182 6100 14188 6112
rect 14143 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 14783 6103 14841 6109
rect 14783 6069 14795 6103
rect 14829 6100 14841 6103
rect 15010 6100 15016 6112
rect 14829 6072 15016 6100
rect 14829 6069 14841 6072
rect 14783 6063 14841 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 16206 6100 16212 6112
rect 16167 6072 16212 6100
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 1104 6010 17756 6032
rect 1104 5958 7288 6010
rect 7340 5958 7352 6010
rect 7404 5958 7416 6010
rect 7468 5958 7480 6010
rect 7532 5958 13595 6010
rect 13647 5958 13659 6010
rect 13711 5958 13723 6010
rect 13775 5958 13787 6010
rect 13839 5958 17756 6010
rect 1104 5936 17756 5958
rect 15378 5828 15384 5840
rect 15339 5800 15384 5828
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 12526 5692 12532 5704
rect 12487 5664 12532 5692
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 1104 5466 17756 5488
rect 1104 5414 4135 5466
rect 4187 5414 4199 5466
rect 4251 5414 4263 5466
rect 4315 5414 4327 5466
rect 4379 5414 10441 5466
rect 10493 5414 10505 5466
rect 10557 5414 10569 5466
rect 10621 5414 10633 5466
rect 10685 5414 16748 5466
rect 16800 5414 16812 5466
rect 16864 5414 16876 5466
rect 16928 5414 16940 5466
rect 16992 5414 17756 5466
rect 1104 5392 17756 5414
rect 15010 5312 15016 5364
rect 15068 5352 15074 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 15068 5324 15761 5352
rect 15068 5312 15074 5324
rect 15749 5321 15761 5324
rect 15795 5352 15807 5355
rect 15795 5324 16068 5352
rect 15795 5321 15807 5324
rect 15749 5315 15807 5321
rect 15378 5284 15384 5296
rect 15339 5256 15384 5284
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 15470 5216 15476 5228
rect 11931 5188 15476 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 9928 5151 9986 5157
rect 9928 5117 9940 5151
rect 9974 5148 9986 5151
rect 11400 5151 11458 5157
rect 9974 5120 10456 5148
rect 9974 5117 9986 5120
rect 9928 5111 9986 5117
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 10428 5021 10456 5120
rect 11400 5117 11412 5151
rect 11446 5148 11458 5151
rect 11900 5148 11928 5179
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 16040 5225 16068 5324
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5185 16083 5219
rect 16298 5216 16304 5228
rect 16259 5188 16304 5216
rect 16025 5179 16083 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 11446 5120 11928 5148
rect 11446 5117 11458 5120
rect 11400 5111 11458 5117
rect 11609 5083 11667 5089
rect 11609 5049 11621 5083
rect 11655 5080 11667 5083
rect 12710 5080 12716 5092
rect 11655 5052 12716 5080
rect 11655 5049 11667 5052
rect 11609 5043 11667 5049
rect 12710 5040 12716 5052
rect 12768 5040 12774 5092
rect 13449 5083 13507 5089
rect 13449 5049 13461 5083
rect 13495 5080 13507 5083
rect 13633 5083 13691 5089
rect 13633 5080 13645 5083
rect 13495 5052 13645 5080
rect 13495 5049 13507 5052
rect 13449 5043 13507 5049
rect 13633 5049 13645 5052
rect 13679 5080 13691 5083
rect 13998 5080 14004 5092
rect 13679 5052 14004 5080
rect 13679 5049 13691 5052
rect 13633 5043 13691 5049
rect 13998 5040 14004 5052
rect 14056 5040 14062 5092
rect 14274 5080 14280 5092
rect 14235 5052 14280 5080
rect 14274 5040 14280 5052
rect 14332 5040 14338 5092
rect 9999 5015 10057 5021
rect 9999 5012 10011 5015
rect 9364 4984 10011 5012
rect 9364 4972 9370 4984
rect 9999 4981 10011 4984
rect 10045 4981 10057 5015
rect 9999 4975 10057 4981
rect 10413 5015 10471 5021
rect 10413 4981 10425 5015
rect 10459 5012 10471 5015
rect 11238 5012 11244 5024
rect 10459 4984 11244 5012
rect 10459 4981 10471 4984
rect 10413 4975 10471 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12529 5015 12587 5021
rect 12529 5012 12541 5015
rect 12492 4984 12541 5012
rect 12492 4972 12498 4984
rect 12529 4981 12541 4984
rect 12575 4981 12587 5015
rect 12529 4975 12587 4981
rect 1104 4922 17756 4944
rect 1104 4870 7288 4922
rect 7340 4870 7352 4922
rect 7404 4870 7416 4922
rect 7468 4870 7480 4922
rect 7532 4870 13595 4922
rect 13647 4870 13659 4922
rect 13711 4870 13723 4922
rect 13775 4870 13787 4922
rect 13839 4870 17756 4922
rect 1104 4848 17756 4870
rect 10091 4811 10149 4817
rect 10091 4777 10103 4811
rect 10137 4808 10149 4811
rect 12342 4808 12348 4820
rect 10137 4780 12204 4808
rect 12303 4780 12348 4808
rect 10137 4777 10149 4780
rect 10091 4771 10149 4777
rect 12176 4684 12204 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 13725 4743 13783 4749
rect 13725 4709 13737 4743
rect 13771 4740 13783 4743
rect 13906 4740 13912 4752
rect 13771 4712 13912 4740
rect 13771 4709 13783 4712
rect 13725 4703 13783 4709
rect 13906 4700 13912 4712
rect 13964 4700 13970 4752
rect 13998 4700 14004 4752
rect 14056 4740 14062 4752
rect 14369 4743 14427 4749
rect 14369 4740 14381 4743
rect 14056 4712 14381 4740
rect 14056 4700 14062 4712
rect 14369 4709 14381 4712
rect 14415 4740 14427 4743
rect 15654 4740 15660 4752
rect 14415 4712 15660 4740
rect 14415 4709 14427 4712
rect 14369 4703 14427 4709
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 10020 4675 10078 4681
rect 10020 4641 10032 4675
rect 10066 4672 10078 4675
rect 10226 4672 10232 4684
rect 10066 4644 10232 4672
rect 10066 4641 10078 4644
rect 10020 4635 10078 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 11032 4675 11090 4681
rect 11032 4641 11044 4675
rect 11078 4672 11090 4675
rect 11146 4672 11152 4684
rect 11078 4644 11152 4672
rect 11078 4641 11090 4644
rect 11032 4635 11090 4641
rect 11146 4632 11152 4644
rect 11204 4632 11210 4684
rect 12158 4672 12164 4684
rect 12071 4644 12164 4672
rect 12158 4632 12164 4644
rect 12216 4632 12222 4684
rect 14826 4564 14832 4616
rect 14884 4604 14890 4616
rect 15562 4604 15568 4616
rect 14884 4576 15568 4604
rect 14884 4564 14890 4576
rect 15562 4564 15568 4576
rect 15620 4564 15626 4616
rect 15746 4564 15752 4616
rect 15804 4604 15810 4616
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15804 4576 15853 4604
rect 15804 4564 15810 4576
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 11103 4471 11161 4477
rect 11103 4468 11115 4471
rect 10928 4440 11115 4468
rect 10928 4428 10934 4440
rect 11103 4437 11115 4440
rect 11149 4437 11161 4471
rect 11103 4431 11161 4437
rect 1104 4378 17756 4400
rect 1104 4326 4135 4378
rect 4187 4326 4199 4378
rect 4251 4326 4263 4378
rect 4315 4326 4327 4378
rect 4379 4326 10441 4378
rect 10493 4326 10505 4378
rect 10557 4326 10569 4378
rect 10621 4326 10633 4378
rect 10685 4326 16748 4378
rect 16800 4326 16812 4378
rect 16864 4326 16876 4378
rect 16928 4326 16940 4378
rect 16992 4326 17756 4378
rect 1104 4304 17756 4326
rect 1854 4264 1860 4276
rect 1815 4236 1860 4264
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 12158 4264 12164 4276
rect 12119 4236 12164 4264
rect 12158 4224 12164 4236
rect 12216 4224 12222 4276
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12584 4236 12633 4264
rect 12584 4224 12590 4236
rect 12621 4233 12633 4236
rect 12667 4233 12679 4267
rect 13906 4264 13912 4276
rect 13867 4236 13912 4264
rect 12621 4227 12679 4233
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 10137 4131 10195 4137
rect 2924 4100 9295 4128
rect 2924 4088 2930 4100
rect 1464 4063 1522 4069
rect 1464 4029 1476 4063
rect 1510 4060 1522 4063
rect 1854 4060 1860 4072
rect 1510 4032 1860 4060
rect 1510 4029 1522 4032
rect 1464 4023 1522 4029
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 9267 4069 9295 4100
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10226 4128 10232 4140
rect 10183 4100 10232 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10226 4088 10232 4100
rect 10284 4128 10290 4140
rect 12636 4128 12664 4227
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 16025 4267 16083 4273
rect 16025 4264 16037 4267
rect 15620 4236 16037 4264
rect 15620 4224 15626 4236
rect 16025 4233 16037 4236
rect 16071 4233 16083 4267
rect 16025 4227 16083 4233
rect 12710 4156 12716 4208
rect 12768 4196 12774 4208
rect 14829 4199 14887 4205
rect 14829 4196 14841 4199
rect 12768 4168 14841 4196
rect 12768 4156 12774 4168
rect 14829 4165 14841 4168
rect 14875 4165 14887 4199
rect 14829 4159 14887 4165
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 10284 4100 12020 4128
rect 12636 4100 12909 4128
rect 10284 4088 10290 4100
rect 5388 4063 5446 4069
rect 5388 4060 5400 4063
rect 4028 4032 5400 4060
rect 4028 4020 4034 4032
rect 5388 4029 5400 4032
rect 5434 4060 5446 4063
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5434 4032 5825 4060
rect 5434 4029 5446 4032
rect 5388 4023 5446 4029
rect 5813 4029 5825 4032
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 9252 4063 9310 4069
rect 9252 4029 9264 4063
rect 9298 4060 9310 4063
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9298 4032 9689 4060
rect 9298 4029 9310 4032
rect 9252 4023 9310 4029
rect 9677 4029 9689 4032
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 11400 4063 11458 4069
rect 11400 4029 11412 4063
rect 11446 4060 11458 4063
rect 11446 4032 11928 4060
rect 11446 4029 11458 4032
rect 11400 4023 11458 4029
rect 1535 3927 1593 3933
rect 1535 3893 1547 3927
rect 1581 3924 1593 3927
rect 2130 3924 2136 3936
rect 1581 3896 2136 3924
rect 1581 3893 1593 3896
rect 1535 3887 1593 3893
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 5491 3927 5549 3933
rect 5491 3893 5503 3927
rect 5537 3924 5549 3927
rect 6270 3924 6276 3936
rect 5537 3896 6276 3924
rect 5537 3893 5549 3896
rect 5491 3887 5549 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 7006 3924 7012 3936
rect 6967 3896 7012 3924
rect 7006 3884 7012 3896
rect 7064 3884 7070 3936
rect 9355 3927 9413 3933
rect 9355 3893 9367 3927
rect 9401 3924 9413 3927
rect 9582 3924 9588 3936
rect 9401 3896 9588 3924
rect 9401 3893 9413 3896
rect 9355 3887 9413 3893
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11054 3924 11060 3936
rect 11015 3896 11060 3924
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 11330 3884 11336 3936
rect 11388 3924 11394 3936
rect 11900 3933 11928 4032
rect 11992 3992 12020 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 14844 4128 14872 4159
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14844 4100 15117 4128
rect 12897 4091 12955 4097
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15746 4128 15752 4140
rect 15707 4100 15752 4128
rect 15105 4091 15163 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 13541 3995 13599 4001
rect 13541 3992 13553 3995
rect 11992 3964 13553 3992
rect 13541 3961 13553 3964
rect 13587 3992 13599 3995
rect 14274 3992 14280 4004
rect 13587 3964 14280 3992
rect 13587 3961 13599 3964
rect 13541 3955 13599 3961
rect 14274 3952 14280 3964
rect 14332 3952 14338 4004
rect 11471 3927 11529 3933
rect 11471 3924 11483 3927
rect 11388 3896 11483 3924
rect 11388 3884 11394 3896
rect 11471 3893 11483 3896
rect 11517 3893 11529 3927
rect 11471 3887 11529 3893
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12342 3924 12348 3936
rect 11931 3896 12348 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 1104 3834 17756 3856
rect 1104 3782 7288 3834
rect 7340 3782 7352 3834
rect 7404 3782 7416 3834
rect 7468 3782 7480 3834
rect 7532 3782 13595 3834
rect 13647 3782 13659 3834
rect 13711 3782 13723 3834
rect 13775 3782 13787 3834
rect 13839 3782 17756 3834
rect 1104 3760 17756 3782
rect 2130 3652 2136 3664
rect 2091 3624 2136 3652
rect 2130 3612 2136 3624
rect 2188 3612 2194 3664
rect 6270 3652 6276 3664
rect 6231 3624 6276 3652
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 9582 3612 9588 3664
rect 9640 3652 9646 3664
rect 10137 3655 10195 3661
rect 10137 3652 10149 3655
rect 9640 3624 10149 3652
rect 9640 3612 9646 3624
rect 10137 3621 10149 3624
rect 10183 3652 10195 3655
rect 10226 3652 10232 3664
rect 10183 3624 10232 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 15381 3655 15439 3661
rect 15381 3621 15393 3655
rect 15427 3652 15439 3655
rect 15746 3652 15752 3664
rect 15427 3624 15752 3652
rect 15427 3621 15439 3624
rect 15381 3615 15439 3621
rect 15746 3612 15752 3624
rect 15804 3612 15810 3664
rect 7742 3584 7748 3596
rect 7703 3556 7748 3584
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 12986 3544 12992 3596
rect 13044 3584 13050 3596
rect 13814 3584 13820 3596
rect 13044 3556 13820 3584
rect 13044 3544 13050 3556
rect 13814 3544 13820 3556
rect 13872 3584 13878 3596
rect 13872 3556 13917 3584
rect 13872 3544 13878 3556
rect 2774 3516 2780 3528
rect 2735 3488 2780 3516
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 3936 3488 4169 3516
rect 3936 3476 3942 3488
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 4798 3516 4804 3528
rect 4759 3488 4804 3516
rect 4157 3479 4215 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 6914 3516 6920 3528
rect 6875 3488 6920 3516
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 10781 3519 10839 3525
rect 10781 3485 10793 3519
rect 10827 3516 10839 3519
rect 11422 3516 11428 3528
rect 10827 3488 11428 3516
rect 10827 3485 10839 3488
rect 10781 3479 10839 3485
rect 11422 3476 11428 3488
rect 11480 3516 11486 3528
rect 11701 3519 11759 3525
rect 11701 3516 11713 3519
rect 11480 3488 11713 3516
rect 11480 3476 11486 3488
rect 11701 3485 11713 3488
rect 11747 3485 11759 3519
rect 12342 3516 12348 3528
rect 12303 3488 12348 3516
rect 11701 3479 11759 3485
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 14550 3476 14556 3528
rect 14608 3516 14614 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 14608 3488 15669 3516
rect 14608 3476 14614 3488
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 15657 3479 15715 3485
rect 7929 3383 7987 3389
rect 7929 3349 7941 3383
rect 7975 3380 7987 3383
rect 8202 3380 8208 3392
rect 7975 3352 8208 3380
rect 7975 3349 7987 3352
rect 7929 3343 7987 3349
rect 8202 3340 8208 3352
rect 8260 3340 8266 3392
rect 13998 3380 14004 3392
rect 13959 3352 14004 3380
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 1104 3290 17756 3312
rect 1104 3238 4135 3290
rect 4187 3238 4199 3290
rect 4251 3238 4263 3290
rect 4315 3238 4327 3290
rect 4379 3238 10441 3290
rect 10493 3238 10505 3290
rect 10557 3238 10569 3290
rect 10621 3238 10633 3290
rect 10685 3238 16748 3290
rect 16800 3238 16812 3290
rect 16864 3238 16876 3290
rect 16928 3238 16940 3290
rect 16992 3238 17756 3290
rect 1104 3216 17756 3238
rect 2130 3176 2136 3188
rect 2091 3148 2136 3176
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 10226 3176 10232 3188
rect 10187 3148 10232 3176
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10318 3136 10324 3188
rect 10376 3176 10382 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 10376 3148 12173 3176
rect 10376 3136 10382 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 2774 3068 2780 3120
rect 2832 3108 2838 3120
rect 3786 3108 3792 3120
rect 2832 3080 3792 3108
rect 2832 3068 2838 3080
rect 3786 3068 3792 3080
rect 3844 3108 3850 3120
rect 3973 3111 4031 3117
rect 3973 3108 3985 3111
rect 3844 3080 3985 3108
rect 3844 3068 3850 3080
rect 3973 3077 3985 3080
rect 4019 3077 4031 3111
rect 9861 3111 9919 3117
rect 9861 3108 9873 3111
rect 3973 3071 4031 3077
rect 7392 3080 9873 3108
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 3878 3040 3884 3052
rect 2363 3012 3884 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 3878 3000 3884 3012
rect 3936 3040 3942 3052
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 3936 3012 4353 3040
rect 3936 3000 3942 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 7392 3049 7420 3080
rect 9861 3077 9873 3080
rect 9907 3077 9919 3111
rect 11422 3108 11428 3120
rect 11383 3080 11428 3108
rect 9861 3071 9919 3077
rect 11422 3068 11428 3080
rect 11480 3108 11486 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 11480 3080 11805 3108
rect 11480 3068 11486 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 11793 3071 11851 3077
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 6972 3012 7205 3040
rect 6972 3000 6978 3012
rect 7193 3009 7205 3012
rect 7239 3040 7251 3043
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7239 3012 7389 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9306 3040 9312 3052
rect 9171 3012 9312 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10870 3040 10876 3052
rect 10735 3012 10876 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 4928 2975 4986 2981
rect 4928 2972 4940 2975
rect 4856 2944 4940 2972
rect 4856 2932 4862 2944
rect 4928 2941 4940 2944
rect 4974 2972 4986 2975
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 4974 2944 5365 2972
rect 4974 2941 4986 2944
rect 4928 2935 4986 2941
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2873 3479 2907
rect 5031 2907 5089 2913
rect 5031 2904 5043 2907
rect 3421 2867 3479 2873
rect 4126 2876 5043 2904
rect 3142 2836 3148 2848
rect 3103 2808 3148 2836
rect 3142 2796 3148 2808
rect 3200 2836 3206 2848
rect 3436 2836 3464 2867
rect 3200 2808 3464 2836
rect 3200 2796 3206 2808
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4126 2836 4154 2876
rect 5031 2873 5043 2876
rect 5077 2873 5089 2907
rect 8018 2904 8024 2916
rect 7979 2876 8024 2904
rect 5031 2867 5089 2873
rect 8018 2864 8024 2876
rect 8076 2864 8082 2916
rect 12176 2904 12204 3139
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 13872 3148 13917 3176
rect 13872 3136 13878 3148
rect 14090 3136 14096 3188
rect 14148 3176 14154 3188
rect 14185 3179 14243 3185
rect 14185 3176 14197 3179
rect 14148 3148 14197 3176
rect 14148 3136 14154 3148
rect 14185 3145 14197 3148
rect 14231 3145 14243 3179
rect 14185 3139 14243 3145
rect 15473 3179 15531 3185
rect 15473 3145 15485 3179
rect 15519 3176 15531 3179
rect 15746 3176 15752 3188
rect 15519 3148 15752 3176
rect 15519 3145 15531 3148
rect 15473 3139 15531 3145
rect 12342 3000 12348 3052
rect 12400 3040 12406 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12400 3012 12817 3040
rect 12400 3000 12406 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 14200 3040 14228 3139
rect 15746 3136 15752 3148
rect 15804 3136 15810 3188
rect 14461 3043 14519 3049
rect 14461 3040 14473 3043
rect 14200 3012 14473 3040
rect 12805 3003 12863 3009
rect 14461 3009 14473 3012
rect 14507 3009 14519 3043
rect 14461 3003 14519 3009
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14608 3012 14749 3040
rect 14608 3000 14614 3012
rect 14737 3009 14749 3012
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16025 3043 16083 3049
rect 16025 3040 16037 3043
rect 15887 3012 16037 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16025 3009 16037 3012
rect 16071 3040 16083 3043
rect 16298 3040 16304 3052
rect 16071 3012 16304 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 12529 2907 12587 2913
rect 12529 2904 12541 2907
rect 12176 2876 12541 2904
rect 12529 2873 12541 2876
rect 12575 2873 12587 2907
rect 12529 2867 12587 2873
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 13906 2904 13912 2916
rect 13504 2876 13912 2904
rect 13504 2864 13510 2876
rect 13906 2864 13912 2876
rect 13964 2904 13970 2916
rect 16669 2907 16727 2913
rect 16669 2904 16681 2907
rect 13964 2876 16681 2904
rect 13964 2864 13970 2876
rect 16669 2873 16681 2876
rect 16715 2873 16727 2907
rect 16669 2867 16727 2873
rect 3568 2808 4154 2836
rect 3568 2796 3574 2808
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7742 2836 7748 2848
rect 6972 2808 7748 2836
rect 6972 2796 6978 2808
rect 7742 2796 7748 2808
rect 7800 2836 7806 2848
rect 8297 2839 8355 2845
rect 8297 2836 8309 2839
rect 7800 2808 8309 2836
rect 7800 2796 7806 2808
rect 8297 2805 8309 2808
rect 8343 2805 8355 2839
rect 8297 2799 8355 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 18506 2836 18512 2848
rect 11112 2808 18512 2836
rect 11112 2796 11118 2808
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 1104 2746 17756 2768
rect 1104 2694 7288 2746
rect 7340 2694 7352 2746
rect 7404 2694 7416 2746
rect 7468 2694 7480 2746
rect 7532 2694 13595 2746
rect 13647 2694 13659 2746
rect 13711 2694 13723 2746
rect 13775 2694 13787 2746
rect 13839 2694 17756 2746
rect 1104 2672 17756 2694
rect 1995 2635 2053 2641
rect 1995 2601 2007 2635
rect 2041 2632 2053 2635
rect 3142 2632 3148 2644
rect 2041 2604 3148 2632
rect 2041 2601 2053 2604
rect 1995 2595 2053 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 3510 2632 3516 2644
rect 3471 2604 3516 2632
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3786 2632 3792 2644
rect 3747 2604 3792 2632
rect 3786 2592 3792 2604
rect 3844 2632 3850 2644
rect 5951 2635 6009 2641
rect 3844 2604 4200 2632
rect 3844 2592 3850 2604
rect 1924 2499 1982 2505
rect 1924 2465 1936 2499
rect 1970 2496 1982 2499
rect 2869 2499 2927 2505
rect 1970 2468 2452 2496
rect 1970 2465 1982 2468
rect 1924 2459 1982 2465
rect 2424 2301 2452 2468
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3528 2496 3556 2592
rect 4172 2573 4200 2604
rect 5951 2601 5963 2635
rect 5997 2632 6009 2635
rect 6914 2632 6920 2644
rect 5997 2604 6920 2632
rect 5997 2601 6009 2604
rect 5951 2595 6009 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 7064 2604 7113 2632
rect 7064 2592 7070 2604
rect 7101 2601 7113 2604
rect 7147 2632 7159 2635
rect 10505 2635 10563 2641
rect 7147 2604 7420 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2533 4215 2567
rect 4798 2564 4804 2576
rect 4759 2536 4804 2564
rect 4157 2527 4215 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7392 2573 7420 2604
rect 10505 2601 10517 2635
rect 10551 2632 10563 2635
rect 12158 2632 12164 2644
rect 10551 2604 12164 2632
rect 10551 2601 10563 2604
rect 10505 2595 10563 2601
rect 12158 2592 12164 2604
rect 12216 2592 12222 2644
rect 12434 2632 12440 2644
rect 12395 2604 12440 2632
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 15286 2592 15292 2644
rect 15344 2632 15350 2644
rect 15749 2635 15807 2641
rect 15749 2632 15761 2635
rect 15344 2604 15761 2632
rect 15344 2592 15350 2604
rect 15749 2601 15761 2604
rect 15795 2601 15807 2635
rect 15749 2595 15807 2601
rect 7377 2567 7435 2573
rect 7377 2533 7389 2567
rect 7423 2533 7435 2567
rect 8018 2564 8024 2576
rect 7979 2536 8024 2564
rect 7377 2527 7435 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 10962 2564 10968 2576
rect 10336 2536 10968 2564
rect 2915 2468 3556 2496
rect 5880 2499 5938 2505
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 5880 2465 5892 2499
rect 5926 2496 5938 2499
rect 5926 2468 6408 2496
rect 5926 2465 5938 2468
rect 5880 2459 5938 2465
rect 6380 2437 6408 2468
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2428 6423 2431
rect 8036 2428 8064 2524
rect 10336 2505 10364 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 12452 2564 12480 2592
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 12452 2536 13001 2564
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 12989 2527 13047 2533
rect 13633 2567 13691 2573
rect 13633 2533 13645 2567
rect 13679 2564 13691 2567
rect 13906 2564 13912 2576
rect 13679 2536 13912 2564
rect 13679 2533 13691 2536
rect 13633 2527 13691 2533
rect 13906 2524 13912 2536
rect 13964 2524 13970 2576
rect 15764 2564 15792 2595
rect 16025 2567 16083 2573
rect 16025 2564 16037 2567
rect 15764 2536 16037 2564
rect 16025 2533 16037 2536
rect 16071 2533 16083 2567
rect 16025 2527 16083 2533
rect 10321 2499 10379 2505
rect 10321 2465 10333 2499
rect 10367 2465 10379 2499
rect 10321 2459 10379 2465
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 11425 2499 11483 2505
rect 11425 2496 11437 2499
rect 11388 2468 11437 2496
rect 11388 2456 11394 2468
rect 11425 2465 11437 2468
rect 11471 2496 11483 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11471 2468 11989 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 16298 2428 16304 2440
rect 6411 2400 8064 2428
rect 16259 2400 16304 2428
rect 6411 2397 6423 2400
rect 6365 2391 6423 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 3053 2363 3111 2369
rect 3053 2329 3065 2363
rect 3099 2360 3111 2363
rect 4522 2360 4528 2372
rect 3099 2332 4528 2360
rect 3099 2329 3111 2332
rect 3053 2323 3111 2329
rect 4522 2320 4528 2332
rect 4580 2320 4586 2372
rect 11609 2363 11667 2369
rect 11609 2329 11621 2363
rect 11655 2360 11667 2363
rect 13078 2360 13084 2372
rect 11655 2332 13084 2360
rect 11655 2329 11667 2332
rect 11609 2323 11667 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 2409 2295 2467 2301
rect 2409 2261 2421 2295
rect 2455 2292 2467 2295
rect 2682 2292 2688 2304
rect 2455 2264 2688 2292
rect 2455 2261 2467 2264
rect 2409 2255 2467 2261
rect 2682 2252 2688 2264
rect 2740 2252 2746 2304
rect 1104 2202 17756 2224
rect 1104 2150 4135 2202
rect 4187 2150 4199 2202
rect 4251 2150 4263 2202
rect 4315 2150 4327 2202
rect 4379 2150 10441 2202
rect 10493 2150 10505 2202
rect 10557 2150 10569 2202
rect 10621 2150 10633 2202
rect 10685 2150 16748 2202
rect 16800 2150 16812 2202
rect 16864 2150 16876 2202
rect 16928 2150 16940 2202
rect 16992 2150 17756 2202
rect 1104 2128 17756 2150
rect 1486 76 1492 128
rect 1544 116 1550 128
rect 2406 116 2412 128
rect 1544 88 2412 116
rect 1544 76 1550 88
rect 2406 76 2412 88
rect 2464 76 2470 128
<< via1 >>
rect 12440 20544 12492 20596
rect 13176 20544 13228 20596
rect 4135 18470 4187 18522
rect 4199 18470 4251 18522
rect 4263 18470 4315 18522
rect 4327 18470 4379 18522
rect 10441 18470 10493 18522
rect 10505 18470 10557 18522
rect 10569 18470 10621 18522
rect 10633 18470 10685 18522
rect 16748 18470 16800 18522
rect 16812 18470 16864 18522
rect 16876 18470 16928 18522
rect 16940 18470 16992 18522
rect 14188 18411 14240 18420
rect 14188 18377 14197 18411
rect 14197 18377 14231 18411
rect 14231 18377 14240 18411
rect 14188 18368 14240 18377
rect 18236 18368 18288 18420
rect 7472 18275 7524 18284
rect 4896 18164 4948 18216
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 18420 18300 18472 18352
rect 17040 18232 17092 18284
rect 9404 18164 9456 18216
rect 14188 18164 14240 18216
rect 8944 18096 8996 18148
rect 18512 18096 18564 18148
rect 5540 18028 5592 18080
rect 5632 18028 5684 18080
rect 6276 18028 6328 18080
rect 8116 18028 8168 18080
rect 9772 18028 9824 18080
rect 13912 18028 13964 18080
rect 16028 18028 16080 18080
rect 7288 17926 7340 17978
rect 7352 17926 7404 17978
rect 7416 17926 7468 17978
rect 7480 17926 7532 17978
rect 13595 17926 13647 17978
rect 13659 17926 13711 17978
rect 13723 17926 13775 17978
rect 13787 17926 13839 17978
rect 1216 17756 1268 17808
rect 5632 17799 5684 17808
rect 5632 17765 5641 17799
rect 5641 17765 5675 17799
rect 5675 17765 5684 17799
rect 5632 17756 5684 17765
rect 8392 17756 8444 17808
rect 4436 17688 4488 17740
rect 11888 17688 11940 17740
rect 12624 17688 12676 17740
rect 14188 17688 14240 17740
rect 4804 17620 4856 17672
rect 7656 17620 7708 17672
rect 15752 17620 15804 17672
rect 15660 17552 15712 17604
rect 1860 17484 1912 17536
rect 3976 17484 4028 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 9128 17484 9180 17536
rect 10324 17484 10376 17536
rect 12992 17484 13044 17536
rect 4135 17382 4187 17434
rect 4199 17382 4251 17434
rect 4263 17382 4315 17434
rect 4327 17382 4379 17434
rect 10441 17382 10493 17434
rect 10505 17382 10557 17434
rect 10569 17382 10621 17434
rect 10633 17382 10685 17434
rect 16748 17382 16800 17434
rect 16812 17382 16864 17434
rect 16876 17382 16928 17434
rect 16940 17382 16992 17434
rect 1216 17280 1268 17332
rect 4436 17280 4488 17332
rect 5632 17280 5684 17332
rect 5816 17323 5868 17332
rect 5816 17289 5825 17323
rect 5825 17289 5859 17323
rect 5859 17289 5868 17323
rect 5816 17280 5868 17289
rect 10232 17280 10284 17332
rect 11888 17280 11940 17332
rect 12624 17323 12676 17332
rect 12624 17289 12633 17323
rect 12633 17289 12667 17323
rect 12667 17289 12676 17323
rect 12624 17280 12676 17289
rect 12992 17323 13044 17332
rect 12992 17289 13001 17323
rect 13001 17289 13035 17323
rect 13035 17289 13044 17323
rect 12992 17280 13044 17289
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 15752 17323 15804 17332
rect 15752 17289 15761 17323
rect 15761 17289 15795 17323
rect 15795 17289 15804 17323
rect 15752 17280 15804 17289
rect 1860 17187 1912 17196
rect 1860 17153 1869 17187
rect 1869 17153 1903 17187
rect 1903 17153 1912 17187
rect 1860 17144 1912 17153
rect 3976 17144 4028 17196
rect 4804 17187 4856 17196
rect 4804 17153 4813 17187
rect 4813 17153 4847 17187
rect 4847 17153 4856 17187
rect 4804 17144 4856 17153
rect 8024 17144 8076 17196
rect 8484 17144 8536 17196
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10600 17187 10652 17196
rect 10600 17153 10609 17187
rect 10609 17153 10643 17187
rect 10643 17153 10652 17187
rect 10600 17144 10652 17153
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 16120 17144 16172 17196
rect 5540 17076 5592 17128
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 2504 17051 2556 17060
rect 2504 17017 2513 17051
rect 2513 17017 2547 17051
rect 2547 17017 2556 17051
rect 2504 17008 2556 17017
rect 8392 17008 8444 17060
rect 14004 17008 14056 17060
rect 15476 17051 15528 17060
rect 15476 17017 15485 17051
rect 15485 17017 15519 17051
rect 15519 17017 15528 17051
rect 15476 17008 15528 17017
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 15292 16940 15344 16992
rect 7288 16838 7340 16890
rect 7352 16838 7404 16890
rect 7416 16838 7468 16890
rect 7480 16838 7532 16890
rect 13595 16838 13647 16890
rect 13659 16838 13711 16890
rect 13723 16838 13775 16890
rect 13787 16838 13839 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 16028 16736 16080 16788
rect 2504 16711 2556 16720
rect 2504 16677 2513 16711
rect 2513 16677 2547 16711
rect 2547 16677 2556 16711
rect 2504 16668 2556 16677
rect 4896 16711 4948 16720
rect 4896 16677 4905 16711
rect 4905 16677 4939 16711
rect 4939 16677 4948 16711
rect 4896 16668 4948 16677
rect 6276 16668 6328 16720
rect 8116 16711 8168 16720
rect 8116 16677 8125 16711
rect 8125 16677 8159 16711
rect 8159 16677 8168 16711
rect 8116 16668 8168 16677
rect 9772 16711 9824 16720
rect 9772 16677 9781 16711
rect 9781 16677 9815 16711
rect 9815 16677 9824 16711
rect 9772 16668 9824 16677
rect 9864 16668 9916 16720
rect 10600 16668 10652 16720
rect 13912 16668 13964 16720
rect 1584 16600 1636 16652
rect 4436 16532 4488 16584
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 8392 16575 8444 16584
rect 8392 16541 8401 16575
rect 8401 16541 8435 16575
rect 8435 16541 8444 16575
rect 8392 16532 8444 16541
rect 14004 16575 14056 16584
rect 14004 16541 14013 16575
rect 14013 16541 14047 16575
rect 14047 16541 14056 16575
rect 14004 16532 14056 16541
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 8024 16464 8076 16516
rect 2044 16396 2096 16448
rect 2136 16396 2188 16448
rect 4135 16294 4187 16346
rect 4199 16294 4251 16346
rect 4263 16294 4315 16346
rect 4327 16294 4379 16346
rect 10441 16294 10493 16346
rect 10505 16294 10557 16346
rect 10569 16294 10621 16346
rect 10633 16294 10685 16346
rect 16748 16294 16800 16346
rect 16812 16294 16864 16346
rect 16876 16294 16928 16346
rect 16940 16294 16992 16346
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 7656 16235 7708 16244
rect 7656 16201 7665 16235
rect 7665 16201 7699 16235
rect 7699 16201 7708 16235
rect 7656 16192 7708 16201
rect 2504 16099 2556 16108
rect 2504 16065 2513 16099
rect 2513 16065 2547 16099
rect 2547 16065 2556 16099
rect 2504 16056 2556 16065
rect 3608 16056 3660 16108
rect 4252 16056 4304 16108
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 8116 16192 8168 16244
rect 9772 16192 9824 16244
rect 13912 16192 13964 16244
rect 14004 16192 14056 16244
rect 8024 16056 8076 16108
rect 9864 16056 9916 16108
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 2136 15963 2188 15972
rect 2136 15929 2145 15963
rect 2145 15929 2179 15963
rect 2179 15929 2188 15963
rect 2136 15920 2188 15929
rect 4252 15963 4304 15972
rect 4252 15929 4261 15963
rect 4261 15929 4295 15963
rect 4295 15929 4304 15963
rect 4252 15920 4304 15929
rect 6276 15920 6328 15972
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 3608 15895 3660 15904
rect 3608 15861 3617 15895
rect 3617 15861 3651 15895
rect 3651 15861 3660 15895
rect 3608 15852 3660 15861
rect 4436 15852 4488 15904
rect 7288 15750 7340 15802
rect 7352 15750 7404 15802
rect 7416 15750 7468 15802
rect 7480 15750 7532 15802
rect 13595 15750 13647 15802
rect 13659 15750 13711 15802
rect 13723 15750 13775 15802
rect 13787 15750 13839 15802
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 2044 15580 2096 15632
rect 3608 15580 3660 15632
rect 8392 15580 8444 15632
rect 15292 15580 15344 15632
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6552 15444 6604 15496
rect 9956 15444 10008 15496
rect 15660 15444 15712 15496
rect 8668 15419 8720 15428
rect 8668 15385 8677 15419
rect 8677 15385 8711 15419
rect 8711 15385 8720 15419
rect 8668 15376 8720 15385
rect 4135 15206 4187 15258
rect 4199 15206 4251 15258
rect 4263 15206 4315 15258
rect 4327 15206 4379 15258
rect 10441 15206 10493 15258
rect 10505 15206 10557 15258
rect 10569 15206 10621 15258
rect 10633 15206 10685 15258
rect 16748 15206 16800 15258
rect 16812 15206 16864 15258
rect 16876 15206 16928 15258
rect 16940 15206 16992 15258
rect 2136 15104 2188 15156
rect 6092 15147 6144 15156
rect 6092 15113 6101 15147
rect 6101 15113 6135 15147
rect 6135 15113 6144 15147
rect 6092 15104 6144 15113
rect 6552 15147 6604 15156
rect 6552 15113 6561 15147
rect 6561 15113 6595 15147
rect 6595 15113 6604 15147
rect 6552 15104 6604 15113
rect 7104 15104 7156 15156
rect 8392 15104 8444 15156
rect 15292 15104 15344 15156
rect 6828 15036 6880 15088
rect 2044 14968 2096 15020
rect 1676 14900 1728 14952
rect 1492 14832 1544 14884
rect 6552 14900 6604 14952
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 16304 15011 16356 15020
rect 16304 14977 16313 15011
rect 16313 14977 16347 15011
rect 16347 14977 16356 15011
rect 16304 14968 16356 14977
rect 112 14764 164 14816
rect 3056 14764 3108 14816
rect 5632 14764 5684 14816
rect 7932 14832 7984 14884
rect 8944 14764 8996 14816
rect 16212 14764 16264 14816
rect 7288 14662 7340 14714
rect 7352 14662 7404 14714
rect 7416 14662 7468 14714
rect 7480 14662 7532 14714
rect 13595 14662 13647 14714
rect 13659 14662 13711 14714
rect 13723 14662 13775 14714
rect 13787 14662 13839 14714
rect 3056 14492 3108 14544
rect 4804 14560 4856 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 16120 14492 16172 14544
rect 5632 14424 5684 14476
rect 8668 14424 8720 14476
rect 9680 14467 9732 14476
rect 9680 14433 9724 14467
rect 9724 14433 9732 14467
rect 9680 14424 9732 14433
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 4528 14399 4580 14408
rect 4528 14365 4537 14399
rect 4537 14365 4571 14399
rect 4571 14365 4580 14399
rect 4528 14356 4580 14365
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 1676 14263 1728 14272
rect 1676 14229 1685 14263
rect 1685 14229 1719 14263
rect 1719 14229 1728 14263
rect 1676 14220 1728 14229
rect 5080 14220 5132 14272
rect 9312 14220 9364 14272
rect 4135 14118 4187 14170
rect 4199 14118 4251 14170
rect 4263 14118 4315 14170
rect 4327 14118 4379 14170
rect 10441 14118 10493 14170
rect 10505 14118 10557 14170
rect 10569 14118 10621 14170
rect 10633 14118 10685 14170
rect 16748 14118 16800 14170
rect 16812 14118 16864 14170
rect 16876 14118 16928 14170
rect 16940 14118 16992 14170
rect 3056 14016 3108 14068
rect 4804 14059 4856 14068
rect 4804 14025 4813 14059
rect 4813 14025 4847 14059
rect 4847 14025 4856 14059
rect 4804 14016 4856 14025
rect 5632 14016 5684 14068
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 9680 14059 9732 14068
rect 9680 14025 9689 14059
rect 9689 14025 9723 14059
rect 9723 14025 9732 14059
rect 9680 14016 9732 14025
rect 16120 14016 16172 14068
rect 16488 14059 16540 14068
rect 16488 14025 16497 14059
rect 16497 14025 16531 14059
rect 16531 14025 16540 14059
rect 16488 14016 16540 14025
rect 2320 13991 2372 14000
rect 2320 13957 2329 13991
rect 2329 13957 2363 13991
rect 2363 13957 2372 13991
rect 2320 13948 2372 13957
rect 1952 13880 2004 13932
rect 4528 13923 4580 13932
rect 4528 13889 4537 13923
rect 4537 13889 4571 13923
rect 4571 13889 4580 13923
rect 4528 13880 4580 13889
rect 9312 13812 9364 13864
rect 16212 13812 16264 13864
rect 3884 13787 3936 13796
rect 3884 13753 3893 13787
rect 3893 13753 3927 13787
rect 3927 13753 3936 13787
rect 3884 13744 3936 13753
rect 9036 13676 9088 13728
rect 14648 13719 14700 13728
rect 14648 13685 14657 13719
rect 14657 13685 14691 13719
rect 14691 13685 14700 13719
rect 14648 13676 14700 13685
rect 7288 13574 7340 13626
rect 7352 13574 7404 13626
rect 7416 13574 7468 13626
rect 7480 13574 7532 13626
rect 13595 13574 13647 13626
rect 13659 13574 13711 13626
rect 13723 13574 13775 13626
rect 13787 13574 13839 13626
rect 1952 13472 2004 13524
rect 2044 13447 2096 13456
rect 2044 13413 2053 13447
rect 2053 13413 2087 13447
rect 2087 13413 2096 13447
rect 2044 13404 2096 13413
rect 2688 13404 2740 13456
rect 14648 13404 14700 13456
rect 15752 13404 15804 13456
rect 16028 13447 16080 13456
rect 16028 13413 16037 13447
rect 16037 13413 16071 13447
rect 16071 13413 16080 13447
rect 16028 13404 16080 13413
rect 4528 13336 4580 13388
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 3240 13132 3292 13184
rect 4135 13030 4187 13082
rect 4199 13030 4251 13082
rect 4263 13030 4315 13082
rect 4327 13030 4379 13082
rect 10441 13030 10493 13082
rect 10505 13030 10557 13082
rect 10569 13030 10621 13082
rect 10633 13030 10685 13082
rect 16748 13030 16800 13082
rect 16812 13030 16864 13082
rect 16876 13030 16928 13082
rect 16940 13030 16992 13082
rect 1676 12928 1728 12980
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 4528 12928 4580 12980
rect 15752 12971 15804 12980
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 16028 12928 16080 12980
rect 112 12860 164 12912
rect 3884 12792 3936 12844
rect 17132 12860 17184 12912
rect 2320 12724 2372 12776
rect 3240 12724 3292 12776
rect 7288 12486 7340 12538
rect 7352 12486 7404 12538
rect 7416 12486 7468 12538
rect 7480 12486 7532 12538
rect 13595 12486 13647 12538
rect 13659 12486 13711 12538
rect 13723 12486 13775 12538
rect 13787 12486 13839 12538
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 4135 11942 4187 11994
rect 4199 11942 4251 11994
rect 4263 11942 4315 11994
rect 4327 11942 4379 11994
rect 10441 11942 10493 11994
rect 10505 11942 10557 11994
rect 10569 11942 10621 11994
rect 10633 11942 10685 11994
rect 16748 11942 16800 11994
rect 16812 11942 16864 11994
rect 16876 11942 16928 11994
rect 16940 11942 16992 11994
rect 1676 11840 1728 11892
rect 1676 11636 1728 11688
rect 7288 11398 7340 11450
rect 7352 11398 7404 11450
rect 7416 11398 7468 11450
rect 7480 11398 7532 11450
rect 13595 11398 13647 11450
rect 13659 11398 13711 11450
rect 13723 11398 13775 11450
rect 13787 11398 13839 11450
rect 4620 11160 4672 11212
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 16120 11092 16172 11144
rect 3608 10956 3660 11008
rect 4135 10854 4187 10906
rect 4199 10854 4251 10906
rect 4263 10854 4315 10906
rect 4327 10854 4379 10906
rect 10441 10854 10493 10906
rect 10505 10854 10557 10906
rect 10569 10854 10621 10906
rect 10633 10854 10685 10906
rect 16748 10854 16800 10906
rect 16812 10854 16864 10906
rect 16876 10854 16928 10906
rect 16940 10854 16992 10906
rect 4620 10795 4672 10804
rect 4620 10761 4629 10795
rect 4629 10761 4663 10795
rect 4663 10761 4672 10795
rect 4620 10752 4672 10761
rect 16028 10752 16080 10804
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 3792 10616 3844 10668
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 112 10548 164 10600
rect 1584 10548 1636 10600
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 2780 10480 2832 10532
rect 1584 10412 1636 10421
rect 7288 10310 7340 10362
rect 7352 10310 7404 10362
rect 7416 10310 7468 10362
rect 7480 10310 7532 10362
rect 13595 10310 13647 10362
rect 13659 10310 13711 10362
rect 13723 10310 13775 10362
rect 13787 10310 13839 10362
rect 16028 10208 16080 10260
rect 2044 10072 2096 10124
rect 15384 10115 15436 10124
rect 15384 10081 15402 10115
rect 15402 10081 15436 10115
rect 15384 10072 15436 10081
rect 15936 10072 15988 10124
rect 17040 10072 17092 10124
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 1492 9868 1544 9920
rect 16120 9868 16172 9920
rect 4135 9766 4187 9818
rect 4199 9766 4251 9818
rect 4263 9766 4315 9818
rect 4327 9766 4379 9818
rect 10441 9766 10493 9818
rect 10505 9766 10557 9818
rect 10569 9766 10621 9818
rect 10633 9766 10685 9818
rect 16748 9766 16800 9818
rect 16812 9766 16864 9818
rect 16876 9766 16928 9818
rect 16940 9766 16992 9818
rect 1308 9664 1360 9716
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 2780 9664 2832 9716
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 3792 9571 3844 9580
rect 2504 9528 2556 9537
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 1492 9460 1544 9512
rect 12440 9664 12492 9716
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 16120 9707 16172 9716
rect 16120 9673 16129 9707
rect 16129 9673 16163 9707
rect 16163 9673 16172 9707
rect 16120 9664 16172 9673
rect 18420 9596 18472 9648
rect 16120 9460 16172 9512
rect 2964 9435 3016 9444
rect 2964 9401 2973 9435
rect 2973 9401 3007 9435
rect 3007 9401 3016 9435
rect 2964 9392 3016 9401
rect 6368 9324 6420 9376
rect 17040 9324 17092 9376
rect 7288 9222 7340 9274
rect 7352 9222 7404 9274
rect 7416 9222 7468 9274
rect 7480 9222 7532 9274
rect 13595 9222 13647 9274
rect 13659 9222 13711 9274
rect 13723 9222 13775 9274
rect 13787 9222 13839 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 2964 9120 3016 9172
rect 16488 9163 16540 9172
rect 16488 9129 16497 9163
rect 16497 9129 16531 9163
rect 16531 9129 16540 9163
rect 16488 9120 16540 9129
rect 6368 9095 6420 9104
rect 6368 9061 6377 9095
rect 6377 9061 6411 9095
rect 6411 9061 6420 9095
rect 6368 9052 6420 9061
rect 15200 9027 15252 9036
rect 15200 8993 15209 9027
rect 15209 8993 15243 9027
rect 15243 8993 15252 9027
rect 15200 8984 15252 8993
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 5908 8916 5960 8968
rect 2596 8823 2648 8832
rect 2596 8789 2605 8823
rect 2605 8789 2639 8823
rect 2639 8789 2648 8823
rect 2596 8780 2648 8789
rect 4135 8678 4187 8730
rect 4199 8678 4251 8730
rect 4263 8678 4315 8730
rect 4327 8678 4379 8730
rect 10441 8678 10493 8730
rect 10505 8678 10557 8730
rect 10569 8678 10621 8730
rect 10633 8678 10685 8730
rect 16748 8678 16800 8730
rect 16812 8678 16864 8730
rect 16876 8678 16928 8730
rect 16940 8678 16992 8730
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 15200 8576 15252 8628
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 16304 8576 16356 8628
rect 16396 8440 16448 8492
rect 2596 8236 2648 8288
rect 3240 8236 3292 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 7288 8134 7340 8186
rect 7352 8134 7404 8186
rect 7416 8134 7468 8186
rect 7480 8134 7532 8186
rect 13595 8134 13647 8186
rect 13659 8134 13711 8186
rect 13723 8134 13775 8186
rect 13787 8134 13839 8186
rect 4988 8032 5040 8084
rect 5908 7964 5960 8016
rect 6368 8007 6420 8016
rect 6368 7973 6377 8007
rect 6377 7973 6411 8007
rect 6411 7973 6420 8007
rect 6368 7964 6420 7973
rect 4436 7939 4488 7948
rect 4436 7905 4445 7939
rect 4445 7905 4479 7939
rect 4479 7905 4488 7939
rect 4436 7896 4488 7905
rect 14832 7896 14884 7948
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 16304 7828 16356 7880
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 15384 7692 15436 7744
rect 4135 7590 4187 7642
rect 4199 7590 4251 7642
rect 4263 7590 4315 7642
rect 4327 7590 4379 7642
rect 10441 7590 10493 7642
rect 10505 7590 10557 7642
rect 10569 7590 10621 7642
rect 10633 7590 10685 7642
rect 16748 7590 16800 7642
rect 16812 7590 16864 7642
rect 16876 7590 16928 7642
rect 16940 7590 16992 7642
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 14464 7531 14516 7540
rect 14464 7497 14473 7531
rect 14473 7497 14507 7531
rect 14507 7497 14516 7531
rect 14464 7488 14516 7497
rect 14832 7531 14884 7540
rect 14832 7497 14841 7531
rect 14841 7497 14875 7531
rect 14875 7497 14884 7531
rect 14832 7488 14884 7497
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 14464 7284 14516 7336
rect 15476 7284 15528 7336
rect 14832 7216 14884 7268
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 7288 7046 7340 7098
rect 7352 7046 7404 7098
rect 7416 7046 7468 7098
rect 7480 7046 7532 7098
rect 13595 7046 13647 7098
rect 13659 7046 13711 7098
rect 13723 7046 13775 7098
rect 13787 7046 13839 7098
rect 6368 6919 6420 6928
rect 6368 6885 6377 6919
rect 6377 6885 6411 6919
rect 6411 6885 6420 6919
rect 6368 6876 6420 6885
rect 6828 6876 6880 6928
rect 7012 6919 7064 6928
rect 7012 6885 7021 6919
rect 7021 6885 7055 6919
rect 7055 6885 7064 6919
rect 7012 6876 7064 6885
rect 7840 6851 7892 6860
rect 7840 6817 7884 6851
rect 7884 6817 7892 6851
rect 7840 6808 7892 6817
rect 13452 6808 13504 6860
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 14464 6672 14516 6724
rect 7472 6604 7524 6656
rect 10968 6604 11020 6656
rect 15292 6604 15344 6656
rect 4135 6502 4187 6554
rect 4199 6502 4251 6554
rect 4263 6502 4315 6554
rect 4327 6502 4379 6554
rect 10441 6502 10493 6554
rect 10505 6502 10557 6554
rect 10569 6502 10621 6554
rect 10633 6502 10685 6554
rect 16748 6502 16800 6554
rect 16812 6502 16864 6554
rect 16876 6502 16928 6554
rect 16940 6502 16992 6554
rect 6368 6443 6420 6452
rect 6368 6409 6377 6443
rect 6377 6409 6411 6443
rect 6411 6409 6420 6443
rect 6368 6400 6420 6409
rect 7472 6443 7524 6452
rect 7472 6409 7481 6443
rect 7481 6409 7515 6443
rect 7515 6409 7524 6443
rect 7472 6400 7524 6409
rect 7840 6443 7892 6452
rect 7840 6409 7849 6443
rect 7849 6409 7883 6443
rect 7883 6409 7892 6443
rect 7840 6400 7892 6409
rect 15936 6400 15988 6452
rect 7472 6196 7524 6248
rect 14556 6264 14608 6316
rect 17132 6332 17184 6384
rect 14464 6128 14516 6180
rect 17224 6264 17276 6316
rect 7104 6060 7156 6112
rect 12992 6060 13044 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 13912 6060 13964 6112
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 15016 6060 15068 6112
rect 16212 6103 16264 6112
rect 16212 6069 16221 6103
rect 16221 6069 16255 6103
rect 16255 6069 16264 6103
rect 16212 6060 16264 6069
rect 7288 5958 7340 6010
rect 7352 5958 7404 6010
rect 7416 5958 7468 6010
rect 7480 5958 7532 6010
rect 13595 5958 13647 6010
rect 13659 5958 13711 6010
rect 13723 5958 13775 6010
rect 13787 5958 13839 6010
rect 15384 5831 15436 5840
rect 15384 5797 15393 5831
rect 15393 5797 15427 5831
rect 15427 5797 15436 5831
rect 15384 5788 15436 5797
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 4135 5414 4187 5466
rect 4199 5414 4251 5466
rect 4263 5414 4315 5466
rect 4327 5414 4379 5466
rect 10441 5414 10493 5466
rect 10505 5414 10557 5466
rect 10569 5414 10621 5466
rect 10633 5414 10685 5466
rect 16748 5414 16800 5466
rect 16812 5414 16864 5466
rect 16876 5414 16928 5466
rect 16940 5414 16992 5466
rect 15016 5312 15068 5364
rect 15384 5287 15436 5296
rect 15384 5253 15393 5287
rect 15393 5253 15427 5287
rect 15427 5253 15436 5287
rect 15384 5244 15436 5253
rect 9312 4972 9364 5024
rect 15476 5176 15528 5228
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 12716 5040 12768 5092
rect 14004 5040 14056 5092
rect 14280 5083 14332 5092
rect 14280 5049 14289 5083
rect 14289 5049 14323 5083
rect 14323 5049 14332 5083
rect 14280 5040 14332 5049
rect 11244 4972 11296 5024
rect 12440 4972 12492 5024
rect 7288 4870 7340 4922
rect 7352 4870 7404 4922
rect 7416 4870 7468 4922
rect 7480 4870 7532 4922
rect 13595 4870 13647 4922
rect 13659 4870 13711 4922
rect 13723 4870 13775 4922
rect 13787 4870 13839 4922
rect 12348 4811 12400 4820
rect 12348 4777 12357 4811
rect 12357 4777 12391 4811
rect 12391 4777 12400 4811
rect 12348 4768 12400 4777
rect 13912 4700 13964 4752
rect 14004 4700 14056 4752
rect 15660 4700 15712 4752
rect 10232 4632 10284 4684
rect 11152 4632 11204 4684
rect 12164 4675 12216 4684
rect 12164 4641 12173 4675
rect 12173 4641 12207 4675
rect 12207 4641 12216 4675
rect 12164 4632 12216 4641
rect 14832 4564 14884 4616
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 15752 4564 15804 4616
rect 10876 4428 10928 4480
rect 4135 4326 4187 4378
rect 4199 4326 4251 4378
rect 4263 4326 4315 4378
rect 4327 4326 4379 4378
rect 10441 4326 10493 4378
rect 10505 4326 10557 4378
rect 10569 4326 10621 4378
rect 10633 4326 10685 4378
rect 16748 4326 16800 4378
rect 16812 4326 16864 4378
rect 16876 4326 16928 4378
rect 16940 4326 16992 4378
rect 1860 4267 1912 4276
rect 1860 4233 1869 4267
rect 1869 4233 1903 4267
rect 1903 4233 1912 4267
rect 1860 4224 1912 4233
rect 12164 4267 12216 4276
rect 12164 4233 12173 4267
rect 12173 4233 12207 4267
rect 12207 4233 12216 4267
rect 12164 4224 12216 4233
rect 12532 4224 12584 4276
rect 13912 4267 13964 4276
rect 2872 4088 2924 4140
rect 1860 4020 1912 4072
rect 3976 4020 4028 4072
rect 10232 4088 10284 4140
rect 13912 4233 13921 4267
rect 13921 4233 13955 4267
rect 13955 4233 13964 4267
rect 13912 4224 13964 4233
rect 15568 4224 15620 4276
rect 12716 4156 12768 4208
rect 2136 3884 2188 3936
rect 6276 3884 6328 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 9588 3884 9640 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11060 3927 11112 3936
rect 11060 3893 11069 3927
rect 11069 3893 11103 3927
rect 11103 3893 11112 3927
rect 11060 3884 11112 3893
rect 11336 3884 11388 3936
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 14280 3952 14332 4004
rect 12348 3884 12400 3936
rect 7288 3782 7340 3834
rect 7352 3782 7404 3834
rect 7416 3782 7468 3834
rect 7480 3782 7532 3834
rect 13595 3782 13647 3834
rect 13659 3782 13711 3834
rect 13723 3782 13775 3834
rect 13787 3782 13839 3834
rect 2136 3655 2188 3664
rect 2136 3621 2145 3655
rect 2145 3621 2179 3655
rect 2179 3621 2188 3655
rect 2136 3612 2188 3621
rect 6276 3655 6328 3664
rect 6276 3621 6285 3655
rect 6285 3621 6319 3655
rect 6319 3621 6328 3655
rect 6276 3612 6328 3621
rect 9588 3612 9640 3664
rect 10232 3612 10284 3664
rect 15752 3612 15804 3664
rect 7748 3587 7800 3596
rect 7748 3553 7757 3587
rect 7757 3553 7791 3587
rect 7791 3553 7800 3587
rect 7748 3544 7800 3553
rect 12992 3544 13044 3596
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 3884 3476 3936 3528
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 11428 3476 11480 3528
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 14556 3476 14608 3528
rect 8208 3340 8260 3392
rect 14004 3383 14056 3392
rect 14004 3349 14013 3383
rect 14013 3349 14047 3383
rect 14047 3349 14056 3383
rect 14004 3340 14056 3349
rect 4135 3238 4187 3290
rect 4199 3238 4251 3290
rect 4263 3238 4315 3290
rect 4327 3238 4379 3290
rect 10441 3238 10493 3290
rect 10505 3238 10557 3290
rect 10569 3238 10621 3290
rect 10633 3238 10685 3290
rect 16748 3238 16800 3290
rect 16812 3238 16864 3290
rect 16876 3238 16928 3290
rect 16940 3238 16992 3290
rect 2136 3179 2188 3188
rect 2136 3145 2145 3179
rect 2145 3145 2179 3179
rect 2179 3145 2188 3179
rect 2136 3136 2188 3145
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 10232 3179 10284 3188
rect 10232 3145 10241 3179
rect 10241 3145 10275 3179
rect 10275 3145 10284 3179
rect 10232 3136 10284 3145
rect 10324 3136 10376 3188
rect 2780 3068 2832 3120
rect 3792 3068 3844 3120
rect 3884 3000 3936 3052
rect 6920 3000 6972 3052
rect 11428 3111 11480 3120
rect 11428 3077 11437 3111
rect 11437 3077 11471 3111
rect 11471 3077 11480 3111
rect 11428 3068 11480 3077
rect 9312 3043 9364 3052
rect 9312 3009 9321 3043
rect 9321 3009 9355 3043
rect 9355 3009 9364 3043
rect 9312 3000 9364 3009
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 4804 2932 4856 2984
rect 3148 2839 3200 2848
rect 3148 2805 3157 2839
rect 3157 2805 3191 2839
rect 3191 2805 3200 2839
rect 3148 2796 3200 2805
rect 3516 2796 3568 2848
rect 8024 2907 8076 2916
rect 8024 2873 8033 2907
rect 8033 2873 8067 2907
rect 8067 2873 8076 2907
rect 8024 2864 8076 2873
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14096 3136 14148 3188
rect 12348 3000 12400 3052
rect 15752 3136 15804 3188
rect 14556 3000 14608 3052
rect 16304 3000 16356 3052
rect 13452 2864 13504 2916
rect 13912 2864 13964 2916
rect 6920 2796 6972 2848
rect 7748 2796 7800 2848
rect 11060 2796 11112 2848
rect 18512 2796 18564 2848
rect 7288 2694 7340 2746
rect 7352 2694 7404 2746
rect 7416 2694 7468 2746
rect 7480 2694 7532 2746
rect 13595 2694 13647 2746
rect 13659 2694 13711 2746
rect 13723 2694 13775 2746
rect 13787 2694 13839 2746
rect 3148 2592 3200 2644
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 3792 2635 3844 2644
rect 3792 2601 3801 2635
rect 3801 2601 3835 2635
rect 3835 2601 3844 2635
rect 3792 2592 3844 2601
rect 6920 2592 6972 2644
rect 7012 2592 7064 2644
rect 4804 2567 4856 2576
rect 4804 2533 4813 2567
rect 4813 2533 4847 2567
rect 4847 2533 4856 2567
rect 4804 2524 4856 2533
rect 12164 2592 12216 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 15292 2592 15344 2644
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 10968 2567 11020 2576
rect 10968 2533 10977 2567
rect 10977 2533 11011 2567
rect 11011 2533 11020 2567
rect 10968 2524 11020 2533
rect 13912 2524 13964 2576
rect 11336 2456 11388 2508
rect 16304 2431 16356 2440
rect 16304 2397 16313 2431
rect 16313 2397 16347 2431
rect 16347 2397 16356 2431
rect 16304 2388 16356 2397
rect 4528 2320 4580 2372
rect 13084 2320 13136 2372
rect 2688 2252 2740 2304
rect 4135 2150 4187 2202
rect 4199 2150 4251 2202
rect 4263 2150 4315 2202
rect 4327 2150 4379 2202
rect 10441 2150 10493 2202
rect 10505 2150 10557 2202
rect 10569 2150 10621 2202
rect 10633 2150 10685 2202
rect 16748 2150 16800 2202
rect 16812 2150 16864 2202
rect 16876 2150 16928 2202
rect 16940 2150 16992 2202
rect 1492 76 1544 128
rect 2412 76 2464 128
<< metal2 >>
rect 570 20583 626 21063
rect 1766 20583 1822 21063
rect 3054 20618 3110 21063
rect 2884 20590 3110 20618
rect 1214 19544 1270 19553
rect 1214 19479 1270 19488
rect 1228 17814 1256 19479
rect 1216 17808 1268 17814
rect 1780 17785 1808 20583
rect 1216 17750 1268 17756
rect 1766 17776 1822 17785
rect 1228 17338 1256 17750
rect 1766 17711 1822 17720
rect 1766 17640 1822 17649
rect 1766 17575 1822 17584
rect 1216 17332 1268 17338
rect 1216 17274 1268 17280
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 15910 1624 16594
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1492 14884 1544 14890
rect 1492 14826 1544 14832
rect 112 14816 164 14822
rect 112 14758 164 14764
rect 124 14385 152 14758
rect 110 14376 166 14385
rect 110 14311 166 14320
rect 1504 13814 1532 14826
rect 1412 13786 1532 13814
rect 112 12912 164 12918
rect 112 12854 164 12860
rect 124 12481 152 12854
rect 110 12472 166 12481
rect 110 12407 166 12416
rect 112 10600 164 10606
rect 112 10542 164 10548
rect 124 6769 152 10542
rect 1306 10024 1362 10033
rect 1306 9959 1362 9968
rect 1320 9722 1348 9959
rect 1308 9716 1360 9722
rect 1308 9658 1360 9664
rect 110 6760 166 6769
rect 110 6695 166 6704
rect 1412 626 1440 13786
rect 1596 10606 1624 15846
rect 1676 14952 1728 14958
rect 1676 14894 1728 14900
rect 1688 14278 1716 14894
rect 1676 14272 1728 14278
rect 1676 14214 1728 14220
rect 1688 12986 1716 14214
rect 1780 13814 1808 17575
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1872 17202 1900 17478
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1872 16794 1900 17138
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 2516 16726 2544 17002
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 2056 15638 2084 16390
rect 2148 15978 2176 16390
rect 2516 16114 2544 16662
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2136 15972 2188 15978
rect 2136 15914 2188 15920
rect 2044 15632 2096 15638
rect 2044 15574 2096 15580
rect 2056 15026 2084 15574
rect 2148 15162 2176 15914
rect 2136 15156 2188 15162
rect 2136 15098 2188 15104
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1780 13786 1900 13814
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11898 1716 12174
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9518 1532 9862
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1596 9178 1624 10406
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1688 4049 1716 11630
rect 1872 4282 1900 13786
rect 1964 13530 1992 13874
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2044 13456 2096 13462
rect 2044 13398 2096 13404
rect 2056 12986 2084 13398
rect 2332 13326 2360 13942
rect 2700 13462 2728 14350
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2332 12986 2360 13262
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2056 12238 2084 12922
rect 2332 12782 2360 12922
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2056 9722 2084 10066
rect 2792 10062 2820 10474
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 2516 9586 2544 9998
rect 2792 9722 2820 9998
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8294 2636 8774
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1872 4078 1900 4218
rect 2884 4146 2912 20590
rect 3054 20583 3110 20590
rect 4342 20618 4398 21063
rect 5538 20618 5594 21063
rect 4342 20590 4476 20618
rect 4342 20583 4398 20590
rect 4109 18524 4405 18544
rect 4165 18522 4189 18524
rect 4245 18522 4269 18524
rect 4325 18522 4349 18524
rect 4187 18470 4189 18522
rect 4251 18470 4263 18522
rect 4325 18470 4327 18522
rect 4165 18468 4189 18470
rect 4245 18468 4269 18470
rect 4325 18468 4349 18470
rect 4109 18448 4405 18468
rect 4448 17746 4476 20590
rect 5538 20590 5856 20618
rect 5538 20583 5594 20590
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3988 17202 4016 17478
rect 4109 17436 4405 17456
rect 4165 17434 4189 17436
rect 4245 17434 4269 17436
rect 4325 17434 4349 17436
rect 4187 17382 4189 17434
rect 4251 17382 4263 17434
rect 4325 17382 4327 17434
rect 4165 17380 4189 17382
rect 4245 17380 4269 17382
rect 4325 17380 4349 17382
rect 4109 17360 4405 17380
rect 4448 17338 4476 17682
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4816 17202 4844 17614
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4109 16348 4405 16368
rect 4165 16346 4189 16348
rect 4245 16346 4269 16348
rect 4325 16346 4349 16348
rect 4187 16294 4189 16346
rect 4251 16294 4263 16346
rect 4325 16294 4327 16346
rect 4165 16292 4189 16294
rect 4245 16292 4269 16294
rect 4325 16292 4349 16294
rect 4109 16272 4405 16292
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 3620 15910 3648 16050
rect 4264 15978 4292 16050
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4448 15910 4476 16526
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 3620 15638 3648 15846
rect 3974 15736 4030 15745
rect 3974 15671 4030 15680
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 3068 14550 3096 14758
rect 3056 14544 3108 14550
rect 3056 14486 3108 14492
rect 3068 14074 3096 14486
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3884 13796 3936 13802
rect 3884 13738 3936 13744
rect 3240 13184 3292 13190
rect 3240 13126 3292 13132
rect 3252 12986 3280 13126
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3252 12782 3280 12922
rect 3896 12850 3924 13738
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10674 3648 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3804 9586 3832 10610
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 9178 3004 9386
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 1860 4072 1912 4078
rect 1674 4040 1730 4049
rect 1860 4014 1912 4020
rect 1674 3975 1730 3984
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3670 2176 3878
rect 2136 3664 2188 3670
rect 2136 3606 2188 3612
rect 2148 3194 2176 3606
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2792 3126 2820 3470
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3160 2650 3188 2790
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 1412 598 1532 626
rect 478 0 534 480
rect 1398 0 1454 480
rect 1504 134 1532 598
rect 1492 128 1544 134
rect 1492 70 1544 76
rect 2410 128 2466 480
rect 2410 76 2412 128
rect 2464 76 2466 128
rect 2700 105 2728 2246
rect 2410 0 2466 76
rect 2686 96 2742 105
rect 3252 82 3280 8230
rect 3988 4078 4016 15671
rect 4109 15260 4405 15280
rect 4165 15258 4189 15260
rect 4245 15258 4269 15260
rect 4325 15258 4349 15260
rect 4187 15206 4189 15258
rect 4251 15206 4263 15258
rect 4325 15206 4327 15258
rect 4165 15204 4189 15206
rect 4245 15204 4269 15206
rect 4325 15204 4349 15206
rect 4109 15184 4405 15204
rect 4816 14618 4844 17138
rect 4908 16726 4936 18158
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5552 17134 5580 18022
rect 5644 17814 5672 18022
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5644 17338 5672 17750
rect 5828 17338 5856 20590
rect 6826 20583 6882 21063
rect 8114 20618 8170 21063
rect 8114 20590 8432 20618
rect 8114 20583 8170 20590
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 5816 17332 5868 17338
rect 5816 17274 5868 17280
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 6288 16726 6316 18022
rect 4896 16720 4948 16726
rect 6276 16720 6328 16726
rect 4896 16662 4948 16668
rect 6196 16680 6276 16708
rect 4908 16114 4936 16662
rect 6196 16250 6224 16680
rect 6276 16662 6328 16668
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 6288 15978 6316 16526
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6104 15162 6132 15438
rect 6564 15162 6592 15438
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6564 14958 6592 15098
rect 6840 15094 6868 20583
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 18193 7512 18226
rect 7470 18184 7526 18193
rect 7470 18119 7526 18128
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7262 17980 7558 18000
rect 7318 17978 7342 17980
rect 7398 17978 7422 17980
rect 7478 17978 7502 17980
rect 7340 17926 7342 17978
rect 7404 17926 7416 17978
rect 7478 17926 7480 17978
rect 7318 17924 7342 17926
rect 7398 17924 7422 17926
rect 7478 17924 7502 17926
rect 7262 17904 7558 17924
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 15162 7144 16934
rect 7262 16892 7558 16912
rect 7318 16890 7342 16892
rect 7398 16890 7422 16892
rect 7478 16890 7502 16892
rect 7340 16838 7342 16890
rect 7404 16838 7416 16890
rect 7478 16838 7480 16890
rect 7318 16836 7342 16838
rect 7398 16836 7422 16838
rect 7478 16836 7502 16838
rect 7262 16816 7558 16836
rect 7668 16250 7696 17614
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 16522 8064 17138
rect 8128 16726 8156 18022
rect 8404 17814 8432 20590
rect 9402 20583 9458 21063
rect 10598 20618 10654 21063
rect 10244 20590 10654 20618
rect 9416 18222 9444 20583
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 17202 8524 17478
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8392 17060 8444 17066
rect 8392 17002 8444 17008
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 8036 16114 8064 16458
rect 8128 16250 8156 16662
rect 8404 16590 8432 17002
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8024 16108 8076 16114
rect 8024 16050 8076 16056
rect 7262 15804 7558 15824
rect 7318 15802 7342 15804
rect 7398 15802 7422 15804
rect 7478 15802 7502 15804
rect 7340 15750 7342 15802
rect 7404 15750 7416 15802
rect 7478 15750 7480 15802
rect 7318 15748 7342 15750
rect 7398 15748 7422 15750
rect 7478 15748 7502 15750
rect 7262 15728 7558 15748
rect 8404 15638 8432 16526
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8404 15162 8432 15574
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 8680 15026 8708 15370
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4109 14172 4405 14192
rect 4165 14170 4189 14172
rect 4245 14170 4269 14172
rect 4325 14170 4349 14172
rect 4187 14118 4189 14170
rect 4251 14118 4263 14170
rect 4325 14118 4327 14170
rect 4165 14116 4189 14118
rect 4245 14116 4269 14118
rect 4325 14116 4349 14118
rect 4109 14096 4405 14116
rect 4540 13938 4568 14350
rect 4816 14074 4844 14554
rect 5644 14482 5672 14758
rect 7262 14716 7558 14736
rect 7318 14714 7342 14716
rect 7398 14714 7422 14716
rect 7478 14714 7502 14716
rect 7340 14662 7342 14714
rect 7404 14662 7416 14714
rect 7478 14662 7480 14714
rect 7318 14660 7342 14662
rect 7398 14660 7422 14662
rect 7478 14660 7502 14662
rect 7262 14640 7558 14660
rect 7944 14618 7972 14826
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8680 14482 8708 14962
rect 8956 14822 8984 18090
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17134 9168 17478
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9784 16726 9812 18022
rect 10244 17338 10272 20590
rect 10598 20583 10654 20590
rect 11886 20583 11942 21063
rect 12440 20596 12492 20602
rect 10415 18524 10711 18544
rect 10471 18522 10495 18524
rect 10551 18522 10575 18524
rect 10631 18522 10655 18524
rect 10493 18470 10495 18522
rect 10557 18470 10569 18522
rect 10631 18470 10633 18522
rect 10471 18468 10495 18470
rect 10551 18468 10575 18470
rect 10631 18468 10655 18470
rect 10415 18448 10711 18468
rect 11900 17746 11928 20583
rect 13174 20596 13230 21063
rect 14462 20618 14518 21063
rect 13174 20583 13176 20596
rect 12440 20538 12492 20544
rect 13228 20583 13230 20596
rect 14200 20590 14518 20618
rect 13176 20538 13228 20544
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10336 17202 10364 17478
rect 10415 17436 10711 17456
rect 10471 17434 10495 17436
rect 10551 17434 10575 17436
rect 10631 17434 10655 17436
rect 10493 17382 10495 17434
rect 10557 17382 10569 17434
rect 10631 17382 10633 17434
rect 10471 17380 10495 17382
rect 10551 17380 10575 17382
rect 10631 17380 10655 17382
rect 10415 17360 10711 17380
rect 11900 17338 11928 17682
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10612 16726 10640 17138
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9864 16720 9916 16726
rect 9864 16662 9916 16668
rect 10600 16720 10652 16726
rect 10600 16662 10652 16668
rect 9784 16250 9812 16662
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9876 16114 9904 16662
rect 10415 16348 10711 16368
rect 10471 16346 10495 16348
rect 10551 16346 10575 16348
rect 10631 16346 10655 16348
rect 10493 16294 10495 16346
rect 10557 16294 10569 16346
rect 10631 16294 10633 16346
rect 10471 16292 10495 16294
rect 10551 16292 10575 16294
rect 10631 16292 10655 16294
rect 10415 16272 10711 16292
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9876 15706 9904 16050
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9968 15502 9996 16050
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 10415 15260 10711 15280
rect 10471 15258 10495 15260
rect 10551 15258 10575 15260
rect 10631 15258 10655 15260
rect 10493 15206 10495 15258
rect 10557 15206 10569 15258
rect 10631 15206 10633 15258
rect 10471 15204 10495 15206
rect 10551 15204 10575 15206
rect 10631 15204 10655 15206
rect 10415 15184 10711 15204
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4540 13394 4568 13874
rect 4528 13388 4580 13394
rect 4528 13330 4580 13336
rect 4109 13084 4405 13104
rect 4165 13082 4189 13084
rect 4245 13082 4269 13084
rect 4325 13082 4349 13084
rect 4187 13030 4189 13082
rect 4251 13030 4263 13082
rect 4325 13030 4327 13082
rect 4165 13028 4189 13030
rect 4245 13028 4269 13030
rect 4325 13028 4349 13030
rect 4109 13008 4405 13028
rect 4540 12986 4568 13330
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4109 11996 4405 12016
rect 4165 11994 4189 11996
rect 4245 11994 4269 11996
rect 4325 11994 4349 11996
rect 4187 11942 4189 11994
rect 4251 11942 4263 11994
rect 4325 11942 4327 11994
rect 4165 11940 4189 11942
rect 4245 11940 4269 11942
rect 4325 11940 4349 11942
rect 4109 11920 4405 11940
rect 4618 11656 4674 11665
rect 4618 11591 4674 11600
rect 4632 11218 4660 11591
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4109 10908 4405 10928
rect 4165 10906 4189 10908
rect 4245 10906 4269 10908
rect 4325 10906 4349 10908
rect 4187 10854 4189 10906
rect 4251 10854 4263 10906
rect 4325 10854 4327 10906
rect 4165 10852 4189 10854
rect 4245 10852 4269 10854
rect 4325 10852 4349 10854
rect 4109 10832 4405 10852
rect 4632 10810 4660 11154
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4109 9820 4405 9840
rect 4165 9818 4189 9820
rect 4245 9818 4269 9820
rect 4325 9818 4349 9820
rect 4187 9766 4189 9818
rect 4251 9766 4263 9818
rect 4325 9766 4327 9818
rect 4165 9764 4189 9766
rect 4245 9764 4269 9766
rect 4325 9764 4349 9766
rect 4109 9744 4405 9764
rect 4109 8732 4405 8752
rect 4165 8730 4189 8732
rect 4245 8730 4269 8732
rect 4325 8730 4349 8732
rect 4187 8678 4189 8730
rect 4251 8678 4263 8730
rect 4325 8678 4327 8730
rect 4165 8676 4189 8678
rect 4245 8676 4269 8678
rect 4325 8676 4349 8678
rect 4109 8656 4405 8676
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4434 8120 4490 8129
rect 5000 8090 5028 8230
rect 4434 8055 4490 8064
rect 4988 8084 5040 8090
rect 4448 7954 4476 8055
rect 4988 8026 5040 8032
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4109 7644 4405 7664
rect 4165 7642 4189 7644
rect 4245 7642 4269 7644
rect 4325 7642 4349 7644
rect 4187 7590 4189 7642
rect 4251 7590 4263 7642
rect 4325 7590 4327 7642
rect 4165 7588 4189 7590
rect 4245 7588 4269 7590
rect 4325 7588 4349 7590
rect 4109 7568 4405 7588
rect 4448 7546 4476 7890
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4109 6556 4405 6576
rect 4165 6554 4189 6556
rect 4245 6554 4269 6556
rect 4325 6554 4349 6556
rect 4187 6502 4189 6554
rect 4251 6502 4263 6554
rect 4325 6502 4327 6554
rect 4165 6500 4189 6502
rect 4245 6500 4269 6502
rect 4325 6500 4349 6502
rect 4109 6480 4405 6500
rect 4109 5468 4405 5488
rect 4165 5466 4189 5468
rect 4245 5466 4269 5468
rect 4325 5466 4349 5468
rect 4187 5414 4189 5466
rect 4251 5414 4263 5466
rect 4325 5414 4327 5466
rect 4165 5412 4189 5414
rect 4245 5412 4269 5414
rect 4325 5412 4349 5414
rect 4109 5392 4405 5412
rect 4109 4380 4405 4400
rect 4165 4378 4189 4380
rect 4245 4378 4269 4380
rect 4325 4378 4349 4380
rect 4187 4326 4189 4378
rect 4251 4326 4263 4378
rect 4325 4326 4327 4378
rect 4165 4324 4189 4326
rect 4245 4324 4269 4326
rect 4325 4324 4349 4326
rect 4109 4304 4405 4324
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2650 3556 2790
rect 3804 2650 3832 3062
rect 3896 3058 3924 3470
rect 4109 3292 4405 3312
rect 4165 3290 4189 3292
rect 4245 3290 4269 3292
rect 4325 3290 4349 3292
rect 4187 3238 4189 3290
rect 4251 3238 4263 3290
rect 4325 3238 4327 3290
rect 4165 3236 4189 3238
rect 4245 3236 4269 3238
rect 4325 3236 4349 3238
rect 4109 3216 4405 3236
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4816 2990 4844 3470
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4816 2582 4844 2926
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4109 2204 4405 2224
rect 4165 2202 4189 2204
rect 4245 2202 4269 2204
rect 4325 2202 4349 2204
rect 4187 2150 4189 2202
rect 4251 2150 4263 2202
rect 4325 2150 4327 2202
rect 4165 2148 4189 2150
rect 4245 2148 4269 2150
rect 4325 2148 4349 2150
rect 4109 2128 4405 2148
rect 3422 82 3478 480
rect 3252 54 3478 82
rect 2686 31 2742 40
rect 3422 0 3478 54
rect 4434 82 4490 480
rect 4540 82 4568 2314
rect 4434 54 4568 82
rect 5092 82 5120 14214
rect 5644 14074 5672 14418
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9324 14074 9352 14214
rect 9692 14074 9720 14418
rect 10415 14172 10711 14192
rect 10471 14170 10495 14172
rect 10551 14170 10575 14172
rect 10631 14170 10655 14172
rect 10493 14118 10495 14170
rect 10557 14118 10569 14170
rect 10631 14118 10633 14170
rect 10471 14116 10495 14118
rect 10551 14116 10575 14118
rect 10631 14116 10655 14118
rect 10415 14096 10711 14116
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9324 13870 9352 14010
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 7262 13628 7558 13648
rect 7318 13626 7342 13628
rect 7398 13626 7422 13628
rect 7478 13626 7502 13628
rect 7340 13574 7342 13626
rect 7404 13574 7416 13626
rect 7478 13574 7480 13626
rect 7318 13572 7342 13574
rect 7398 13572 7422 13574
rect 7478 13572 7502 13574
rect 7262 13552 7558 13572
rect 7262 12540 7558 12560
rect 7318 12538 7342 12540
rect 7398 12538 7422 12540
rect 7478 12538 7502 12540
rect 7340 12486 7342 12538
rect 7404 12486 7416 12538
rect 7478 12486 7480 12538
rect 7318 12484 7342 12486
rect 7398 12484 7422 12486
rect 7478 12484 7502 12486
rect 7262 12464 7558 12484
rect 7262 11452 7558 11472
rect 7318 11450 7342 11452
rect 7398 11450 7422 11452
rect 7478 11450 7502 11452
rect 7340 11398 7342 11450
rect 7404 11398 7416 11450
rect 7478 11398 7480 11450
rect 7318 11396 7342 11398
rect 7398 11396 7422 11398
rect 7478 11396 7502 11398
rect 7262 11376 7558 11396
rect 7262 10364 7558 10384
rect 7318 10362 7342 10364
rect 7398 10362 7422 10364
rect 7478 10362 7502 10364
rect 7340 10310 7342 10362
rect 7404 10310 7416 10362
rect 7478 10310 7480 10362
rect 7318 10308 7342 10310
rect 7398 10308 7422 10310
rect 7478 10308 7502 10310
rect 7262 10288 7558 10308
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 9110 6408 9318
rect 7262 9276 7558 9296
rect 7318 9274 7342 9276
rect 7398 9274 7422 9276
rect 7478 9274 7502 9276
rect 7340 9222 7342 9274
rect 7404 9222 7416 9274
rect 7478 9222 7480 9274
rect 7318 9220 7342 9222
rect 7398 9220 7422 9222
rect 7478 9220 7502 9222
rect 7262 9200 7558 9220
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8498 5948 8910
rect 6380 8634 6408 9046
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5920 8022 5948 8434
rect 7262 8188 7558 8208
rect 7318 8186 7342 8188
rect 7398 8186 7422 8188
rect 7478 8186 7502 8188
rect 7340 8134 7342 8186
rect 7404 8134 7416 8186
rect 7478 8134 7480 8186
rect 7318 8132 7342 8134
rect 7398 8132 7422 8134
rect 7478 8132 7502 8134
rect 7262 8112 7558 8132
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6380 7546 6408 7958
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 6934 6868 7142
rect 7024 6934 7052 7822
rect 7262 7100 7558 7120
rect 7318 7098 7342 7100
rect 7398 7098 7422 7100
rect 7478 7098 7502 7100
rect 7340 7046 7342 7098
rect 7404 7046 7416 7098
rect 7478 7046 7480 7098
rect 7318 7044 7342 7046
rect 7398 7044 7422 7046
rect 7478 7044 7502 7046
rect 7262 7024 7558 7044
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6380 6458 6408 6870
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6458 7512 6598
rect 7852 6458 7880 6802
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7484 6254 7512 6394
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6288 3670 6316 3878
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6288 3194 6316 3606
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6932 3058 6960 3470
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2650 6960 2790
rect 7024 2650 7052 3878
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 6734 2000 6790 2009
rect 6734 1935 6790 1944
rect 5446 82 5502 480
rect 5092 54 5502 82
rect 4434 0 4490 54
rect 5446 0 5502 54
rect 6458 82 6514 480
rect 6748 82 6776 1935
rect 6458 54 6776 82
rect 7116 82 7144 6054
rect 7262 6012 7558 6032
rect 7318 6010 7342 6012
rect 7398 6010 7422 6012
rect 7478 6010 7502 6012
rect 7340 5958 7342 6010
rect 7404 5958 7416 6010
rect 7478 5958 7480 6010
rect 7318 5956 7342 5958
rect 7398 5956 7422 5958
rect 7478 5956 7502 5958
rect 7262 5936 7558 5956
rect 7262 4924 7558 4944
rect 7318 4922 7342 4924
rect 7398 4922 7422 4924
rect 7478 4922 7502 4924
rect 7340 4870 7342 4922
rect 7404 4870 7416 4922
rect 7478 4870 7480 4922
rect 7318 4868 7342 4870
rect 7398 4868 7422 4870
rect 7478 4868 7502 4870
rect 7262 4848 7558 4868
rect 7262 3836 7558 3856
rect 7318 3834 7342 3836
rect 7398 3834 7422 3836
rect 7478 3834 7502 3836
rect 7340 3782 7342 3834
rect 7404 3782 7416 3834
rect 7478 3782 7480 3834
rect 7318 3780 7342 3782
rect 7398 3780 7422 3782
rect 7478 3780 7502 3782
rect 7262 3760 7558 3780
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7760 2854 7788 3538
rect 8208 3392 8260 3398
rect 8208 3334 8260 3340
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7262 2748 7558 2768
rect 7318 2746 7342 2748
rect 7398 2746 7422 2748
rect 7478 2746 7502 2748
rect 7340 2694 7342 2746
rect 7404 2694 7416 2746
rect 7478 2694 7480 2746
rect 7318 2692 7342 2694
rect 7398 2692 7422 2694
rect 7478 2692 7502 2694
rect 7262 2672 7558 2692
rect 8036 2582 8064 2858
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7378 82 7434 480
rect 7116 54 7434 82
rect 8220 82 8248 3334
rect 8390 82 8446 480
rect 8220 54 8446 82
rect 9048 82 9076 13670
rect 10415 13084 10711 13104
rect 10471 13082 10495 13084
rect 10551 13082 10575 13084
rect 10631 13082 10655 13084
rect 10493 13030 10495 13082
rect 10557 13030 10569 13082
rect 10631 13030 10633 13082
rect 10471 13028 10495 13030
rect 10551 13028 10575 13030
rect 10631 13028 10655 13030
rect 10415 13008 10711 13028
rect 10415 11996 10711 12016
rect 10471 11994 10495 11996
rect 10551 11994 10575 11996
rect 10631 11994 10655 11996
rect 10493 11942 10495 11994
rect 10557 11942 10569 11994
rect 10631 11942 10633 11994
rect 10471 11940 10495 11942
rect 10551 11940 10575 11942
rect 10631 11940 10655 11942
rect 10415 11920 10711 11940
rect 10415 10908 10711 10928
rect 10471 10906 10495 10908
rect 10551 10906 10575 10908
rect 10631 10906 10655 10908
rect 10493 10854 10495 10906
rect 10557 10854 10569 10906
rect 10631 10854 10633 10906
rect 10471 10852 10495 10854
rect 10551 10852 10575 10854
rect 10631 10852 10655 10854
rect 10415 10832 10711 10852
rect 10415 9820 10711 9840
rect 10471 9818 10495 9820
rect 10551 9818 10575 9820
rect 10631 9818 10655 9820
rect 10493 9766 10495 9818
rect 10557 9766 10569 9818
rect 10631 9766 10633 9818
rect 10471 9764 10495 9766
rect 10551 9764 10575 9766
rect 10631 9764 10655 9766
rect 10415 9744 10711 9764
rect 12452 9722 12480 20538
rect 13188 20507 13216 20538
rect 14200 18426 14228 20590
rect 14462 20583 14518 20590
rect 15212 20590 15608 20618
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14200 18222 14228 18362
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13912 18080 13964 18086
rect 13912 18022 13964 18028
rect 13569 17980 13865 18000
rect 13625 17978 13649 17980
rect 13705 17978 13729 17980
rect 13785 17978 13809 17980
rect 13647 17926 13649 17978
rect 13711 17926 13723 17978
rect 13785 17926 13787 17978
rect 13625 17924 13649 17926
rect 13705 17924 13729 17926
rect 13785 17924 13809 17926
rect 13569 17904 13865 17924
rect 12622 17776 12678 17785
rect 12622 17711 12624 17720
rect 12676 17711 12678 17720
rect 12624 17682 12676 17688
rect 12636 17338 12664 17682
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17338 13032 17478
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13569 16892 13865 16912
rect 13625 16890 13649 16892
rect 13705 16890 13729 16892
rect 13785 16890 13809 16892
rect 13647 16838 13649 16890
rect 13711 16838 13723 16890
rect 13785 16838 13787 16890
rect 13625 16836 13649 16838
rect 13705 16836 13729 16838
rect 13785 16836 13809 16838
rect 13569 16816 13865 16836
rect 13924 16726 13952 18022
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14200 17338 14228 17682
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13924 16250 13952 16662
rect 14016 16590 14044 17002
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 14016 16250 14044 16526
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 13569 15804 13865 15824
rect 13625 15802 13649 15804
rect 13705 15802 13729 15804
rect 13785 15802 13809 15804
rect 13647 15750 13649 15802
rect 13711 15750 13723 15802
rect 13785 15750 13787 15802
rect 13625 15748 13649 15750
rect 13705 15748 13729 15750
rect 13785 15748 13809 15750
rect 13569 15728 13865 15748
rect 13569 14716 13865 14736
rect 13625 14714 13649 14716
rect 13705 14714 13729 14716
rect 13785 14714 13809 14716
rect 13647 14662 13649 14714
rect 13711 14662 13723 14714
rect 13785 14662 13787 14714
rect 13625 14660 13649 14662
rect 13705 14660 13729 14662
rect 13785 14660 13809 14662
rect 13569 14640 13865 14660
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 13569 13628 13865 13648
rect 13625 13626 13649 13628
rect 13705 13626 13729 13628
rect 13785 13626 13809 13628
rect 13647 13574 13649 13626
rect 13711 13574 13723 13626
rect 13785 13574 13787 13626
rect 13625 13572 13649 13574
rect 13705 13572 13729 13574
rect 13785 13572 13809 13574
rect 13569 13552 13865 13572
rect 14660 13462 14688 13670
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 13569 12540 13865 12560
rect 13625 12538 13649 12540
rect 13705 12538 13729 12540
rect 13785 12538 13809 12540
rect 13647 12486 13649 12538
rect 13711 12486 13723 12538
rect 13785 12486 13787 12538
rect 13625 12484 13649 12486
rect 13705 12484 13729 12486
rect 13785 12484 13809 12486
rect 13569 12464 13865 12484
rect 15212 11665 15240 20590
rect 15580 20584 15608 20590
rect 15658 20584 15714 21063
rect 15580 20583 15714 20584
rect 16946 20618 17002 21063
rect 16946 20590 17080 20618
rect 16946 20583 17002 20590
rect 15580 20556 15700 20583
rect 16722 18524 17018 18544
rect 16778 18522 16802 18524
rect 16858 18522 16882 18524
rect 16938 18522 16962 18524
rect 16800 18470 16802 18522
rect 16864 18470 16876 18522
rect 16938 18470 16940 18522
rect 16778 18468 16802 18470
rect 16858 18468 16882 18470
rect 16938 18468 16962 18470
rect 16722 18448 17018 18468
rect 17052 18290 17080 20590
rect 18234 20583 18290 21063
rect 18248 18426 18276 20583
rect 18510 20360 18566 20369
rect 18510 20295 18566 20304
rect 18418 19136 18474 19145
rect 18418 19071 18474 19080
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18432 18358 18460 19071
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 18524 18154 18552 20295
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15476 17060 15528 17066
rect 15476 17002 15528 17008
rect 15292 16992 15344 16998
rect 15488 16969 15516 17002
rect 15292 16934 15344 16940
rect 15474 16960 15530 16969
rect 15304 15638 15332 16934
rect 15474 16895 15530 16904
rect 15672 16114 15700 17546
rect 15764 17338 15792 17614
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 16040 17202 16068 18022
rect 16722 17436 17018 17456
rect 16778 17434 16802 17436
rect 16858 17434 16882 17436
rect 16938 17434 16962 17436
rect 16800 17382 16802 17434
rect 16864 17382 16876 17434
rect 16938 17382 16940 17434
rect 16778 17380 16802 17382
rect 16858 17380 16882 17382
rect 16938 17380 16962 17382
rect 16722 17360 17018 17380
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 16040 16794 16068 17138
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15292 15632 15344 15638
rect 15292 15574 15344 15580
rect 15304 15162 15332 15574
rect 15672 15502 15700 16050
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15764 12986 15792 13398
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15198 11656 15254 11665
rect 15198 11591 15254 11600
rect 13569 11452 13865 11472
rect 13625 11450 13649 11452
rect 13705 11450 13729 11452
rect 13785 11450 13809 11452
rect 13647 11398 13649 11450
rect 13711 11398 13723 11450
rect 13785 11398 13787 11450
rect 13625 11396 13649 11398
rect 13705 11396 13729 11398
rect 13785 11396 13809 11398
rect 13569 11376 13865 11396
rect 14830 11248 14886 11257
rect 14830 11183 14886 11192
rect 13569 10364 13865 10384
rect 13625 10362 13649 10364
rect 13705 10362 13729 10364
rect 13785 10362 13809 10364
rect 13647 10310 13649 10362
rect 13711 10310 13723 10362
rect 13785 10310 13787 10362
rect 13625 10308 13649 10310
rect 13705 10308 13729 10310
rect 13785 10308 13809 10310
rect 13569 10288 13865 10308
rect 14462 10024 14518 10033
rect 14462 9959 14518 9968
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 13569 9276 13865 9296
rect 13625 9274 13649 9276
rect 13705 9274 13729 9276
rect 13785 9274 13809 9276
rect 13647 9222 13649 9274
rect 13711 9222 13723 9274
rect 13785 9222 13787 9274
rect 13625 9220 13649 9222
rect 13705 9220 13729 9222
rect 13785 9220 13809 9222
rect 13569 9200 13865 9220
rect 10415 8732 10711 8752
rect 10471 8730 10495 8732
rect 10551 8730 10575 8732
rect 10631 8730 10655 8732
rect 10493 8678 10495 8730
rect 10557 8678 10569 8730
rect 10631 8678 10633 8730
rect 10471 8676 10495 8678
rect 10551 8676 10575 8678
rect 10631 8676 10655 8678
rect 10415 8656 10711 8676
rect 13569 8188 13865 8208
rect 13625 8186 13649 8188
rect 13705 8186 13729 8188
rect 13785 8186 13809 8188
rect 13647 8134 13649 8186
rect 13711 8134 13723 8186
rect 13785 8134 13787 8186
rect 13625 8132 13649 8134
rect 13705 8132 13729 8134
rect 13785 8132 13809 8134
rect 13569 8112 13865 8132
rect 10415 7644 10711 7664
rect 10471 7642 10495 7644
rect 10551 7642 10575 7644
rect 10631 7642 10655 7644
rect 10493 7590 10495 7642
rect 10557 7590 10569 7642
rect 10631 7590 10633 7642
rect 10471 7588 10495 7590
rect 10551 7588 10575 7590
rect 10631 7588 10655 7590
rect 10415 7568 10711 7588
rect 14476 7546 14504 9959
rect 14844 7954 14872 11183
rect 15948 10674 15976 16050
rect 16040 13462 16068 16526
rect 16132 14550 16160 17138
rect 16722 16348 17018 16368
rect 16778 16346 16802 16348
rect 16858 16346 16882 16348
rect 16938 16346 16962 16348
rect 16800 16294 16802 16346
rect 16864 16294 16876 16346
rect 16938 16294 16940 16346
rect 16778 16292 16802 16294
rect 16858 16292 16882 16294
rect 16938 16292 16962 16294
rect 16722 16272 17018 16292
rect 16722 15260 17018 15280
rect 16778 15258 16802 15260
rect 16858 15258 16882 15260
rect 16938 15258 16962 15260
rect 16800 15206 16802 15258
rect 16864 15206 16876 15258
rect 16938 15206 16940 15258
rect 16778 15204 16802 15206
rect 16858 15204 16882 15206
rect 16938 15204 16962 15206
rect 16722 15184 17018 15204
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 16132 14074 16160 14486
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16040 12986 16068 13398
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16132 11150 16160 14010
rect 16224 13870 16252 14758
rect 16316 14414 16344 14962
rect 16486 14920 16542 14929
rect 16486 14855 16542 14864
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16500 14074 16528 14855
rect 16722 14172 17018 14192
rect 16778 14170 16802 14172
rect 16858 14170 16882 14172
rect 16938 14170 16962 14172
rect 16800 14118 16802 14170
rect 16864 14118 16876 14170
rect 16938 14118 16940 14170
rect 16778 14116 16802 14118
rect 16858 14116 16882 14118
rect 16938 14116 16962 14118
rect 16722 14096 17018 14116
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16040 10810 16068 11086
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10130 15976 10610
rect 16040 10266 16068 10746
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15396 9722 15424 10066
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9722 16160 9862
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16132 9518 16160 9658
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16500 9178 16528 13631
rect 16722 13084 17018 13104
rect 16778 13082 16802 13084
rect 16858 13082 16882 13084
rect 16938 13082 16962 13084
rect 16800 13030 16802 13082
rect 16864 13030 16876 13082
rect 16938 13030 16940 13082
rect 16778 13028 16802 13030
rect 16858 13028 16882 13030
rect 16938 13028 16962 13030
rect 16722 13008 17018 13028
rect 17130 13016 17186 13025
rect 17130 12951 17186 12960
rect 17144 12918 17172 12951
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 16722 11996 17018 12016
rect 16778 11994 16802 11996
rect 16858 11994 16882 11996
rect 16938 11994 16962 11996
rect 16800 11942 16802 11994
rect 16864 11942 16876 11994
rect 16938 11942 16940 11994
rect 16778 11940 16802 11942
rect 16858 11940 16882 11942
rect 16938 11940 16962 11942
rect 16722 11920 17018 11940
rect 16722 10908 17018 10928
rect 16778 10906 16802 10908
rect 16858 10906 16882 10908
rect 16938 10906 16962 10908
rect 16800 10854 16802 10906
rect 16864 10854 16876 10906
rect 16938 10854 16940 10906
rect 16778 10852 16802 10854
rect 16858 10852 16882 10854
rect 16938 10852 16962 10854
rect 16722 10832 17018 10852
rect 17040 10124 17092 10130
rect 17040 10066 17092 10072
rect 16722 9820 17018 9840
rect 16778 9818 16802 9820
rect 16858 9818 16882 9820
rect 16938 9818 16962 9820
rect 16800 9766 16802 9818
rect 16864 9766 16876 9818
rect 16938 9766 16940 9818
rect 16778 9764 16802 9766
rect 16858 9764 16882 9766
rect 16938 9764 16962 9766
rect 16722 9744 17018 9764
rect 17052 9382 17080 10066
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 15212 8634 15240 8978
rect 16316 8634 16344 8978
rect 16722 8732 17018 8752
rect 16778 8730 16802 8732
rect 16858 8730 16882 8732
rect 16938 8730 16962 8732
rect 16800 8678 16802 8730
rect 16864 8678 16876 8730
rect 16938 8678 16940 8730
rect 16778 8676 16802 8678
rect 16858 8676 16882 8678
rect 16938 8676 16962 8678
rect 16722 8656 17018 8676
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 15474 7984 15530 7993
rect 14832 7948 14884 7954
rect 15474 7919 15530 7928
rect 14832 7890 14884 7896
rect 14844 7546 14872 7890
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14476 7342 14504 7482
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 13569 7100 13865 7120
rect 13625 7098 13649 7100
rect 13705 7098 13729 7100
rect 13785 7098 13809 7100
rect 13647 7046 13649 7098
rect 13711 7046 13723 7098
rect 13785 7046 13787 7098
rect 13625 7044 13649 7046
rect 13705 7044 13729 7046
rect 13785 7044 13809 7046
rect 13569 7024 13865 7044
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10415 6556 10711 6576
rect 10471 6554 10495 6556
rect 10551 6554 10575 6556
rect 10631 6554 10655 6556
rect 10493 6502 10495 6554
rect 10557 6502 10569 6554
rect 10631 6502 10633 6554
rect 10471 6500 10495 6502
rect 10551 6500 10575 6502
rect 10631 6500 10655 6502
rect 10415 6480 10711 6500
rect 10415 5468 10711 5488
rect 10471 5466 10495 5468
rect 10551 5466 10575 5468
rect 10631 5466 10655 5468
rect 10493 5414 10495 5466
rect 10557 5414 10569 5466
rect 10631 5414 10633 5466
rect 10471 5412 10495 5414
rect 10551 5412 10575 5414
rect 10631 5412 10655 5414
rect 10415 5392 10711 5412
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 3058 9352 4966
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 4146 10272 4626
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10415 4380 10711 4400
rect 10471 4378 10495 4380
rect 10551 4378 10575 4380
rect 10631 4378 10655 4380
rect 10493 4326 10495 4378
rect 10557 4326 10569 4378
rect 10631 4326 10633 4378
rect 10471 4324 10495 4326
rect 10551 4324 10575 4326
rect 10631 4324 10655 4326
rect 10415 4304 10711 4324
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 9600 3670 9628 3878
rect 9588 3664 9640 3670
rect 9588 3606 9640 3612
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10244 3194 10272 3606
rect 10336 3194 10364 3878
rect 10415 3292 10711 3312
rect 10471 3290 10495 3292
rect 10551 3290 10575 3292
rect 10631 3290 10655 3292
rect 10493 3238 10495 3290
rect 10557 3238 10569 3290
rect 10631 3238 10633 3290
rect 10471 3236 10495 3238
rect 10551 3236 10575 3238
rect 10631 3236 10655 3238
rect 10415 3216 10711 3236
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10888 3058 10916 4422
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2582 11008 6598
rect 13464 6118 13492 6802
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14476 6186 14504 6666
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12346 5128 12402 5137
rect 12346 5063 12402 5072
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4684 11204 4690
rect 11072 4644 11152 4672
rect 11072 3942 11100 4644
rect 11152 4626 11204 4632
rect 11256 4154 11284 4966
rect 12360 4826 12388 5063
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 12176 4282 12204 4626
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 11164 4126 11284 4154
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 2854 11100 3878
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10415 2204 10711 2224
rect 10471 2202 10495 2204
rect 10551 2202 10575 2204
rect 10631 2202 10655 2204
rect 10493 2150 10495 2202
rect 10557 2150 10569 2202
rect 10631 2150 10633 2202
rect 10471 2148 10495 2150
rect 10551 2148 10575 2150
rect 10631 2148 10655 2150
rect 10415 2128 10711 2148
rect 9402 82 9458 480
rect 9048 54 9458 82
rect 6458 0 6514 54
rect 7378 0 7434 54
rect 8390 0 8446 54
rect 9402 0 9458 54
rect 10414 96 10470 480
rect 11164 82 11192 4126
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 11348 2514 11376 3878
rect 12360 3534 12388 3878
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 11440 3126 11468 3470
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 12360 3058 12388 3470
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12452 2650 12480 4966
rect 12544 4282 12572 5646
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12728 4214 12756 5034
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 13004 3602 13032 6054
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 13464 2922 13492 6054
rect 13569 6012 13865 6032
rect 13625 6010 13649 6012
rect 13705 6010 13729 6012
rect 13785 6010 13809 6012
rect 13647 5958 13649 6010
rect 13711 5958 13723 6010
rect 13785 5958 13787 6010
rect 13625 5956 13649 5958
rect 13705 5956 13729 5958
rect 13785 5956 13809 5958
rect 13569 5936 13865 5956
rect 13569 4924 13865 4944
rect 13625 4922 13649 4924
rect 13705 4922 13729 4924
rect 13785 4922 13809 4924
rect 13647 4870 13649 4922
rect 13711 4870 13723 4922
rect 13785 4870 13787 4922
rect 13625 4868 13649 4870
rect 13705 4868 13729 4870
rect 13785 4868 13809 4870
rect 13569 4848 13865 4868
rect 13924 4758 13952 6054
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14004 5092 14056 5098
rect 14004 5034 14056 5040
rect 14016 4758 14044 5034
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 14004 4752 14056 4758
rect 14004 4694 14056 4700
rect 13924 4282 13952 4694
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 13569 3836 13865 3856
rect 13625 3834 13649 3836
rect 13705 3834 13729 3836
rect 13785 3834 13809 3836
rect 13647 3782 13649 3834
rect 13711 3782 13723 3834
rect 13785 3782 13787 3834
rect 13625 3780 13649 3782
rect 13705 3780 13729 3782
rect 13785 3780 13809 3782
rect 13569 3760 13865 3780
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13832 3194 13860 3538
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13569 2748 13865 2768
rect 13625 2746 13649 2748
rect 13705 2746 13729 2748
rect 13785 2746 13809 2748
rect 13647 2694 13649 2746
rect 13711 2694 13723 2746
rect 13785 2694 13787 2746
rect 13625 2692 13649 2694
rect 13705 2692 13729 2694
rect 13785 2692 13809 2694
rect 13569 2672 13865 2692
rect 12164 2644 12216 2650
rect 12164 2586 12216 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 11426 82 11482 480
rect 11164 54 11482 82
rect 12176 82 12204 2586
rect 13924 2582 13952 2858
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 12438 82 12494 480
rect 12176 54 12494 82
rect 13096 82 13124 2314
rect 14016 2009 14044 3334
rect 14108 3194 14136 5646
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14002 2000 14058 2009
rect 14002 1935 14058 1944
rect 13358 82 13414 480
rect 13096 54 13414 82
rect 14200 82 14228 6054
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 14292 4010 14320 5034
rect 14280 4004 14332 4010
rect 14280 3946 14332 3952
rect 14568 3534 14596 6258
rect 14844 4622 14872 7210
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 15028 5370 15056 6054
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 3058 14596 3470
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 15304 2650 15332 6598
rect 15396 5846 15424 7686
rect 15488 7546 15516 7919
rect 16408 7886 16436 8434
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15488 7342 15516 7482
rect 16316 7410 16344 7822
rect 16722 7644 17018 7664
rect 16778 7642 16802 7644
rect 16858 7642 16882 7644
rect 16938 7642 16962 7644
rect 16800 7590 16802 7642
rect 16864 7590 16876 7642
rect 16938 7590 16940 7642
rect 16778 7588 16802 7590
rect 16858 7588 16882 7590
rect 16938 7588 16962 7590
rect 16722 7568 17018 7588
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 16316 6798 16344 7346
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15948 6458 15976 6734
rect 16722 6556 17018 6576
rect 16778 6554 16802 6556
rect 16858 6554 16882 6556
rect 16938 6554 16962 6556
rect 16800 6502 16802 6554
rect 16864 6502 16876 6554
rect 16938 6502 16940 6554
rect 16778 6500 16802 6502
rect 16858 6500 16882 6502
rect 16938 6500 16962 6502
rect 16722 6480 17018 6500
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16212 6112 16264 6118
rect 17052 6089 17080 9318
rect 18432 9217 18460 9590
rect 18418 9208 18474 9217
rect 18418 9143 18474 9152
rect 17130 6488 17186 6497
rect 17130 6423 17186 6432
rect 17144 6390 17172 6423
rect 17132 6384 17184 6390
rect 17132 6326 17184 6332
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 16212 6054 16264 6060
rect 17038 6080 17094 6089
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15396 5302 15424 5782
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15292 2644 15344 2650
rect 15292 2586 15344 2592
rect 14370 82 14426 480
rect 14200 54 14426 82
rect 10414 0 10470 40
rect 11426 0 11482 54
rect 12438 0 12494 54
rect 13358 0 13414 54
rect 14370 0 14426 54
rect 15382 82 15438 480
rect 15488 82 15516 5170
rect 15672 4758 15700 5646
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15752 4616 15804 4622
rect 15752 4558 15804 4564
rect 15580 4282 15608 4558
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15764 4146 15792 4558
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15764 3670 15792 4082
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15764 3194 15792 3606
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15382 54 15516 82
rect 16224 82 16252 6054
rect 17038 6015 17094 6024
rect 16722 5468 17018 5488
rect 16778 5466 16802 5468
rect 16858 5466 16882 5468
rect 16938 5466 16962 5468
rect 16800 5414 16802 5466
rect 16864 5414 16876 5466
rect 16938 5414 16940 5466
rect 16778 5412 16802 5414
rect 16858 5412 16882 5414
rect 16938 5412 16962 5414
rect 16722 5392 17018 5412
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16316 3058 16344 5170
rect 16722 4380 17018 4400
rect 16778 4378 16802 4380
rect 16858 4378 16882 4380
rect 16938 4378 16962 4380
rect 16800 4326 16802 4378
rect 16864 4326 16876 4378
rect 16938 4326 16940 4378
rect 16778 4324 16802 4326
rect 16858 4324 16882 4326
rect 16938 4324 16962 4326
rect 16722 4304 17018 4324
rect 16722 3292 17018 3312
rect 16778 3290 16802 3292
rect 16858 3290 16882 3292
rect 16938 3290 16962 3292
rect 16800 3238 16802 3290
rect 16864 3238 16876 3290
rect 16938 3238 16940 3290
rect 16778 3236 16802 3238
rect 16858 3236 16882 3238
rect 16938 3236 16962 3238
rect 16722 3216 17018 3236
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16316 2446 16344 2994
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 16722 2204 17018 2224
rect 16778 2202 16802 2204
rect 16858 2202 16882 2204
rect 16938 2202 16962 2204
rect 16800 2150 16802 2202
rect 16864 2150 16876 2202
rect 16938 2150 16940 2202
rect 16778 2148 16802 2150
rect 16858 2148 16882 2150
rect 16938 2148 16962 2150
rect 16722 2128 17018 2148
rect 16394 82 16450 480
rect 16224 54 16450 82
rect 17236 82 17264 6258
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 17406 82 17462 480
rect 17236 54 17462 82
rect 15382 0 15438 54
rect 16394 0 16450 54
rect 17406 0 17462 54
rect 18418 82 18474 480
rect 18524 82 18552 2790
rect 18418 54 18552 82
rect 18418 0 18474 54
<< via2 >>
rect 1214 19488 1270 19544
rect 1766 17720 1822 17776
rect 1766 17584 1822 17640
rect 110 14320 166 14376
rect 110 12416 166 12472
rect 1306 9968 1362 10024
rect 110 6704 166 6760
rect 4109 18522 4165 18524
rect 4189 18522 4245 18524
rect 4269 18522 4325 18524
rect 4349 18522 4405 18524
rect 4109 18470 4135 18522
rect 4135 18470 4165 18522
rect 4189 18470 4199 18522
rect 4199 18470 4245 18522
rect 4269 18470 4315 18522
rect 4315 18470 4325 18522
rect 4349 18470 4379 18522
rect 4379 18470 4405 18522
rect 4109 18468 4165 18470
rect 4189 18468 4245 18470
rect 4269 18468 4325 18470
rect 4349 18468 4405 18470
rect 4109 17434 4165 17436
rect 4189 17434 4245 17436
rect 4269 17434 4325 17436
rect 4349 17434 4405 17436
rect 4109 17382 4135 17434
rect 4135 17382 4165 17434
rect 4189 17382 4199 17434
rect 4199 17382 4245 17434
rect 4269 17382 4315 17434
rect 4315 17382 4325 17434
rect 4349 17382 4379 17434
rect 4379 17382 4405 17434
rect 4109 17380 4165 17382
rect 4189 17380 4245 17382
rect 4269 17380 4325 17382
rect 4349 17380 4405 17382
rect 4109 16346 4165 16348
rect 4189 16346 4245 16348
rect 4269 16346 4325 16348
rect 4349 16346 4405 16348
rect 4109 16294 4135 16346
rect 4135 16294 4165 16346
rect 4189 16294 4199 16346
rect 4199 16294 4245 16346
rect 4269 16294 4315 16346
rect 4315 16294 4325 16346
rect 4349 16294 4379 16346
rect 4379 16294 4405 16346
rect 4109 16292 4165 16294
rect 4189 16292 4245 16294
rect 4269 16292 4325 16294
rect 4349 16292 4405 16294
rect 3974 15680 4030 15736
rect 1674 3984 1730 4040
rect 2686 40 2742 96
rect 4109 15258 4165 15260
rect 4189 15258 4245 15260
rect 4269 15258 4325 15260
rect 4349 15258 4405 15260
rect 4109 15206 4135 15258
rect 4135 15206 4165 15258
rect 4189 15206 4199 15258
rect 4199 15206 4245 15258
rect 4269 15206 4315 15258
rect 4315 15206 4325 15258
rect 4349 15206 4379 15258
rect 4379 15206 4405 15258
rect 4109 15204 4165 15206
rect 4189 15204 4245 15206
rect 4269 15204 4325 15206
rect 4349 15204 4405 15206
rect 7470 18128 7526 18184
rect 7262 17978 7318 17980
rect 7342 17978 7398 17980
rect 7422 17978 7478 17980
rect 7502 17978 7558 17980
rect 7262 17926 7288 17978
rect 7288 17926 7318 17978
rect 7342 17926 7352 17978
rect 7352 17926 7398 17978
rect 7422 17926 7468 17978
rect 7468 17926 7478 17978
rect 7502 17926 7532 17978
rect 7532 17926 7558 17978
rect 7262 17924 7318 17926
rect 7342 17924 7398 17926
rect 7422 17924 7478 17926
rect 7502 17924 7558 17926
rect 7262 16890 7318 16892
rect 7342 16890 7398 16892
rect 7422 16890 7478 16892
rect 7502 16890 7558 16892
rect 7262 16838 7288 16890
rect 7288 16838 7318 16890
rect 7342 16838 7352 16890
rect 7352 16838 7398 16890
rect 7422 16838 7468 16890
rect 7468 16838 7478 16890
rect 7502 16838 7532 16890
rect 7532 16838 7558 16890
rect 7262 16836 7318 16838
rect 7342 16836 7398 16838
rect 7422 16836 7478 16838
rect 7502 16836 7558 16838
rect 7262 15802 7318 15804
rect 7342 15802 7398 15804
rect 7422 15802 7478 15804
rect 7502 15802 7558 15804
rect 7262 15750 7288 15802
rect 7288 15750 7318 15802
rect 7342 15750 7352 15802
rect 7352 15750 7398 15802
rect 7422 15750 7468 15802
rect 7468 15750 7478 15802
rect 7502 15750 7532 15802
rect 7532 15750 7558 15802
rect 7262 15748 7318 15750
rect 7342 15748 7398 15750
rect 7422 15748 7478 15750
rect 7502 15748 7558 15750
rect 4109 14170 4165 14172
rect 4189 14170 4245 14172
rect 4269 14170 4325 14172
rect 4349 14170 4405 14172
rect 4109 14118 4135 14170
rect 4135 14118 4165 14170
rect 4189 14118 4199 14170
rect 4199 14118 4245 14170
rect 4269 14118 4315 14170
rect 4315 14118 4325 14170
rect 4349 14118 4379 14170
rect 4379 14118 4405 14170
rect 4109 14116 4165 14118
rect 4189 14116 4245 14118
rect 4269 14116 4325 14118
rect 4349 14116 4405 14118
rect 7262 14714 7318 14716
rect 7342 14714 7398 14716
rect 7422 14714 7478 14716
rect 7502 14714 7558 14716
rect 7262 14662 7288 14714
rect 7288 14662 7318 14714
rect 7342 14662 7352 14714
rect 7352 14662 7398 14714
rect 7422 14662 7468 14714
rect 7468 14662 7478 14714
rect 7502 14662 7532 14714
rect 7532 14662 7558 14714
rect 7262 14660 7318 14662
rect 7342 14660 7398 14662
rect 7422 14660 7478 14662
rect 7502 14660 7558 14662
rect 10415 18522 10471 18524
rect 10495 18522 10551 18524
rect 10575 18522 10631 18524
rect 10655 18522 10711 18524
rect 10415 18470 10441 18522
rect 10441 18470 10471 18522
rect 10495 18470 10505 18522
rect 10505 18470 10551 18522
rect 10575 18470 10621 18522
rect 10621 18470 10631 18522
rect 10655 18470 10685 18522
rect 10685 18470 10711 18522
rect 10415 18468 10471 18470
rect 10495 18468 10551 18470
rect 10575 18468 10631 18470
rect 10655 18468 10711 18470
rect 10415 17434 10471 17436
rect 10495 17434 10551 17436
rect 10575 17434 10631 17436
rect 10655 17434 10711 17436
rect 10415 17382 10441 17434
rect 10441 17382 10471 17434
rect 10495 17382 10505 17434
rect 10505 17382 10551 17434
rect 10575 17382 10621 17434
rect 10621 17382 10631 17434
rect 10655 17382 10685 17434
rect 10685 17382 10711 17434
rect 10415 17380 10471 17382
rect 10495 17380 10551 17382
rect 10575 17380 10631 17382
rect 10655 17380 10711 17382
rect 10415 16346 10471 16348
rect 10495 16346 10551 16348
rect 10575 16346 10631 16348
rect 10655 16346 10711 16348
rect 10415 16294 10441 16346
rect 10441 16294 10471 16346
rect 10495 16294 10505 16346
rect 10505 16294 10551 16346
rect 10575 16294 10621 16346
rect 10621 16294 10631 16346
rect 10655 16294 10685 16346
rect 10685 16294 10711 16346
rect 10415 16292 10471 16294
rect 10495 16292 10551 16294
rect 10575 16292 10631 16294
rect 10655 16292 10711 16294
rect 10415 15258 10471 15260
rect 10495 15258 10551 15260
rect 10575 15258 10631 15260
rect 10655 15258 10711 15260
rect 10415 15206 10441 15258
rect 10441 15206 10471 15258
rect 10495 15206 10505 15258
rect 10505 15206 10551 15258
rect 10575 15206 10621 15258
rect 10621 15206 10631 15258
rect 10655 15206 10685 15258
rect 10685 15206 10711 15258
rect 10415 15204 10471 15206
rect 10495 15204 10551 15206
rect 10575 15204 10631 15206
rect 10655 15204 10711 15206
rect 4109 13082 4165 13084
rect 4189 13082 4245 13084
rect 4269 13082 4325 13084
rect 4349 13082 4405 13084
rect 4109 13030 4135 13082
rect 4135 13030 4165 13082
rect 4189 13030 4199 13082
rect 4199 13030 4245 13082
rect 4269 13030 4315 13082
rect 4315 13030 4325 13082
rect 4349 13030 4379 13082
rect 4379 13030 4405 13082
rect 4109 13028 4165 13030
rect 4189 13028 4245 13030
rect 4269 13028 4325 13030
rect 4349 13028 4405 13030
rect 4109 11994 4165 11996
rect 4189 11994 4245 11996
rect 4269 11994 4325 11996
rect 4349 11994 4405 11996
rect 4109 11942 4135 11994
rect 4135 11942 4165 11994
rect 4189 11942 4199 11994
rect 4199 11942 4245 11994
rect 4269 11942 4315 11994
rect 4315 11942 4325 11994
rect 4349 11942 4379 11994
rect 4379 11942 4405 11994
rect 4109 11940 4165 11942
rect 4189 11940 4245 11942
rect 4269 11940 4325 11942
rect 4349 11940 4405 11942
rect 4618 11600 4674 11656
rect 4109 10906 4165 10908
rect 4189 10906 4245 10908
rect 4269 10906 4325 10908
rect 4349 10906 4405 10908
rect 4109 10854 4135 10906
rect 4135 10854 4165 10906
rect 4189 10854 4199 10906
rect 4199 10854 4245 10906
rect 4269 10854 4315 10906
rect 4315 10854 4325 10906
rect 4349 10854 4379 10906
rect 4379 10854 4405 10906
rect 4109 10852 4165 10854
rect 4189 10852 4245 10854
rect 4269 10852 4325 10854
rect 4349 10852 4405 10854
rect 4109 9818 4165 9820
rect 4189 9818 4245 9820
rect 4269 9818 4325 9820
rect 4349 9818 4405 9820
rect 4109 9766 4135 9818
rect 4135 9766 4165 9818
rect 4189 9766 4199 9818
rect 4199 9766 4245 9818
rect 4269 9766 4315 9818
rect 4315 9766 4325 9818
rect 4349 9766 4379 9818
rect 4379 9766 4405 9818
rect 4109 9764 4165 9766
rect 4189 9764 4245 9766
rect 4269 9764 4325 9766
rect 4349 9764 4405 9766
rect 4109 8730 4165 8732
rect 4189 8730 4245 8732
rect 4269 8730 4325 8732
rect 4349 8730 4405 8732
rect 4109 8678 4135 8730
rect 4135 8678 4165 8730
rect 4189 8678 4199 8730
rect 4199 8678 4245 8730
rect 4269 8678 4315 8730
rect 4315 8678 4325 8730
rect 4349 8678 4379 8730
rect 4379 8678 4405 8730
rect 4109 8676 4165 8678
rect 4189 8676 4245 8678
rect 4269 8676 4325 8678
rect 4349 8676 4405 8678
rect 4434 8064 4490 8120
rect 4109 7642 4165 7644
rect 4189 7642 4245 7644
rect 4269 7642 4325 7644
rect 4349 7642 4405 7644
rect 4109 7590 4135 7642
rect 4135 7590 4165 7642
rect 4189 7590 4199 7642
rect 4199 7590 4245 7642
rect 4269 7590 4315 7642
rect 4315 7590 4325 7642
rect 4349 7590 4379 7642
rect 4379 7590 4405 7642
rect 4109 7588 4165 7590
rect 4189 7588 4245 7590
rect 4269 7588 4325 7590
rect 4349 7588 4405 7590
rect 4109 6554 4165 6556
rect 4189 6554 4245 6556
rect 4269 6554 4325 6556
rect 4349 6554 4405 6556
rect 4109 6502 4135 6554
rect 4135 6502 4165 6554
rect 4189 6502 4199 6554
rect 4199 6502 4245 6554
rect 4269 6502 4315 6554
rect 4315 6502 4325 6554
rect 4349 6502 4379 6554
rect 4379 6502 4405 6554
rect 4109 6500 4165 6502
rect 4189 6500 4245 6502
rect 4269 6500 4325 6502
rect 4349 6500 4405 6502
rect 4109 5466 4165 5468
rect 4189 5466 4245 5468
rect 4269 5466 4325 5468
rect 4349 5466 4405 5468
rect 4109 5414 4135 5466
rect 4135 5414 4165 5466
rect 4189 5414 4199 5466
rect 4199 5414 4245 5466
rect 4269 5414 4315 5466
rect 4315 5414 4325 5466
rect 4349 5414 4379 5466
rect 4379 5414 4405 5466
rect 4109 5412 4165 5414
rect 4189 5412 4245 5414
rect 4269 5412 4325 5414
rect 4349 5412 4405 5414
rect 4109 4378 4165 4380
rect 4189 4378 4245 4380
rect 4269 4378 4325 4380
rect 4349 4378 4405 4380
rect 4109 4326 4135 4378
rect 4135 4326 4165 4378
rect 4189 4326 4199 4378
rect 4199 4326 4245 4378
rect 4269 4326 4315 4378
rect 4315 4326 4325 4378
rect 4349 4326 4379 4378
rect 4379 4326 4405 4378
rect 4109 4324 4165 4326
rect 4189 4324 4245 4326
rect 4269 4324 4325 4326
rect 4349 4324 4405 4326
rect 4109 3290 4165 3292
rect 4189 3290 4245 3292
rect 4269 3290 4325 3292
rect 4349 3290 4405 3292
rect 4109 3238 4135 3290
rect 4135 3238 4165 3290
rect 4189 3238 4199 3290
rect 4199 3238 4245 3290
rect 4269 3238 4315 3290
rect 4315 3238 4325 3290
rect 4349 3238 4379 3290
rect 4379 3238 4405 3290
rect 4109 3236 4165 3238
rect 4189 3236 4245 3238
rect 4269 3236 4325 3238
rect 4349 3236 4405 3238
rect 4109 2202 4165 2204
rect 4189 2202 4245 2204
rect 4269 2202 4325 2204
rect 4349 2202 4405 2204
rect 4109 2150 4135 2202
rect 4135 2150 4165 2202
rect 4189 2150 4199 2202
rect 4199 2150 4245 2202
rect 4269 2150 4315 2202
rect 4315 2150 4325 2202
rect 4349 2150 4379 2202
rect 4379 2150 4405 2202
rect 4109 2148 4165 2150
rect 4189 2148 4245 2150
rect 4269 2148 4325 2150
rect 4349 2148 4405 2150
rect 10415 14170 10471 14172
rect 10495 14170 10551 14172
rect 10575 14170 10631 14172
rect 10655 14170 10711 14172
rect 10415 14118 10441 14170
rect 10441 14118 10471 14170
rect 10495 14118 10505 14170
rect 10505 14118 10551 14170
rect 10575 14118 10621 14170
rect 10621 14118 10631 14170
rect 10655 14118 10685 14170
rect 10685 14118 10711 14170
rect 10415 14116 10471 14118
rect 10495 14116 10551 14118
rect 10575 14116 10631 14118
rect 10655 14116 10711 14118
rect 7262 13626 7318 13628
rect 7342 13626 7398 13628
rect 7422 13626 7478 13628
rect 7502 13626 7558 13628
rect 7262 13574 7288 13626
rect 7288 13574 7318 13626
rect 7342 13574 7352 13626
rect 7352 13574 7398 13626
rect 7422 13574 7468 13626
rect 7468 13574 7478 13626
rect 7502 13574 7532 13626
rect 7532 13574 7558 13626
rect 7262 13572 7318 13574
rect 7342 13572 7398 13574
rect 7422 13572 7478 13574
rect 7502 13572 7558 13574
rect 7262 12538 7318 12540
rect 7342 12538 7398 12540
rect 7422 12538 7478 12540
rect 7502 12538 7558 12540
rect 7262 12486 7288 12538
rect 7288 12486 7318 12538
rect 7342 12486 7352 12538
rect 7352 12486 7398 12538
rect 7422 12486 7468 12538
rect 7468 12486 7478 12538
rect 7502 12486 7532 12538
rect 7532 12486 7558 12538
rect 7262 12484 7318 12486
rect 7342 12484 7398 12486
rect 7422 12484 7478 12486
rect 7502 12484 7558 12486
rect 7262 11450 7318 11452
rect 7342 11450 7398 11452
rect 7422 11450 7478 11452
rect 7502 11450 7558 11452
rect 7262 11398 7288 11450
rect 7288 11398 7318 11450
rect 7342 11398 7352 11450
rect 7352 11398 7398 11450
rect 7422 11398 7468 11450
rect 7468 11398 7478 11450
rect 7502 11398 7532 11450
rect 7532 11398 7558 11450
rect 7262 11396 7318 11398
rect 7342 11396 7398 11398
rect 7422 11396 7478 11398
rect 7502 11396 7558 11398
rect 7262 10362 7318 10364
rect 7342 10362 7398 10364
rect 7422 10362 7478 10364
rect 7502 10362 7558 10364
rect 7262 10310 7288 10362
rect 7288 10310 7318 10362
rect 7342 10310 7352 10362
rect 7352 10310 7398 10362
rect 7422 10310 7468 10362
rect 7468 10310 7478 10362
rect 7502 10310 7532 10362
rect 7532 10310 7558 10362
rect 7262 10308 7318 10310
rect 7342 10308 7398 10310
rect 7422 10308 7478 10310
rect 7502 10308 7558 10310
rect 7262 9274 7318 9276
rect 7342 9274 7398 9276
rect 7422 9274 7478 9276
rect 7502 9274 7558 9276
rect 7262 9222 7288 9274
rect 7288 9222 7318 9274
rect 7342 9222 7352 9274
rect 7352 9222 7398 9274
rect 7422 9222 7468 9274
rect 7468 9222 7478 9274
rect 7502 9222 7532 9274
rect 7532 9222 7558 9274
rect 7262 9220 7318 9222
rect 7342 9220 7398 9222
rect 7422 9220 7478 9222
rect 7502 9220 7558 9222
rect 7262 8186 7318 8188
rect 7342 8186 7398 8188
rect 7422 8186 7478 8188
rect 7502 8186 7558 8188
rect 7262 8134 7288 8186
rect 7288 8134 7318 8186
rect 7342 8134 7352 8186
rect 7352 8134 7398 8186
rect 7422 8134 7468 8186
rect 7468 8134 7478 8186
rect 7502 8134 7532 8186
rect 7532 8134 7558 8186
rect 7262 8132 7318 8134
rect 7342 8132 7398 8134
rect 7422 8132 7478 8134
rect 7502 8132 7558 8134
rect 7262 7098 7318 7100
rect 7342 7098 7398 7100
rect 7422 7098 7478 7100
rect 7502 7098 7558 7100
rect 7262 7046 7288 7098
rect 7288 7046 7318 7098
rect 7342 7046 7352 7098
rect 7352 7046 7398 7098
rect 7422 7046 7468 7098
rect 7468 7046 7478 7098
rect 7502 7046 7532 7098
rect 7532 7046 7558 7098
rect 7262 7044 7318 7046
rect 7342 7044 7398 7046
rect 7422 7044 7478 7046
rect 7502 7044 7558 7046
rect 6734 1944 6790 2000
rect 7262 6010 7318 6012
rect 7342 6010 7398 6012
rect 7422 6010 7478 6012
rect 7502 6010 7558 6012
rect 7262 5958 7288 6010
rect 7288 5958 7318 6010
rect 7342 5958 7352 6010
rect 7352 5958 7398 6010
rect 7422 5958 7468 6010
rect 7468 5958 7478 6010
rect 7502 5958 7532 6010
rect 7532 5958 7558 6010
rect 7262 5956 7318 5958
rect 7342 5956 7398 5958
rect 7422 5956 7478 5958
rect 7502 5956 7558 5958
rect 7262 4922 7318 4924
rect 7342 4922 7398 4924
rect 7422 4922 7478 4924
rect 7502 4922 7558 4924
rect 7262 4870 7288 4922
rect 7288 4870 7318 4922
rect 7342 4870 7352 4922
rect 7352 4870 7398 4922
rect 7422 4870 7468 4922
rect 7468 4870 7478 4922
rect 7502 4870 7532 4922
rect 7532 4870 7558 4922
rect 7262 4868 7318 4870
rect 7342 4868 7398 4870
rect 7422 4868 7478 4870
rect 7502 4868 7558 4870
rect 7262 3834 7318 3836
rect 7342 3834 7398 3836
rect 7422 3834 7478 3836
rect 7502 3834 7558 3836
rect 7262 3782 7288 3834
rect 7288 3782 7318 3834
rect 7342 3782 7352 3834
rect 7352 3782 7398 3834
rect 7422 3782 7468 3834
rect 7468 3782 7478 3834
rect 7502 3782 7532 3834
rect 7532 3782 7558 3834
rect 7262 3780 7318 3782
rect 7342 3780 7398 3782
rect 7422 3780 7478 3782
rect 7502 3780 7558 3782
rect 7262 2746 7318 2748
rect 7342 2746 7398 2748
rect 7422 2746 7478 2748
rect 7502 2746 7558 2748
rect 7262 2694 7288 2746
rect 7288 2694 7318 2746
rect 7342 2694 7352 2746
rect 7352 2694 7398 2746
rect 7422 2694 7468 2746
rect 7468 2694 7478 2746
rect 7502 2694 7532 2746
rect 7532 2694 7558 2746
rect 7262 2692 7318 2694
rect 7342 2692 7398 2694
rect 7422 2692 7478 2694
rect 7502 2692 7558 2694
rect 10415 13082 10471 13084
rect 10495 13082 10551 13084
rect 10575 13082 10631 13084
rect 10655 13082 10711 13084
rect 10415 13030 10441 13082
rect 10441 13030 10471 13082
rect 10495 13030 10505 13082
rect 10505 13030 10551 13082
rect 10575 13030 10621 13082
rect 10621 13030 10631 13082
rect 10655 13030 10685 13082
rect 10685 13030 10711 13082
rect 10415 13028 10471 13030
rect 10495 13028 10551 13030
rect 10575 13028 10631 13030
rect 10655 13028 10711 13030
rect 10415 11994 10471 11996
rect 10495 11994 10551 11996
rect 10575 11994 10631 11996
rect 10655 11994 10711 11996
rect 10415 11942 10441 11994
rect 10441 11942 10471 11994
rect 10495 11942 10505 11994
rect 10505 11942 10551 11994
rect 10575 11942 10621 11994
rect 10621 11942 10631 11994
rect 10655 11942 10685 11994
rect 10685 11942 10711 11994
rect 10415 11940 10471 11942
rect 10495 11940 10551 11942
rect 10575 11940 10631 11942
rect 10655 11940 10711 11942
rect 10415 10906 10471 10908
rect 10495 10906 10551 10908
rect 10575 10906 10631 10908
rect 10655 10906 10711 10908
rect 10415 10854 10441 10906
rect 10441 10854 10471 10906
rect 10495 10854 10505 10906
rect 10505 10854 10551 10906
rect 10575 10854 10621 10906
rect 10621 10854 10631 10906
rect 10655 10854 10685 10906
rect 10685 10854 10711 10906
rect 10415 10852 10471 10854
rect 10495 10852 10551 10854
rect 10575 10852 10631 10854
rect 10655 10852 10711 10854
rect 10415 9818 10471 9820
rect 10495 9818 10551 9820
rect 10575 9818 10631 9820
rect 10655 9818 10711 9820
rect 10415 9766 10441 9818
rect 10441 9766 10471 9818
rect 10495 9766 10505 9818
rect 10505 9766 10551 9818
rect 10575 9766 10621 9818
rect 10621 9766 10631 9818
rect 10655 9766 10685 9818
rect 10685 9766 10711 9818
rect 10415 9764 10471 9766
rect 10495 9764 10551 9766
rect 10575 9764 10631 9766
rect 10655 9764 10711 9766
rect 13569 17978 13625 17980
rect 13649 17978 13705 17980
rect 13729 17978 13785 17980
rect 13809 17978 13865 17980
rect 13569 17926 13595 17978
rect 13595 17926 13625 17978
rect 13649 17926 13659 17978
rect 13659 17926 13705 17978
rect 13729 17926 13775 17978
rect 13775 17926 13785 17978
rect 13809 17926 13839 17978
rect 13839 17926 13865 17978
rect 13569 17924 13625 17926
rect 13649 17924 13705 17926
rect 13729 17924 13785 17926
rect 13809 17924 13865 17926
rect 12622 17740 12678 17776
rect 12622 17720 12624 17740
rect 12624 17720 12676 17740
rect 12676 17720 12678 17740
rect 13569 16890 13625 16892
rect 13649 16890 13705 16892
rect 13729 16890 13785 16892
rect 13809 16890 13865 16892
rect 13569 16838 13595 16890
rect 13595 16838 13625 16890
rect 13649 16838 13659 16890
rect 13659 16838 13705 16890
rect 13729 16838 13775 16890
rect 13775 16838 13785 16890
rect 13809 16838 13839 16890
rect 13839 16838 13865 16890
rect 13569 16836 13625 16838
rect 13649 16836 13705 16838
rect 13729 16836 13785 16838
rect 13809 16836 13865 16838
rect 13569 15802 13625 15804
rect 13649 15802 13705 15804
rect 13729 15802 13785 15804
rect 13809 15802 13865 15804
rect 13569 15750 13595 15802
rect 13595 15750 13625 15802
rect 13649 15750 13659 15802
rect 13659 15750 13705 15802
rect 13729 15750 13775 15802
rect 13775 15750 13785 15802
rect 13809 15750 13839 15802
rect 13839 15750 13865 15802
rect 13569 15748 13625 15750
rect 13649 15748 13705 15750
rect 13729 15748 13785 15750
rect 13809 15748 13865 15750
rect 13569 14714 13625 14716
rect 13649 14714 13705 14716
rect 13729 14714 13785 14716
rect 13809 14714 13865 14716
rect 13569 14662 13595 14714
rect 13595 14662 13625 14714
rect 13649 14662 13659 14714
rect 13659 14662 13705 14714
rect 13729 14662 13775 14714
rect 13775 14662 13785 14714
rect 13809 14662 13839 14714
rect 13839 14662 13865 14714
rect 13569 14660 13625 14662
rect 13649 14660 13705 14662
rect 13729 14660 13785 14662
rect 13809 14660 13865 14662
rect 13569 13626 13625 13628
rect 13649 13626 13705 13628
rect 13729 13626 13785 13628
rect 13809 13626 13865 13628
rect 13569 13574 13595 13626
rect 13595 13574 13625 13626
rect 13649 13574 13659 13626
rect 13659 13574 13705 13626
rect 13729 13574 13775 13626
rect 13775 13574 13785 13626
rect 13809 13574 13839 13626
rect 13839 13574 13865 13626
rect 13569 13572 13625 13574
rect 13649 13572 13705 13574
rect 13729 13572 13785 13574
rect 13809 13572 13865 13574
rect 13569 12538 13625 12540
rect 13649 12538 13705 12540
rect 13729 12538 13785 12540
rect 13809 12538 13865 12540
rect 13569 12486 13595 12538
rect 13595 12486 13625 12538
rect 13649 12486 13659 12538
rect 13659 12486 13705 12538
rect 13729 12486 13775 12538
rect 13775 12486 13785 12538
rect 13809 12486 13839 12538
rect 13839 12486 13865 12538
rect 13569 12484 13625 12486
rect 13649 12484 13705 12486
rect 13729 12484 13785 12486
rect 13809 12484 13865 12486
rect 16722 18522 16778 18524
rect 16802 18522 16858 18524
rect 16882 18522 16938 18524
rect 16962 18522 17018 18524
rect 16722 18470 16748 18522
rect 16748 18470 16778 18522
rect 16802 18470 16812 18522
rect 16812 18470 16858 18522
rect 16882 18470 16928 18522
rect 16928 18470 16938 18522
rect 16962 18470 16992 18522
rect 16992 18470 17018 18522
rect 16722 18468 16778 18470
rect 16802 18468 16858 18470
rect 16882 18468 16938 18470
rect 16962 18468 17018 18470
rect 18510 20304 18566 20360
rect 18418 19080 18474 19136
rect 15474 16904 15530 16960
rect 16722 17434 16778 17436
rect 16802 17434 16858 17436
rect 16882 17434 16938 17436
rect 16962 17434 17018 17436
rect 16722 17382 16748 17434
rect 16748 17382 16778 17434
rect 16802 17382 16812 17434
rect 16812 17382 16858 17434
rect 16882 17382 16928 17434
rect 16928 17382 16938 17434
rect 16962 17382 16992 17434
rect 16992 17382 17018 17434
rect 16722 17380 16778 17382
rect 16802 17380 16858 17382
rect 16882 17380 16938 17382
rect 16962 17380 17018 17382
rect 15198 11600 15254 11656
rect 13569 11450 13625 11452
rect 13649 11450 13705 11452
rect 13729 11450 13785 11452
rect 13809 11450 13865 11452
rect 13569 11398 13595 11450
rect 13595 11398 13625 11450
rect 13649 11398 13659 11450
rect 13659 11398 13705 11450
rect 13729 11398 13775 11450
rect 13775 11398 13785 11450
rect 13809 11398 13839 11450
rect 13839 11398 13865 11450
rect 13569 11396 13625 11398
rect 13649 11396 13705 11398
rect 13729 11396 13785 11398
rect 13809 11396 13865 11398
rect 14830 11192 14886 11248
rect 13569 10362 13625 10364
rect 13649 10362 13705 10364
rect 13729 10362 13785 10364
rect 13809 10362 13865 10364
rect 13569 10310 13595 10362
rect 13595 10310 13625 10362
rect 13649 10310 13659 10362
rect 13659 10310 13705 10362
rect 13729 10310 13775 10362
rect 13775 10310 13785 10362
rect 13809 10310 13839 10362
rect 13839 10310 13865 10362
rect 13569 10308 13625 10310
rect 13649 10308 13705 10310
rect 13729 10308 13785 10310
rect 13809 10308 13865 10310
rect 14462 9968 14518 10024
rect 13569 9274 13625 9276
rect 13649 9274 13705 9276
rect 13729 9274 13785 9276
rect 13809 9274 13865 9276
rect 13569 9222 13595 9274
rect 13595 9222 13625 9274
rect 13649 9222 13659 9274
rect 13659 9222 13705 9274
rect 13729 9222 13775 9274
rect 13775 9222 13785 9274
rect 13809 9222 13839 9274
rect 13839 9222 13865 9274
rect 13569 9220 13625 9222
rect 13649 9220 13705 9222
rect 13729 9220 13785 9222
rect 13809 9220 13865 9222
rect 10415 8730 10471 8732
rect 10495 8730 10551 8732
rect 10575 8730 10631 8732
rect 10655 8730 10711 8732
rect 10415 8678 10441 8730
rect 10441 8678 10471 8730
rect 10495 8678 10505 8730
rect 10505 8678 10551 8730
rect 10575 8678 10621 8730
rect 10621 8678 10631 8730
rect 10655 8678 10685 8730
rect 10685 8678 10711 8730
rect 10415 8676 10471 8678
rect 10495 8676 10551 8678
rect 10575 8676 10631 8678
rect 10655 8676 10711 8678
rect 13569 8186 13625 8188
rect 13649 8186 13705 8188
rect 13729 8186 13785 8188
rect 13809 8186 13865 8188
rect 13569 8134 13595 8186
rect 13595 8134 13625 8186
rect 13649 8134 13659 8186
rect 13659 8134 13705 8186
rect 13729 8134 13775 8186
rect 13775 8134 13785 8186
rect 13809 8134 13839 8186
rect 13839 8134 13865 8186
rect 13569 8132 13625 8134
rect 13649 8132 13705 8134
rect 13729 8132 13785 8134
rect 13809 8132 13865 8134
rect 10415 7642 10471 7644
rect 10495 7642 10551 7644
rect 10575 7642 10631 7644
rect 10655 7642 10711 7644
rect 10415 7590 10441 7642
rect 10441 7590 10471 7642
rect 10495 7590 10505 7642
rect 10505 7590 10551 7642
rect 10575 7590 10621 7642
rect 10621 7590 10631 7642
rect 10655 7590 10685 7642
rect 10685 7590 10711 7642
rect 10415 7588 10471 7590
rect 10495 7588 10551 7590
rect 10575 7588 10631 7590
rect 10655 7588 10711 7590
rect 16722 16346 16778 16348
rect 16802 16346 16858 16348
rect 16882 16346 16938 16348
rect 16962 16346 17018 16348
rect 16722 16294 16748 16346
rect 16748 16294 16778 16346
rect 16802 16294 16812 16346
rect 16812 16294 16858 16346
rect 16882 16294 16928 16346
rect 16928 16294 16938 16346
rect 16962 16294 16992 16346
rect 16992 16294 17018 16346
rect 16722 16292 16778 16294
rect 16802 16292 16858 16294
rect 16882 16292 16938 16294
rect 16962 16292 17018 16294
rect 16722 15258 16778 15260
rect 16802 15258 16858 15260
rect 16882 15258 16938 15260
rect 16962 15258 17018 15260
rect 16722 15206 16748 15258
rect 16748 15206 16778 15258
rect 16802 15206 16812 15258
rect 16812 15206 16858 15258
rect 16882 15206 16928 15258
rect 16928 15206 16938 15258
rect 16962 15206 16992 15258
rect 16992 15206 17018 15258
rect 16722 15204 16778 15206
rect 16802 15204 16858 15206
rect 16882 15204 16938 15206
rect 16962 15204 17018 15206
rect 16486 14864 16542 14920
rect 16722 14170 16778 14172
rect 16802 14170 16858 14172
rect 16882 14170 16938 14172
rect 16962 14170 17018 14172
rect 16722 14118 16748 14170
rect 16748 14118 16778 14170
rect 16802 14118 16812 14170
rect 16812 14118 16858 14170
rect 16882 14118 16928 14170
rect 16928 14118 16938 14170
rect 16962 14118 16992 14170
rect 16992 14118 17018 14170
rect 16722 14116 16778 14118
rect 16802 14116 16858 14118
rect 16882 14116 16938 14118
rect 16962 14116 17018 14118
rect 16486 13640 16542 13696
rect 16722 13082 16778 13084
rect 16802 13082 16858 13084
rect 16882 13082 16938 13084
rect 16962 13082 17018 13084
rect 16722 13030 16748 13082
rect 16748 13030 16778 13082
rect 16802 13030 16812 13082
rect 16812 13030 16858 13082
rect 16882 13030 16928 13082
rect 16928 13030 16938 13082
rect 16962 13030 16992 13082
rect 16992 13030 17018 13082
rect 16722 13028 16778 13030
rect 16802 13028 16858 13030
rect 16882 13028 16938 13030
rect 16962 13028 17018 13030
rect 17130 12960 17186 13016
rect 16722 11994 16778 11996
rect 16802 11994 16858 11996
rect 16882 11994 16938 11996
rect 16962 11994 17018 11996
rect 16722 11942 16748 11994
rect 16748 11942 16778 11994
rect 16802 11942 16812 11994
rect 16812 11942 16858 11994
rect 16882 11942 16928 11994
rect 16928 11942 16938 11994
rect 16962 11942 16992 11994
rect 16992 11942 17018 11994
rect 16722 11940 16778 11942
rect 16802 11940 16858 11942
rect 16882 11940 16938 11942
rect 16962 11940 17018 11942
rect 16722 10906 16778 10908
rect 16802 10906 16858 10908
rect 16882 10906 16938 10908
rect 16962 10906 17018 10908
rect 16722 10854 16748 10906
rect 16748 10854 16778 10906
rect 16802 10854 16812 10906
rect 16812 10854 16858 10906
rect 16882 10854 16928 10906
rect 16928 10854 16938 10906
rect 16962 10854 16992 10906
rect 16992 10854 17018 10906
rect 16722 10852 16778 10854
rect 16802 10852 16858 10854
rect 16882 10852 16938 10854
rect 16962 10852 17018 10854
rect 16722 9818 16778 9820
rect 16802 9818 16858 9820
rect 16882 9818 16938 9820
rect 16962 9818 17018 9820
rect 16722 9766 16748 9818
rect 16748 9766 16778 9818
rect 16802 9766 16812 9818
rect 16812 9766 16858 9818
rect 16882 9766 16928 9818
rect 16928 9766 16938 9818
rect 16962 9766 16992 9818
rect 16992 9766 17018 9818
rect 16722 9764 16778 9766
rect 16802 9764 16858 9766
rect 16882 9764 16938 9766
rect 16962 9764 17018 9766
rect 16722 8730 16778 8732
rect 16802 8730 16858 8732
rect 16882 8730 16938 8732
rect 16962 8730 17018 8732
rect 16722 8678 16748 8730
rect 16748 8678 16778 8730
rect 16802 8678 16812 8730
rect 16812 8678 16858 8730
rect 16882 8678 16928 8730
rect 16928 8678 16938 8730
rect 16962 8678 16992 8730
rect 16992 8678 17018 8730
rect 16722 8676 16778 8678
rect 16802 8676 16858 8678
rect 16882 8676 16938 8678
rect 16962 8676 17018 8678
rect 15474 7928 15530 7984
rect 13569 7098 13625 7100
rect 13649 7098 13705 7100
rect 13729 7098 13785 7100
rect 13809 7098 13865 7100
rect 13569 7046 13595 7098
rect 13595 7046 13625 7098
rect 13649 7046 13659 7098
rect 13659 7046 13705 7098
rect 13729 7046 13775 7098
rect 13775 7046 13785 7098
rect 13809 7046 13839 7098
rect 13839 7046 13865 7098
rect 13569 7044 13625 7046
rect 13649 7044 13705 7046
rect 13729 7044 13785 7046
rect 13809 7044 13865 7046
rect 10415 6554 10471 6556
rect 10495 6554 10551 6556
rect 10575 6554 10631 6556
rect 10655 6554 10711 6556
rect 10415 6502 10441 6554
rect 10441 6502 10471 6554
rect 10495 6502 10505 6554
rect 10505 6502 10551 6554
rect 10575 6502 10621 6554
rect 10621 6502 10631 6554
rect 10655 6502 10685 6554
rect 10685 6502 10711 6554
rect 10415 6500 10471 6502
rect 10495 6500 10551 6502
rect 10575 6500 10631 6502
rect 10655 6500 10711 6502
rect 10415 5466 10471 5468
rect 10495 5466 10551 5468
rect 10575 5466 10631 5468
rect 10655 5466 10711 5468
rect 10415 5414 10441 5466
rect 10441 5414 10471 5466
rect 10495 5414 10505 5466
rect 10505 5414 10551 5466
rect 10575 5414 10621 5466
rect 10621 5414 10631 5466
rect 10655 5414 10685 5466
rect 10685 5414 10711 5466
rect 10415 5412 10471 5414
rect 10495 5412 10551 5414
rect 10575 5412 10631 5414
rect 10655 5412 10711 5414
rect 10415 4378 10471 4380
rect 10495 4378 10551 4380
rect 10575 4378 10631 4380
rect 10655 4378 10711 4380
rect 10415 4326 10441 4378
rect 10441 4326 10471 4378
rect 10495 4326 10505 4378
rect 10505 4326 10551 4378
rect 10575 4326 10621 4378
rect 10621 4326 10631 4378
rect 10655 4326 10685 4378
rect 10685 4326 10711 4378
rect 10415 4324 10471 4326
rect 10495 4324 10551 4326
rect 10575 4324 10631 4326
rect 10655 4324 10711 4326
rect 10415 3290 10471 3292
rect 10495 3290 10551 3292
rect 10575 3290 10631 3292
rect 10655 3290 10711 3292
rect 10415 3238 10441 3290
rect 10441 3238 10471 3290
rect 10495 3238 10505 3290
rect 10505 3238 10551 3290
rect 10575 3238 10621 3290
rect 10621 3238 10631 3290
rect 10655 3238 10685 3290
rect 10685 3238 10711 3290
rect 10415 3236 10471 3238
rect 10495 3236 10551 3238
rect 10575 3236 10631 3238
rect 10655 3236 10711 3238
rect 12346 5072 12402 5128
rect 10415 2202 10471 2204
rect 10495 2202 10551 2204
rect 10575 2202 10631 2204
rect 10655 2202 10711 2204
rect 10415 2150 10441 2202
rect 10441 2150 10471 2202
rect 10495 2150 10505 2202
rect 10505 2150 10551 2202
rect 10575 2150 10621 2202
rect 10621 2150 10631 2202
rect 10655 2150 10685 2202
rect 10685 2150 10711 2202
rect 10415 2148 10471 2150
rect 10495 2148 10551 2150
rect 10575 2148 10631 2150
rect 10655 2148 10711 2150
rect 10414 40 10470 96
rect 13569 6010 13625 6012
rect 13649 6010 13705 6012
rect 13729 6010 13785 6012
rect 13809 6010 13865 6012
rect 13569 5958 13595 6010
rect 13595 5958 13625 6010
rect 13649 5958 13659 6010
rect 13659 5958 13705 6010
rect 13729 5958 13775 6010
rect 13775 5958 13785 6010
rect 13809 5958 13839 6010
rect 13839 5958 13865 6010
rect 13569 5956 13625 5958
rect 13649 5956 13705 5958
rect 13729 5956 13785 5958
rect 13809 5956 13865 5958
rect 13569 4922 13625 4924
rect 13649 4922 13705 4924
rect 13729 4922 13785 4924
rect 13809 4922 13865 4924
rect 13569 4870 13595 4922
rect 13595 4870 13625 4922
rect 13649 4870 13659 4922
rect 13659 4870 13705 4922
rect 13729 4870 13775 4922
rect 13775 4870 13785 4922
rect 13809 4870 13839 4922
rect 13839 4870 13865 4922
rect 13569 4868 13625 4870
rect 13649 4868 13705 4870
rect 13729 4868 13785 4870
rect 13809 4868 13865 4870
rect 13569 3834 13625 3836
rect 13649 3834 13705 3836
rect 13729 3834 13785 3836
rect 13809 3834 13865 3836
rect 13569 3782 13595 3834
rect 13595 3782 13625 3834
rect 13649 3782 13659 3834
rect 13659 3782 13705 3834
rect 13729 3782 13775 3834
rect 13775 3782 13785 3834
rect 13809 3782 13839 3834
rect 13839 3782 13865 3834
rect 13569 3780 13625 3782
rect 13649 3780 13705 3782
rect 13729 3780 13785 3782
rect 13809 3780 13865 3782
rect 13569 2746 13625 2748
rect 13649 2746 13705 2748
rect 13729 2746 13785 2748
rect 13809 2746 13865 2748
rect 13569 2694 13595 2746
rect 13595 2694 13625 2746
rect 13649 2694 13659 2746
rect 13659 2694 13705 2746
rect 13729 2694 13775 2746
rect 13775 2694 13785 2746
rect 13809 2694 13839 2746
rect 13839 2694 13865 2746
rect 13569 2692 13625 2694
rect 13649 2692 13705 2694
rect 13729 2692 13785 2694
rect 13809 2692 13865 2694
rect 14002 1944 14058 2000
rect 16722 7642 16778 7644
rect 16802 7642 16858 7644
rect 16882 7642 16938 7644
rect 16962 7642 17018 7644
rect 16722 7590 16748 7642
rect 16748 7590 16778 7642
rect 16802 7590 16812 7642
rect 16812 7590 16858 7642
rect 16882 7590 16928 7642
rect 16928 7590 16938 7642
rect 16962 7590 16992 7642
rect 16992 7590 17018 7642
rect 16722 7588 16778 7590
rect 16802 7588 16858 7590
rect 16882 7588 16938 7590
rect 16962 7588 17018 7590
rect 16722 6554 16778 6556
rect 16802 6554 16858 6556
rect 16882 6554 16938 6556
rect 16962 6554 17018 6556
rect 16722 6502 16748 6554
rect 16748 6502 16778 6554
rect 16802 6502 16812 6554
rect 16812 6502 16858 6554
rect 16882 6502 16928 6554
rect 16928 6502 16938 6554
rect 16962 6502 16992 6554
rect 16992 6502 17018 6554
rect 16722 6500 16778 6502
rect 16802 6500 16858 6502
rect 16882 6500 16938 6502
rect 16962 6500 17018 6502
rect 18418 9152 18474 9208
rect 17130 6432 17186 6488
rect 17038 6024 17094 6080
rect 16722 5466 16778 5468
rect 16802 5466 16858 5468
rect 16882 5466 16938 5468
rect 16962 5466 17018 5468
rect 16722 5414 16748 5466
rect 16748 5414 16778 5466
rect 16802 5414 16812 5466
rect 16812 5414 16858 5466
rect 16882 5414 16928 5466
rect 16928 5414 16938 5466
rect 16962 5414 16992 5466
rect 16992 5414 17018 5466
rect 16722 5412 16778 5414
rect 16802 5412 16858 5414
rect 16882 5412 16938 5414
rect 16962 5412 17018 5414
rect 16722 4378 16778 4380
rect 16802 4378 16858 4380
rect 16882 4378 16938 4380
rect 16962 4378 17018 4380
rect 16722 4326 16748 4378
rect 16748 4326 16778 4378
rect 16802 4326 16812 4378
rect 16812 4326 16858 4378
rect 16882 4326 16928 4378
rect 16928 4326 16938 4378
rect 16962 4326 16992 4378
rect 16992 4326 17018 4378
rect 16722 4324 16778 4326
rect 16802 4324 16858 4326
rect 16882 4324 16938 4326
rect 16962 4324 17018 4326
rect 16722 3290 16778 3292
rect 16802 3290 16858 3292
rect 16882 3290 16938 3292
rect 16962 3290 17018 3292
rect 16722 3238 16748 3290
rect 16748 3238 16778 3290
rect 16802 3238 16812 3290
rect 16812 3238 16858 3290
rect 16882 3238 16928 3290
rect 16928 3238 16938 3290
rect 16962 3238 16992 3290
rect 16992 3238 17018 3290
rect 16722 3236 16778 3238
rect 16802 3236 16858 3238
rect 16882 3236 16938 3238
rect 16962 3236 17018 3238
rect 16722 2202 16778 2204
rect 16802 2202 16858 2204
rect 16882 2202 16938 2204
rect 16962 2202 17018 2204
rect 16722 2150 16748 2202
rect 16748 2150 16778 2202
rect 16802 2150 16812 2202
rect 16812 2150 16858 2202
rect 16882 2150 16928 2202
rect 16928 2150 16938 2202
rect 16962 2150 16992 2202
rect 16992 2150 17018 2202
rect 16722 2148 16778 2150
rect 16802 2148 16858 2150
rect 16882 2148 16938 2150
rect 16962 2148 17018 2150
<< metal3 >>
rect 18439 20360 18919 20392
rect 18439 20304 18510 20360
rect 18566 20304 18919 20360
rect 18439 20272 18919 20304
rect 0 20000 480 20120
rect 62 19546 122 20000
rect 1209 19546 1275 19549
rect 62 19544 1275 19546
rect 62 19488 1214 19544
rect 1270 19488 1275 19544
rect 62 19486 1275 19488
rect 1209 19483 1275 19486
rect 18439 19141 18919 19168
rect 18413 19138 18919 19141
rect 18332 19136 18919 19138
rect 18332 19080 18418 19136
rect 18474 19080 18919 19136
rect 18332 19078 18919 19080
rect 18413 19075 18919 19078
rect 18439 19048 18919 19075
rect 4097 18528 4417 18529
rect 4097 18464 4105 18528
rect 4169 18464 4185 18528
rect 4249 18464 4265 18528
rect 4329 18464 4345 18528
rect 4409 18464 4417 18528
rect 4097 18463 4417 18464
rect 10403 18528 10723 18529
rect 10403 18464 10411 18528
rect 10475 18464 10491 18528
rect 10555 18464 10571 18528
rect 10635 18464 10651 18528
rect 10715 18464 10723 18528
rect 10403 18463 10723 18464
rect 16710 18528 17030 18529
rect 16710 18464 16718 18528
rect 16782 18464 16798 18528
rect 16862 18464 16878 18528
rect 16942 18464 16958 18528
rect 17022 18464 17030 18528
rect 16710 18463 17030 18464
rect 0 18096 480 18216
rect 7465 18186 7531 18189
rect 7465 18184 18522 18186
rect 7465 18128 7470 18184
rect 7526 18128 18522 18184
rect 7465 18126 18522 18128
rect 7465 18123 7531 18126
rect 62 17642 122 18096
rect 7250 17984 7570 17985
rect 7250 17920 7258 17984
rect 7322 17920 7338 17984
rect 7402 17920 7418 17984
rect 7482 17920 7498 17984
rect 7562 17920 7570 17984
rect 7250 17919 7570 17920
rect 13557 17984 13877 17985
rect 13557 17920 13565 17984
rect 13629 17920 13645 17984
rect 13709 17920 13725 17984
rect 13789 17920 13805 17984
rect 13869 17920 13877 17984
rect 18462 17944 18522 18126
rect 13557 17919 13877 17920
rect 18439 17824 18919 17944
rect 1761 17778 1827 17781
rect 12617 17778 12683 17781
rect 1761 17776 12683 17778
rect 1761 17720 1766 17776
rect 1822 17720 12622 17776
rect 12678 17720 12683 17776
rect 1761 17718 12683 17720
rect 1761 17715 1827 17718
rect 12617 17715 12683 17718
rect 1761 17642 1827 17645
rect 62 17640 1827 17642
rect 62 17584 1766 17640
rect 1822 17584 1827 17640
rect 62 17582 1827 17584
rect 1761 17579 1827 17582
rect 4097 17440 4417 17441
rect 4097 17376 4105 17440
rect 4169 17376 4185 17440
rect 4249 17376 4265 17440
rect 4329 17376 4345 17440
rect 4409 17376 4417 17440
rect 4097 17375 4417 17376
rect 10403 17440 10723 17441
rect 10403 17376 10411 17440
rect 10475 17376 10491 17440
rect 10555 17376 10571 17440
rect 10635 17376 10651 17440
rect 10715 17376 10723 17440
rect 10403 17375 10723 17376
rect 16710 17440 17030 17441
rect 16710 17376 16718 17440
rect 16782 17376 16798 17440
rect 16862 17376 16878 17440
rect 16942 17376 16958 17440
rect 17022 17376 17030 17440
rect 16710 17375 17030 17376
rect 15469 16962 15535 16965
rect 15469 16960 18522 16962
rect 15469 16904 15474 16960
rect 15530 16904 18522 16960
rect 15469 16902 18522 16904
rect 15469 16899 15535 16902
rect 7250 16896 7570 16897
rect 7250 16832 7258 16896
rect 7322 16832 7338 16896
rect 7402 16832 7418 16896
rect 7482 16832 7498 16896
rect 7562 16832 7570 16896
rect 7250 16831 7570 16832
rect 13557 16896 13877 16897
rect 13557 16832 13565 16896
rect 13629 16832 13645 16896
rect 13709 16832 13725 16896
rect 13789 16832 13805 16896
rect 13869 16832 13877 16896
rect 13557 16831 13877 16832
rect 18462 16720 18522 16902
rect 18439 16600 18919 16720
rect 4097 16352 4417 16353
rect 0 16192 480 16312
rect 4097 16288 4105 16352
rect 4169 16288 4185 16352
rect 4249 16288 4265 16352
rect 4329 16288 4345 16352
rect 4409 16288 4417 16352
rect 4097 16287 4417 16288
rect 10403 16352 10723 16353
rect 10403 16288 10411 16352
rect 10475 16288 10491 16352
rect 10555 16288 10571 16352
rect 10635 16288 10651 16352
rect 10715 16288 10723 16352
rect 10403 16287 10723 16288
rect 16710 16352 17030 16353
rect 16710 16288 16718 16352
rect 16782 16288 16798 16352
rect 16862 16288 16878 16352
rect 16942 16288 16958 16352
rect 17022 16288 17030 16352
rect 16710 16287 17030 16288
rect 62 15738 122 16192
rect 7250 15808 7570 15809
rect 7250 15744 7258 15808
rect 7322 15744 7338 15808
rect 7402 15744 7418 15808
rect 7482 15744 7498 15808
rect 7562 15744 7570 15808
rect 7250 15743 7570 15744
rect 13557 15808 13877 15809
rect 13557 15744 13565 15808
rect 13629 15744 13645 15808
rect 13709 15744 13725 15808
rect 13789 15744 13805 15808
rect 13869 15744 13877 15808
rect 13557 15743 13877 15744
rect 3969 15738 4035 15741
rect 62 15736 4035 15738
rect 62 15680 3974 15736
rect 4030 15680 4035 15736
rect 62 15678 4035 15680
rect 3969 15675 4035 15678
rect 18439 15376 18919 15496
rect 4097 15264 4417 15265
rect 4097 15200 4105 15264
rect 4169 15200 4185 15264
rect 4249 15200 4265 15264
rect 4329 15200 4345 15264
rect 4409 15200 4417 15264
rect 4097 15199 4417 15200
rect 10403 15264 10723 15265
rect 10403 15200 10411 15264
rect 10475 15200 10491 15264
rect 10555 15200 10571 15264
rect 10635 15200 10651 15264
rect 10715 15200 10723 15264
rect 10403 15199 10723 15200
rect 16710 15264 17030 15265
rect 16710 15200 16718 15264
rect 16782 15200 16798 15264
rect 16862 15200 16878 15264
rect 16942 15200 16958 15264
rect 17022 15200 17030 15264
rect 16710 15199 17030 15200
rect 16481 14922 16547 14925
rect 18462 14922 18522 15376
rect 16481 14920 18522 14922
rect 16481 14864 16486 14920
rect 16542 14864 18522 14920
rect 16481 14862 18522 14864
rect 16481 14859 16547 14862
rect 7250 14720 7570 14721
rect 7250 14656 7258 14720
rect 7322 14656 7338 14720
rect 7402 14656 7418 14720
rect 7482 14656 7498 14720
rect 7562 14656 7570 14720
rect 7250 14655 7570 14656
rect 13557 14720 13877 14721
rect 13557 14656 13565 14720
rect 13629 14656 13645 14720
rect 13709 14656 13725 14720
rect 13789 14656 13805 14720
rect 13869 14656 13877 14720
rect 13557 14655 13877 14656
rect 0 14376 480 14408
rect 0 14320 110 14376
rect 166 14320 480 14376
rect 0 14288 480 14320
rect 4097 14176 4417 14177
rect 4097 14112 4105 14176
rect 4169 14112 4185 14176
rect 4249 14112 4265 14176
rect 4329 14112 4345 14176
rect 4409 14112 4417 14176
rect 4097 14111 4417 14112
rect 10403 14176 10723 14177
rect 10403 14112 10411 14176
rect 10475 14112 10491 14176
rect 10555 14112 10571 14176
rect 10635 14112 10651 14176
rect 10715 14112 10723 14176
rect 10403 14111 10723 14112
rect 16710 14176 17030 14177
rect 16710 14112 16718 14176
rect 16782 14112 16798 14176
rect 16862 14112 16878 14176
rect 16942 14112 16958 14176
rect 17022 14112 17030 14176
rect 18439 14152 18919 14272
rect 16710 14111 17030 14112
rect 16481 13698 16547 13701
rect 18462 13698 18522 14152
rect 16481 13696 18522 13698
rect 16481 13640 16486 13696
rect 16542 13640 18522 13696
rect 16481 13638 18522 13640
rect 16481 13635 16547 13638
rect 7250 13632 7570 13633
rect 7250 13568 7258 13632
rect 7322 13568 7338 13632
rect 7402 13568 7418 13632
rect 7482 13568 7498 13632
rect 7562 13568 7570 13632
rect 7250 13567 7570 13568
rect 13557 13632 13877 13633
rect 13557 13568 13565 13632
rect 13629 13568 13645 13632
rect 13709 13568 13725 13632
rect 13789 13568 13805 13632
rect 13869 13568 13877 13632
rect 13557 13567 13877 13568
rect 4097 13088 4417 13089
rect 4097 13024 4105 13088
rect 4169 13024 4185 13088
rect 4249 13024 4265 13088
rect 4329 13024 4345 13088
rect 4409 13024 4417 13088
rect 4097 13023 4417 13024
rect 10403 13088 10723 13089
rect 10403 13024 10411 13088
rect 10475 13024 10491 13088
rect 10555 13024 10571 13088
rect 10635 13024 10651 13088
rect 10715 13024 10723 13088
rect 10403 13023 10723 13024
rect 16710 13088 17030 13089
rect 16710 13024 16718 13088
rect 16782 13024 16798 13088
rect 16862 13024 16878 13088
rect 16942 13024 16958 13088
rect 17022 13024 17030 13088
rect 16710 13023 17030 13024
rect 17125 13018 17191 13021
rect 18439 13018 18919 13048
rect 17125 13016 18919 13018
rect 17125 12960 17130 13016
rect 17186 12960 18919 13016
rect 17125 12958 18919 12960
rect 17125 12955 17191 12958
rect 18439 12928 18919 12958
rect 7250 12544 7570 12545
rect 0 12472 480 12504
rect 7250 12480 7258 12544
rect 7322 12480 7338 12544
rect 7402 12480 7418 12544
rect 7482 12480 7498 12544
rect 7562 12480 7570 12544
rect 7250 12479 7570 12480
rect 13557 12544 13877 12545
rect 13557 12480 13565 12544
rect 13629 12480 13645 12544
rect 13709 12480 13725 12544
rect 13789 12480 13805 12544
rect 13869 12480 13877 12544
rect 13557 12479 13877 12480
rect 0 12416 110 12472
rect 166 12416 480 12472
rect 0 12384 480 12416
rect 4097 12000 4417 12001
rect 4097 11936 4105 12000
rect 4169 11936 4185 12000
rect 4249 11936 4265 12000
rect 4329 11936 4345 12000
rect 4409 11936 4417 12000
rect 4097 11935 4417 11936
rect 10403 12000 10723 12001
rect 10403 11936 10411 12000
rect 10475 11936 10491 12000
rect 10555 11936 10571 12000
rect 10635 11936 10651 12000
rect 10715 11936 10723 12000
rect 10403 11935 10723 11936
rect 16710 12000 17030 12001
rect 16710 11936 16718 12000
rect 16782 11936 16798 12000
rect 16862 11936 16878 12000
rect 16942 11936 16958 12000
rect 17022 11936 17030 12000
rect 16710 11935 17030 11936
rect 18439 11704 18919 11824
rect 4613 11658 4679 11661
rect 15193 11658 15259 11661
rect 4613 11656 15259 11658
rect 4613 11600 4618 11656
rect 4674 11600 15198 11656
rect 15254 11600 15259 11656
rect 4613 11598 15259 11600
rect 4613 11595 4679 11598
rect 15193 11595 15259 11598
rect 7250 11456 7570 11457
rect 7250 11392 7258 11456
rect 7322 11392 7338 11456
rect 7402 11392 7418 11456
rect 7482 11392 7498 11456
rect 7562 11392 7570 11456
rect 7250 11391 7570 11392
rect 13557 11456 13877 11457
rect 13557 11392 13565 11456
rect 13629 11392 13645 11456
rect 13709 11392 13725 11456
rect 13789 11392 13805 11456
rect 13869 11392 13877 11456
rect 13557 11391 13877 11392
rect 14825 11250 14891 11253
rect 18462 11250 18522 11704
rect 14825 11248 18522 11250
rect 14825 11192 14830 11248
rect 14886 11192 18522 11248
rect 14825 11190 18522 11192
rect 14825 11187 14891 11190
rect 4097 10912 4417 10913
rect 4097 10848 4105 10912
rect 4169 10848 4185 10912
rect 4249 10848 4265 10912
rect 4329 10848 4345 10912
rect 4409 10848 4417 10912
rect 4097 10847 4417 10848
rect 10403 10912 10723 10913
rect 10403 10848 10411 10912
rect 10475 10848 10491 10912
rect 10555 10848 10571 10912
rect 10635 10848 10651 10912
rect 10715 10848 10723 10912
rect 10403 10847 10723 10848
rect 16710 10912 17030 10913
rect 16710 10848 16718 10912
rect 16782 10848 16798 10912
rect 16862 10848 16878 10912
rect 16942 10848 16958 10912
rect 17022 10848 17030 10912
rect 16710 10847 17030 10848
rect 0 10480 480 10600
rect 62 10026 122 10480
rect 7250 10368 7570 10369
rect 7250 10304 7258 10368
rect 7322 10304 7338 10368
rect 7402 10304 7418 10368
rect 7482 10304 7498 10368
rect 7562 10304 7570 10368
rect 7250 10303 7570 10304
rect 13557 10368 13877 10369
rect 13557 10304 13565 10368
rect 13629 10304 13645 10368
rect 13709 10304 13725 10368
rect 13789 10304 13805 10368
rect 13869 10304 13877 10368
rect 18439 10344 18919 10464
rect 13557 10303 13877 10304
rect 1301 10026 1367 10029
rect 62 10024 1367 10026
rect 62 9968 1306 10024
rect 1362 9968 1367 10024
rect 62 9966 1367 9968
rect 1301 9963 1367 9966
rect 14457 10026 14523 10029
rect 18462 10026 18522 10344
rect 14457 10024 18522 10026
rect 14457 9968 14462 10024
rect 14518 9968 18522 10024
rect 14457 9966 18522 9968
rect 14457 9963 14523 9966
rect 4097 9824 4417 9825
rect 4097 9760 4105 9824
rect 4169 9760 4185 9824
rect 4249 9760 4265 9824
rect 4329 9760 4345 9824
rect 4409 9760 4417 9824
rect 4097 9759 4417 9760
rect 10403 9824 10723 9825
rect 10403 9760 10411 9824
rect 10475 9760 10491 9824
rect 10555 9760 10571 9824
rect 10635 9760 10651 9824
rect 10715 9760 10723 9824
rect 10403 9759 10723 9760
rect 16710 9824 17030 9825
rect 16710 9760 16718 9824
rect 16782 9760 16798 9824
rect 16862 9760 16878 9824
rect 16942 9760 16958 9824
rect 17022 9760 17030 9824
rect 16710 9759 17030 9760
rect 7250 9280 7570 9281
rect 7250 9216 7258 9280
rect 7322 9216 7338 9280
rect 7402 9216 7418 9280
rect 7482 9216 7498 9280
rect 7562 9216 7570 9280
rect 7250 9215 7570 9216
rect 13557 9280 13877 9281
rect 13557 9216 13565 9280
rect 13629 9216 13645 9280
rect 13709 9216 13725 9280
rect 13789 9216 13805 9280
rect 13869 9216 13877 9280
rect 13557 9215 13877 9216
rect 18439 9213 18919 9240
rect 18413 9210 18919 9213
rect 18332 9208 18919 9210
rect 18332 9152 18418 9208
rect 18474 9152 18919 9208
rect 18332 9150 18919 9152
rect 18413 9147 18919 9150
rect 18439 9120 18919 9147
rect 4097 8736 4417 8737
rect 0 8576 480 8696
rect 4097 8672 4105 8736
rect 4169 8672 4185 8736
rect 4249 8672 4265 8736
rect 4329 8672 4345 8736
rect 4409 8672 4417 8736
rect 4097 8671 4417 8672
rect 10403 8736 10723 8737
rect 10403 8672 10411 8736
rect 10475 8672 10491 8736
rect 10555 8672 10571 8736
rect 10635 8672 10651 8736
rect 10715 8672 10723 8736
rect 10403 8671 10723 8672
rect 16710 8736 17030 8737
rect 16710 8672 16718 8736
rect 16782 8672 16798 8736
rect 16862 8672 16878 8736
rect 16942 8672 16958 8736
rect 17022 8672 17030 8736
rect 16710 8671 17030 8672
rect 62 8122 122 8576
rect 7250 8192 7570 8193
rect 7250 8128 7258 8192
rect 7322 8128 7338 8192
rect 7402 8128 7418 8192
rect 7482 8128 7498 8192
rect 7562 8128 7570 8192
rect 7250 8127 7570 8128
rect 13557 8192 13877 8193
rect 13557 8128 13565 8192
rect 13629 8128 13645 8192
rect 13709 8128 13725 8192
rect 13789 8128 13805 8192
rect 13869 8128 13877 8192
rect 13557 8127 13877 8128
rect 4429 8122 4495 8125
rect 62 8120 4495 8122
rect 62 8064 4434 8120
rect 4490 8064 4495 8120
rect 62 8062 4495 8064
rect 4429 8059 4495 8062
rect 15469 7986 15535 7989
rect 18439 7986 18919 8016
rect 15469 7984 18919 7986
rect 15469 7928 15474 7984
rect 15530 7928 18919 7984
rect 15469 7926 18919 7928
rect 15469 7923 15535 7926
rect 18439 7896 18919 7926
rect 4097 7648 4417 7649
rect 4097 7584 4105 7648
rect 4169 7584 4185 7648
rect 4249 7584 4265 7648
rect 4329 7584 4345 7648
rect 4409 7584 4417 7648
rect 4097 7583 4417 7584
rect 10403 7648 10723 7649
rect 10403 7584 10411 7648
rect 10475 7584 10491 7648
rect 10555 7584 10571 7648
rect 10635 7584 10651 7648
rect 10715 7584 10723 7648
rect 10403 7583 10723 7584
rect 16710 7648 17030 7649
rect 16710 7584 16718 7648
rect 16782 7584 16798 7648
rect 16862 7584 16878 7648
rect 16942 7584 16958 7648
rect 17022 7584 17030 7648
rect 16710 7583 17030 7584
rect 7250 7104 7570 7105
rect 7250 7040 7258 7104
rect 7322 7040 7338 7104
rect 7402 7040 7418 7104
rect 7482 7040 7498 7104
rect 7562 7040 7570 7104
rect 7250 7039 7570 7040
rect 13557 7104 13877 7105
rect 13557 7040 13565 7104
rect 13629 7040 13645 7104
rect 13709 7040 13725 7104
rect 13789 7040 13805 7104
rect 13869 7040 13877 7104
rect 13557 7039 13877 7040
rect 0 6760 480 6792
rect 0 6704 110 6760
rect 166 6704 480 6760
rect 0 6672 480 6704
rect 18439 6672 18919 6792
rect 4097 6560 4417 6561
rect 4097 6496 4105 6560
rect 4169 6496 4185 6560
rect 4249 6496 4265 6560
rect 4329 6496 4345 6560
rect 4409 6496 4417 6560
rect 4097 6495 4417 6496
rect 10403 6560 10723 6561
rect 10403 6496 10411 6560
rect 10475 6496 10491 6560
rect 10555 6496 10571 6560
rect 10635 6496 10651 6560
rect 10715 6496 10723 6560
rect 10403 6495 10723 6496
rect 16710 6560 17030 6561
rect 16710 6496 16718 6560
rect 16782 6496 16798 6560
rect 16862 6496 16878 6560
rect 16942 6496 16958 6560
rect 17022 6496 17030 6560
rect 16710 6495 17030 6496
rect 17125 6490 17191 6493
rect 18462 6490 18522 6672
rect 17125 6488 18522 6490
rect 17125 6432 17130 6488
rect 17186 6432 18522 6488
rect 17125 6430 18522 6432
rect 17125 6427 17191 6430
rect 17033 6082 17099 6085
rect 17033 6080 18522 6082
rect 17033 6024 17038 6080
rect 17094 6024 18522 6080
rect 17033 6022 18522 6024
rect 17033 6019 17099 6022
rect 7250 6016 7570 6017
rect 7250 5952 7258 6016
rect 7322 5952 7338 6016
rect 7402 5952 7418 6016
rect 7482 5952 7498 6016
rect 7562 5952 7570 6016
rect 7250 5951 7570 5952
rect 13557 6016 13877 6017
rect 13557 5952 13565 6016
rect 13629 5952 13645 6016
rect 13709 5952 13725 6016
rect 13789 5952 13805 6016
rect 13869 5952 13877 6016
rect 13557 5951 13877 5952
rect 18462 5568 18522 6022
rect 4097 5472 4417 5473
rect 4097 5408 4105 5472
rect 4169 5408 4185 5472
rect 4249 5408 4265 5472
rect 4329 5408 4345 5472
rect 4409 5408 4417 5472
rect 4097 5407 4417 5408
rect 10403 5472 10723 5473
rect 10403 5408 10411 5472
rect 10475 5408 10491 5472
rect 10555 5408 10571 5472
rect 10635 5408 10651 5472
rect 10715 5408 10723 5472
rect 10403 5407 10723 5408
rect 16710 5472 17030 5473
rect 16710 5408 16718 5472
rect 16782 5408 16798 5472
rect 16862 5408 16878 5472
rect 16942 5408 16958 5472
rect 17022 5408 17030 5472
rect 18439 5448 18919 5568
rect 16710 5407 17030 5408
rect 12341 5130 12407 5133
rect 62 5128 12407 5130
rect 62 5072 12346 5128
rect 12402 5072 12407 5128
rect 62 5070 12407 5072
rect 62 4888 122 5070
rect 12341 5067 12407 5070
rect 7250 4928 7570 4929
rect 0 4768 480 4888
rect 7250 4864 7258 4928
rect 7322 4864 7338 4928
rect 7402 4864 7418 4928
rect 7482 4864 7498 4928
rect 7562 4864 7570 4928
rect 7250 4863 7570 4864
rect 13557 4928 13877 4929
rect 13557 4864 13565 4928
rect 13629 4864 13645 4928
rect 13709 4864 13725 4928
rect 13789 4864 13805 4928
rect 13869 4864 13877 4928
rect 13557 4863 13877 4864
rect 4097 4384 4417 4385
rect 4097 4320 4105 4384
rect 4169 4320 4185 4384
rect 4249 4320 4265 4384
rect 4329 4320 4345 4384
rect 4409 4320 4417 4384
rect 4097 4319 4417 4320
rect 10403 4384 10723 4385
rect 10403 4320 10411 4384
rect 10475 4320 10491 4384
rect 10555 4320 10571 4384
rect 10635 4320 10651 4384
rect 10715 4320 10723 4384
rect 10403 4319 10723 4320
rect 16710 4384 17030 4385
rect 16710 4320 16718 4384
rect 16782 4320 16798 4384
rect 16862 4320 16878 4384
rect 16942 4320 16958 4384
rect 17022 4320 17030 4384
rect 16710 4319 17030 4320
rect 18439 4224 18919 4344
rect 54 3980 60 4044
rect 124 4042 130 4044
rect 1669 4042 1735 4045
rect 124 4040 1735 4042
rect 124 3984 1674 4040
rect 1730 3984 1735 4040
rect 124 3982 1735 3984
rect 124 3980 130 3982
rect 1669 3979 1735 3982
rect 7250 3840 7570 3841
rect 7250 3776 7258 3840
rect 7322 3776 7338 3840
rect 7402 3776 7418 3840
rect 7482 3776 7498 3840
rect 7562 3776 7570 3840
rect 7250 3775 7570 3776
rect 13557 3840 13877 3841
rect 13557 3776 13565 3840
rect 13629 3776 13645 3840
rect 13709 3776 13725 3840
rect 13789 3776 13805 3840
rect 13869 3776 13877 3840
rect 13557 3775 13877 3776
rect 4097 3296 4417 3297
rect 4097 3232 4105 3296
rect 4169 3232 4185 3296
rect 4249 3232 4265 3296
rect 4329 3232 4345 3296
rect 4409 3232 4417 3296
rect 4097 3231 4417 3232
rect 10403 3296 10723 3297
rect 10403 3232 10411 3296
rect 10475 3232 10491 3296
rect 10555 3232 10571 3296
rect 10635 3232 10651 3296
rect 10715 3232 10723 3296
rect 10403 3231 10723 3232
rect 16710 3296 17030 3297
rect 16710 3232 16718 3296
rect 16782 3232 16798 3296
rect 16862 3232 16878 3296
rect 16942 3232 16958 3296
rect 17022 3232 17030 3296
rect 16710 3231 17030 3232
rect 18439 3000 18919 3120
rect 0 2956 480 2984
rect 0 2892 60 2956
rect 124 2892 480 2956
rect 0 2864 480 2892
rect 7250 2752 7570 2753
rect 7250 2688 7258 2752
rect 7322 2688 7338 2752
rect 7402 2688 7418 2752
rect 7482 2688 7498 2752
rect 7562 2688 7570 2752
rect 7250 2687 7570 2688
rect 13557 2752 13877 2753
rect 13557 2688 13565 2752
rect 13629 2688 13645 2752
rect 13709 2688 13725 2752
rect 13789 2688 13805 2752
rect 13869 2688 13877 2752
rect 13557 2687 13877 2688
rect 4097 2208 4417 2209
rect 4097 2144 4105 2208
rect 4169 2144 4185 2208
rect 4249 2144 4265 2208
rect 4329 2144 4345 2208
rect 4409 2144 4417 2208
rect 4097 2143 4417 2144
rect 10403 2208 10723 2209
rect 10403 2144 10411 2208
rect 10475 2144 10491 2208
rect 10555 2144 10571 2208
rect 10635 2144 10651 2208
rect 10715 2144 10723 2208
rect 10403 2143 10723 2144
rect 16710 2208 17030 2209
rect 16710 2144 16718 2208
rect 16782 2144 16798 2208
rect 16862 2144 16878 2208
rect 16942 2144 16958 2208
rect 17022 2144 17030 2208
rect 16710 2143 17030 2144
rect 6729 2002 6795 2005
rect 13997 2002 14063 2005
rect 6729 2000 14063 2002
rect 6729 1944 6734 2000
rect 6790 1944 14002 2000
rect 14058 1944 14063 2000
rect 6729 1942 14063 1944
rect 6729 1939 6795 1942
rect 13997 1939 14063 1942
rect 18439 1776 18919 1896
rect 0 960 480 1080
rect 18439 552 18919 672
rect 2681 98 2747 101
rect 10409 98 10475 101
rect 2681 96 10475 98
rect 2681 40 2686 96
rect 2742 40 10414 96
rect 10470 40 10475 96
rect 2681 38 10475 40
rect 2681 35 2747 38
rect 10409 35 10475 38
<< via3 >>
rect 4105 18524 4169 18528
rect 4105 18468 4109 18524
rect 4109 18468 4165 18524
rect 4165 18468 4169 18524
rect 4105 18464 4169 18468
rect 4185 18524 4249 18528
rect 4185 18468 4189 18524
rect 4189 18468 4245 18524
rect 4245 18468 4249 18524
rect 4185 18464 4249 18468
rect 4265 18524 4329 18528
rect 4265 18468 4269 18524
rect 4269 18468 4325 18524
rect 4325 18468 4329 18524
rect 4265 18464 4329 18468
rect 4345 18524 4409 18528
rect 4345 18468 4349 18524
rect 4349 18468 4405 18524
rect 4405 18468 4409 18524
rect 4345 18464 4409 18468
rect 10411 18524 10475 18528
rect 10411 18468 10415 18524
rect 10415 18468 10471 18524
rect 10471 18468 10475 18524
rect 10411 18464 10475 18468
rect 10491 18524 10555 18528
rect 10491 18468 10495 18524
rect 10495 18468 10551 18524
rect 10551 18468 10555 18524
rect 10491 18464 10555 18468
rect 10571 18524 10635 18528
rect 10571 18468 10575 18524
rect 10575 18468 10631 18524
rect 10631 18468 10635 18524
rect 10571 18464 10635 18468
rect 10651 18524 10715 18528
rect 10651 18468 10655 18524
rect 10655 18468 10711 18524
rect 10711 18468 10715 18524
rect 10651 18464 10715 18468
rect 16718 18524 16782 18528
rect 16718 18468 16722 18524
rect 16722 18468 16778 18524
rect 16778 18468 16782 18524
rect 16718 18464 16782 18468
rect 16798 18524 16862 18528
rect 16798 18468 16802 18524
rect 16802 18468 16858 18524
rect 16858 18468 16862 18524
rect 16798 18464 16862 18468
rect 16878 18524 16942 18528
rect 16878 18468 16882 18524
rect 16882 18468 16938 18524
rect 16938 18468 16942 18524
rect 16878 18464 16942 18468
rect 16958 18524 17022 18528
rect 16958 18468 16962 18524
rect 16962 18468 17018 18524
rect 17018 18468 17022 18524
rect 16958 18464 17022 18468
rect 7258 17980 7322 17984
rect 7258 17924 7262 17980
rect 7262 17924 7318 17980
rect 7318 17924 7322 17980
rect 7258 17920 7322 17924
rect 7338 17980 7402 17984
rect 7338 17924 7342 17980
rect 7342 17924 7398 17980
rect 7398 17924 7402 17980
rect 7338 17920 7402 17924
rect 7418 17980 7482 17984
rect 7418 17924 7422 17980
rect 7422 17924 7478 17980
rect 7478 17924 7482 17980
rect 7418 17920 7482 17924
rect 7498 17980 7562 17984
rect 7498 17924 7502 17980
rect 7502 17924 7558 17980
rect 7558 17924 7562 17980
rect 7498 17920 7562 17924
rect 13565 17980 13629 17984
rect 13565 17924 13569 17980
rect 13569 17924 13625 17980
rect 13625 17924 13629 17980
rect 13565 17920 13629 17924
rect 13645 17980 13709 17984
rect 13645 17924 13649 17980
rect 13649 17924 13705 17980
rect 13705 17924 13709 17980
rect 13645 17920 13709 17924
rect 13725 17980 13789 17984
rect 13725 17924 13729 17980
rect 13729 17924 13785 17980
rect 13785 17924 13789 17980
rect 13725 17920 13789 17924
rect 13805 17980 13869 17984
rect 13805 17924 13809 17980
rect 13809 17924 13865 17980
rect 13865 17924 13869 17980
rect 13805 17920 13869 17924
rect 4105 17436 4169 17440
rect 4105 17380 4109 17436
rect 4109 17380 4165 17436
rect 4165 17380 4169 17436
rect 4105 17376 4169 17380
rect 4185 17436 4249 17440
rect 4185 17380 4189 17436
rect 4189 17380 4245 17436
rect 4245 17380 4249 17436
rect 4185 17376 4249 17380
rect 4265 17436 4329 17440
rect 4265 17380 4269 17436
rect 4269 17380 4325 17436
rect 4325 17380 4329 17436
rect 4265 17376 4329 17380
rect 4345 17436 4409 17440
rect 4345 17380 4349 17436
rect 4349 17380 4405 17436
rect 4405 17380 4409 17436
rect 4345 17376 4409 17380
rect 10411 17436 10475 17440
rect 10411 17380 10415 17436
rect 10415 17380 10471 17436
rect 10471 17380 10475 17436
rect 10411 17376 10475 17380
rect 10491 17436 10555 17440
rect 10491 17380 10495 17436
rect 10495 17380 10551 17436
rect 10551 17380 10555 17436
rect 10491 17376 10555 17380
rect 10571 17436 10635 17440
rect 10571 17380 10575 17436
rect 10575 17380 10631 17436
rect 10631 17380 10635 17436
rect 10571 17376 10635 17380
rect 10651 17436 10715 17440
rect 10651 17380 10655 17436
rect 10655 17380 10711 17436
rect 10711 17380 10715 17436
rect 10651 17376 10715 17380
rect 16718 17436 16782 17440
rect 16718 17380 16722 17436
rect 16722 17380 16778 17436
rect 16778 17380 16782 17436
rect 16718 17376 16782 17380
rect 16798 17436 16862 17440
rect 16798 17380 16802 17436
rect 16802 17380 16858 17436
rect 16858 17380 16862 17436
rect 16798 17376 16862 17380
rect 16878 17436 16942 17440
rect 16878 17380 16882 17436
rect 16882 17380 16938 17436
rect 16938 17380 16942 17436
rect 16878 17376 16942 17380
rect 16958 17436 17022 17440
rect 16958 17380 16962 17436
rect 16962 17380 17018 17436
rect 17018 17380 17022 17436
rect 16958 17376 17022 17380
rect 7258 16892 7322 16896
rect 7258 16836 7262 16892
rect 7262 16836 7318 16892
rect 7318 16836 7322 16892
rect 7258 16832 7322 16836
rect 7338 16892 7402 16896
rect 7338 16836 7342 16892
rect 7342 16836 7398 16892
rect 7398 16836 7402 16892
rect 7338 16832 7402 16836
rect 7418 16892 7482 16896
rect 7418 16836 7422 16892
rect 7422 16836 7478 16892
rect 7478 16836 7482 16892
rect 7418 16832 7482 16836
rect 7498 16892 7562 16896
rect 7498 16836 7502 16892
rect 7502 16836 7558 16892
rect 7558 16836 7562 16892
rect 7498 16832 7562 16836
rect 13565 16892 13629 16896
rect 13565 16836 13569 16892
rect 13569 16836 13625 16892
rect 13625 16836 13629 16892
rect 13565 16832 13629 16836
rect 13645 16892 13709 16896
rect 13645 16836 13649 16892
rect 13649 16836 13705 16892
rect 13705 16836 13709 16892
rect 13645 16832 13709 16836
rect 13725 16892 13789 16896
rect 13725 16836 13729 16892
rect 13729 16836 13785 16892
rect 13785 16836 13789 16892
rect 13725 16832 13789 16836
rect 13805 16892 13869 16896
rect 13805 16836 13809 16892
rect 13809 16836 13865 16892
rect 13865 16836 13869 16892
rect 13805 16832 13869 16836
rect 4105 16348 4169 16352
rect 4105 16292 4109 16348
rect 4109 16292 4165 16348
rect 4165 16292 4169 16348
rect 4105 16288 4169 16292
rect 4185 16348 4249 16352
rect 4185 16292 4189 16348
rect 4189 16292 4245 16348
rect 4245 16292 4249 16348
rect 4185 16288 4249 16292
rect 4265 16348 4329 16352
rect 4265 16292 4269 16348
rect 4269 16292 4325 16348
rect 4325 16292 4329 16348
rect 4265 16288 4329 16292
rect 4345 16348 4409 16352
rect 4345 16292 4349 16348
rect 4349 16292 4405 16348
rect 4405 16292 4409 16348
rect 4345 16288 4409 16292
rect 10411 16348 10475 16352
rect 10411 16292 10415 16348
rect 10415 16292 10471 16348
rect 10471 16292 10475 16348
rect 10411 16288 10475 16292
rect 10491 16348 10555 16352
rect 10491 16292 10495 16348
rect 10495 16292 10551 16348
rect 10551 16292 10555 16348
rect 10491 16288 10555 16292
rect 10571 16348 10635 16352
rect 10571 16292 10575 16348
rect 10575 16292 10631 16348
rect 10631 16292 10635 16348
rect 10571 16288 10635 16292
rect 10651 16348 10715 16352
rect 10651 16292 10655 16348
rect 10655 16292 10711 16348
rect 10711 16292 10715 16348
rect 10651 16288 10715 16292
rect 16718 16348 16782 16352
rect 16718 16292 16722 16348
rect 16722 16292 16778 16348
rect 16778 16292 16782 16348
rect 16718 16288 16782 16292
rect 16798 16348 16862 16352
rect 16798 16292 16802 16348
rect 16802 16292 16858 16348
rect 16858 16292 16862 16348
rect 16798 16288 16862 16292
rect 16878 16348 16942 16352
rect 16878 16292 16882 16348
rect 16882 16292 16938 16348
rect 16938 16292 16942 16348
rect 16878 16288 16942 16292
rect 16958 16348 17022 16352
rect 16958 16292 16962 16348
rect 16962 16292 17018 16348
rect 17018 16292 17022 16348
rect 16958 16288 17022 16292
rect 7258 15804 7322 15808
rect 7258 15748 7262 15804
rect 7262 15748 7318 15804
rect 7318 15748 7322 15804
rect 7258 15744 7322 15748
rect 7338 15804 7402 15808
rect 7338 15748 7342 15804
rect 7342 15748 7398 15804
rect 7398 15748 7402 15804
rect 7338 15744 7402 15748
rect 7418 15804 7482 15808
rect 7418 15748 7422 15804
rect 7422 15748 7478 15804
rect 7478 15748 7482 15804
rect 7418 15744 7482 15748
rect 7498 15804 7562 15808
rect 7498 15748 7502 15804
rect 7502 15748 7558 15804
rect 7558 15748 7562 15804
rect 7498 15744 7562 15748
rect 13565 15804 13629 15808
rect 13565 15748 13569 15804
rect 13569 15748 13625 15804
rect 13625 15748 13629 15804
rect 13565 15744 13629 15748
rect 13645 15804 13709 15808
rect 13645 15748 13649 15804
rect 13649 15748 13705 15804
rect 13705 15748 13709 15804
rect 13645 15744 13709 15748
rect 13725 15804 13789 15808
rect 13725 15748 13729 15804
rect 13729 15748 13785 15804
rect 13785 15748 13789 15804
rect 13725 15744 13789 15748
rect 13805 15804 13869 15808
rect 13805 15748 13809 15804
rect 13809 15748 13865 15804
rect 13865 15748 13869 15804
rect 13805 15744 13869 15748
rect 4105 15260 4169 15264
rect 4105 15204 4109 15260
rect 4109 15204 4165 15260
rect 4165 15204 4169 15260
rect 4105 15200 4169 15204
rect 4185 15260 4249 15264
rect 4185 15204 4189 15260
rect 4189 15204 4245 15260
rect 4245 15204 4249 15260
rect 4185 15200 4249 15204
rect 4265 15260 4329 15264
rect 4265 15204 4269 15260
rect 4269 15204 4325 15260
rect 4325 15204 4329 15260
rect 4265 15200 4329 15204
rect 4345 15260 4409 15264
rect 4345 15204 4349 15260
rect 4349 15204 4405 15260
rect 4405 15204 4409 15260
rect 4345 15200 4409 15204
rect 10411 15260 10475 15264
rect 10411 15204 10415 15260
rect 10415 15204 10471 15260
rect 10471 15204 10475 15260
rect 10411 15200 10475 15204
rect 10491 15260 10555 15264
rect 10491 15204 10495 15260
rect 10495 15204 10551 15260
rect 10551 15204 10555 15260
rect 10491 15200 10555 15204
rect 10571 15260 10635 15264
rect 10571 15204 10575 15260
rect 10575 15204 10631 15260
rect 10631 15204 10635 15260
rect 10571 15200 10635 15204
rect 10651 15260 10715 15264
rect 10651 15204 10655 15260
rect 10655 15204 10711 15260
rect 10711 15204 10715 15260
rect 10651 15200 10715 15204
rect 16718 15260 16782 15264
rect 16718 15204 16722 15260
rect 16722 15204 16778 15260
rect 16778 15204 16782 15260
rect 16718 15200 16782 15204
rect 16798 15260 16862 15264
rect 16798 15204 16802 15260
rect 16802 15204 16858 15260
rect 16858 15204 16862 15260
rect 16798 15200 16862 15204
rect 16878 15260 16942 15264
rect 16878 15204 16882 15260
rect 16882 15204 16938 15260
rect 16938 15204 16942 15260
rect 16878 15200 16942 15204
rect 16958 15260 17022 15264
rect 16958 15204 16962 15260
rect 16962 15204 17018 15260
rect 17018 15204 17022 15260
rect 16958 15200 17022 15204
rect 7258 14716 7322 14720
rect 7258 14660 7262 14716
rect 7262 14660 7318 14716
rect 7318 14660 7322 14716
rect 7258 14656 7322 14660
rect 7338 14716 7402 14720
rect 7338 14660 7342 14716
rect 7342 14660 7398 14716
rect 7398 14660 7402 14716
rect 7338 14656 7402 14660
rect 7418 14716 7482 14720
rect 7418 14660 7422 14716
rect 7422 14660 7478 14716
rect 7478 14660 7482 14716
rect 7418 14656 7482 14660
rect 7498 14716 7562 14720
rect 7498 14660 7502 14716
rect 7502 14660 7558 14716
rect 7558 14660 7562 14716
rect 7498 14656 7562 14660
rect 13565 14716 13629 14720
rect 13565 14660 13569 14716
rect 13569 14660 13625 14716
rect 13625 14660 13629 14716
rect 13565 14656 13629 14660
rect 13645 14716 13709 14720
rect 13645 14660 13649 14716
rect 13649 14660 13705 14716
rect 13705 14660 13709 14716
rect 13645 14656 13709 14660
rect 13725 14716 13789 14720
rect 13725 14660 13729 14716
rect 13729 14660 13785 14716
rect 13785 14660 13789 14716
rect 13725 14656 13789 14660
rect 13805 14716 13869 14720
rect 13805 14660 13809 14716
rect 13809 14660 13865 14716
rect 13865 14660 13869 14716
rect 13805 14656 13869 14660
rect 4105 14172 4169 14176
rect 4105 14116 4109 14172
rect 4109 14116 4165 14172
rect 4165 14116 4169 14172
rect 4105 14112 4169 14116
rect 4185 14172 4249 14176
rect 4185 14116 4189 14172
rect 4189 14116 4245 14172
rect 4245 14116 4249 14172
rect 4185 14112 4249 14116
rect 4265 14172 4329 14176
rect 4265 14116 4269 14172
rect 4269 14116 4325 14172
rect 4325 14116 4329 14172
rect 4265 14112 4329 14116
rect 4345 14172 4409 14176
rect 4345 14116 4349 14172
rect 4349 14116 4405 14172
rect 4405 14116 4409 14172
rect 4345 14112 4409 14116
rect 10411 14172 10475 14176
rect 10411 14116 10415 14172
rect 10415 14116 10471 14172
rect 10471 14116 10475 14172
rect 10411 14112 10475 14116
rect 10491 14172 10555 14176
rect 10491 14116 10495 14172
rect 10495 14116 10551 14172
rect 10551 14116 10555 14172
rect 10491 14112 10555 14116
rect 10571 14172 10635 14176
rect 10571 14116 10575 14172
rect 10575 14116 10631 14172
rect 10631 14116 10635 14172
rect 10571 14112 10635 14116
rect 10651 14172 10715 14176
rect 10651 14116 10655 14172
rect 10655 14116 10711 14172
rect 10711 14116 10715 14172
rect 10651 14112 10715 14116
rect 16718 14172 16782 14176
rect 16718 14116 16722 14172
rect 16722 14116 16778 14172
rect 16778 14116 16782 14172
rect 16718 14112 16782 14116
rect 16798 14172 16862 14176
rect 16798 14116 16802 14172
rect 16802 14116 16858 14172
rect 16858 14116 16862 14172
rect 16798 14112 16862 14116
rect 16878 14172 16942 14176
rect 16878 14116 16882 14172
rect 16882 14116 16938 14172
rect 16938 14116 16942 14172
rect 16878 14112 16942 14116
rect 16958 14172 17022 14176
rect 16958 14116 16962 14172
rect 16962 14116 17018 14172
rect 17018 14116 17022 14172
rect 16958 14112 17022 14116
rect 7258 13628 7322 13632
rect 7258 13572 7262 13628
rect 7262 13572 7318 13628
rect 7318 13572 7322 13628
rect 7258 13568 7322 13572
rect 7338 13628 7402 13632
rect 7338 13572 7342 13628
rect 7342 13572 7398 13628
rect 7398 13572 7402 13628
rect 7338 13568 7402 13572
rect 7418 13628 7482 13632
rect 7418 13572 7422 13628
rect 7422 13572 7478 13628
rect 7478 13572 7482 13628
rect 7418 13568 7482 13572
rect 7498 13628 7562 13632
rect 7498 13572 7502 13628
rect 7502 13572 7558 13628
rect 7558 13572 7562 13628
rect 7498 13568 7562 13572
rect 13565 13628 13629 13632
rect 13565 13572 13569 13628
rect 13569 13572 13625 13628
rect 13625 13572 13629 13628
rect 13565 13568 13629 13572
rect 13645 13628 13709 13632
rect 13645 13572 13649 13628
rect 13649 13572 13705 13628
rect 13705 13572 13709 13628
rect 13645 13568 13709 13572
rect 13725 13628 13789 13632
rect 13725 13572 13729 13628
rect 13729 13572 13785 13628
rect 13785 13572 13789 13628
rect 13725 13568 13789 13572
rect 13805 13628 13869 13632
rect 13805 13572 13809 13628
rect 13809 13572 13865 13628
rect 13865 13572 13869 13628
rect 13805 13568 13869 13572
rect 4105 13084 4169 13088
rect 4105 13028 4109 13084
rect 4109 13028 4165 13084
rect 4165 13028 4169 13084
rect 4105 13024 4169 13028
rect 4185 13084 4249 13088
rect 4185 13028 4189 13084
rect 4189 13028 4245 13084
rect 4245 13028 4249 13084
rect 4185 13024 4249 13028
rect 4265 13084 4329 13088
rect 4265 13028 4269 13084
rect 4269 13028 4325 13084
rect 4325 13028 4329 13084
rect 4265 13024 4329 13028
rect 4345 13084 4409 13088
rect 4345 13028 4349 13084
rect 4349 13028 4405 13084
rect 4405 13028 4409 13084
rect 4345 13024 4409 13028
rect 10411 13084 10475 13088
rect 10411 13028 10415 13084
rect 10415 13028 10471 13084
rect 10471 13028 10475 13084
rect 10411 13024 10475 13028
rect 10491 13084 10555 13088
rect 10491 13028 10495 13084
rect 10495 13028 10551 13084
rect 10551 13028 10555 13084
rect 10491 13024 10555 13028
rect 10571 13084 10635 13088
rect 10571 13028 10575 13084
rect 10575 13028 10631 13084
rect 10631 13028 10635 13084
rect 10571 13024 10635 13028
rect 10651 13084 10715 13088
rect 10651 13028 10655 13084
rect 10655 13028 10711 13084
rect 10711 13028 10715 13084
rect 10651 13024 10715 13028
rect 16718 13084 16782 13088
rect 16718 13028 16722 13084
rect 16722 13028 16778 13084
rect 16778 13028 16782 13084
rect 16718 13024 16782 13028
rect 16798 13084 16862 13088
rect 16798 13028 16802 13084
rect 16802 13028 16858 13084
rect 16858 13028 16862 13084
rect 16798 13024 16862 13028
rect 16878 13084 16942 13088
rect 16878 13028 16882 13084
rect 16882 13028 16938 13084
rect 16938 13028 16942 13084
rect 16878 13024 16942 13028
rect 16958 13084 17022 13088
rect 16958 13028 16962 13084
rect 16962 13028 17018 13084
rect 17018 13028 17022 13084
rect 16958 13024 17022 13028
rect 7258 12540 7322 12544
rect 7258 12484 7262 12540
rect 7262 12484 7318 12540
rect 7318 12484 7322 12540
rect 7258 12480 7322 12484
rect 7338 12540 7402 12544
rect 7338 12484 7342 12540
rect 7342 12484 7398 12540
rect 7398 12484 7402 12540
rect 7338 12480 7402 12484
rect 7418 12540 7482 12544
rect 7418 12484 7422 12540
rect 7422 12484 7478 12540
rect 7478 12484 7482 12540
rect 7418 12480 7482 12484
rect 7498 12540 7562 12544
rect 7498 12484 7502 12540
rect 7502 12484 7558 12540
rect 7558 12484 7562 12540
rect 7498 12480 7562 12484
rect 13565 12540 13629 12544
rect 13565 12484 13569 12540
rect 13569 12484 13625 12540
rect 13625 12484 13629 12540
rect 13565 12480 13629 12484
rect 13645 12540 13709 12544
rect 13645 12484 13649 12540
rect 13649 12484 13705 12540
rect 13705 12484 13709 12540
rect 13645 12480 13709 12484
rect 13725 12540 13789 12544
rect 13725 12484 13729 12540
rect 13729 12484 13785 12540
rect 13785 12484 13789 12540
rect 13725 12480 13789 12484
rect 13805 12540 13869 12544
rect 13805 12484 13809 12540
rect 13809 12484 13865 12540
rect 13865 12484 13869 12540
rect 13805 12480 13869 12484
rect 4105 11996 4169 12000
rect 4105 11940 4109 11996
rect 4109 11940 4165 11996
rect 4165 11940 4169 11996
rect 4105 11936 4169 11940
rect 4185 11996 4249 12000
rect 4185 11940 4189 11996
rect 4189 11940 4245 11996
rect 4245 11940 4249 11996
rect 4185 11936 4249 11940
rect 4265 11996 4329 12000
rect 4265 11940 4269 11996
rect 4269 11940 4325 11996
rect 4325 11940 4329 11996
rect 4265 11936 4329 11940
rect 4345 11996 4409 12000
rect 4345 11940 4349 11996
rect 4349 11940 4405 11996
rect 4405 11940 4409 11996
rect 4345 11936 4409 11940
rect 10411 11996 10475 12000
rect 10411 11940 10415 11996
rect 10415 11940 10471 11996
rect 10471 11940 10475 11996
rect 10411 11936 10475 11940
rect 10491 11996 10555 12000
rect 10491 11940 10495 11996
rect 10495 11940 10551 11996
rect 10551 11940 10555 11996
rect 10491 11936 10555 11940
rect 10571 11996 10635 12000
rect 10571 11940 10575 11996
rect 10575 11940 10631 11996
rect 10631 11940 10635 11996
rect 10571 11936 10635 11940
rect 10651 11996 10715 12000
rect 10651 11940 10655 11996
rect 10655 11940 10711 11996
rect 10711 11940 10715 11996
rect 10651 11936 10715 11940
rect 16718 11996 16782 12000
rect 16718 11940 16722 11996
rect 16722 11940 16778 11996
rect 16778 11940 16782 11996
rect 16718 11936 16782 11940
rect 16798 11996 16862 12000
rect 16798 11940 16802 11996
rect 16802 11940 16858 11996
rect 16858 11940 16862 11996
rect 16798 11936 16862 11940
rect 16878 11996 16942 12000
rect 16878 11940 16882 11996
rect 16882 11940 16938 11996
rect 16938 11940 16942 11996
rect 16878 11936 16942 11940
rect 16958 11996 17022 12000
rect 16958 11940 16962 11996
rect 16962 11940 17018 11996
rect 17018 11940 17022 11996
rect 16958 11936 17022 11940
rect 7258 11452 7322 11456
rect 7258 11396 7262 11452
rect 7262 11396 7318 11452
rect 7318 11396 7322 11452
rect 7258 11392 7322 11396
rect 7338 11452 7402 11456
rect 7338 11396 7342 11452
rect 7342 11396 7398 11452
rect 7398 11396 7402 11452
rect 7338 11392 7402 11396
rect 7418 11452 7482 11456
rect 7418 11396 7422 11452
rect 7422 11396 7478 11452
rect 7478 11396 7482 11452
rect 7418 11392 7482 11396
rect 7498 11452 7562 11456
rect 7498 11396 7502 11452
rect 7502 11396 7558 11452
rect 7558 11396 7562 11452
rect 7498 11392 7562 11396
rect 13565 11452 13629 11456
rect 13565 11396 13569 11452
rect 13569 11396 13625 11452
rect 13625 11396 13629 11452
rect 13565 11392 13629 11396
rect 13645 11452 13709 11456
rect 13645 11396 13649 11452
rect 13649 11396 13705 11452
rect 13705 11396 13709 11452
rect 13645 11392 13709 11396
rect 13725 11452 13789 11456
rect 13725 11396 13729 11452
rect 13729 11396 13785 11452
rect 13785 11396 13789 11452
rect 13725 11392 13789 11396
rect 13805 11452 13869 11456
rect 13805 11396 13809 11452
rect 13809 11396 13865 11452
rect 13865 11396 13869 11452
rect 13805 11392 13869 11396
rect 4105 10908 4169 10912
rect 4105 10852 4109 10908
rect 4109 10852 4165 10908
rect 4165 10852 4169 10908
rect 4105 10848 4169 10852
rect 4185 10908 4249 10912
rect 4185 10852 4189 10908
rect 4189 10852 4245 10908
rect 4245 10852 4249 10908
rect 4185 10848 4249 10852
rect 4265 10908 4329 10912
rect 4265 10852 4269 10908
rect 4269 10852 4325 10908
rect 4325 10852 4329 10908
rect 4265 10848 4329 10852
rect 4345 10908 4409 10912
rect 4345 10852 4349 10908
rect 4349 10852 4405 10908
rect 4405 10852 4409 10908
rect 4345 10848 4409 10852
rect 10411 10908 10475 10912
rect 10411 10852 10415 10908
rect 10415 10852 10471 10908
rect 10471 10852 10475 10908
rect 10411 10848 10475 10852
rect 10491 10908 10555 10912
rect 10491 10852 10495 10908
rect 10495 10852 10551 10908
rect 10551 10852 10555 10908
rect 10491 10848 10555 10852
rect 10571 10908 10635 10912
rect 10571 10852 10575 10908
rect 10575 10852 10631 10908
rect 10631 10852 10635 10908
rect 10571 10848 10635 10852
rect 10651 10908 10715 10912
rect 10651 10852 10655 10908
rect 10655 10852 10711 10908
rect 10711 10852 10715 10908
rect 10651 10848 10715 10852
rect 16718 10908 16782 10912
rect 16718 10852 16722 10908
rect 16722 10852 16778 10908
rect 16778 10852 16782 10908
rect 16718 10848 16782 10852
rect 16798 10908 16862 10912
rect 16798 10852 16802 10908
rect 16802 10852 16858 10908
rect 16858 10852 16862 10908
rect 16798 10848 16862 10852
rect 16878 10908 16942 10912
rect 16878 10852 16882 10908
rect 16882 10852 16938 10908
rect 16938 10852 16942 10908
rect 16878 10848 16942 10852
rect 16958 10908 17022 10912
rect 16958 10852 16962 10908
rect 16962 10852 17018 10908
rect 17018 10852 17022 10908
rect 16958 10848 17022 10852
rect 7258 10364 7322 10368
rect 7258 10308 7262 10364
rect 7262 10308 7318 10364
rect 7318 10308 7322 10364
rect 7258 10304 7322 10308
rect 7338 10364 7402 10368
rect 7338 10308 7342 10364
rect 7342 10308 7398 10364
rect 7398 10308 7402 10364
rect 7338 10304 7402 10308
rect 7418 10364 7482 10368
rect 7418 10308 7422 10364
rect 7422 10308 7478 10364
rect 7478 10308 7482 10364
rect 7418 10304 7482 10308
rect 7498 10364 7562 10368
rect 7498 10308 7502 10364
rect 7502 10308 7558 10364
rect 7558 10308 7562 10364
rect 7498 10304 7562 10308
rect 13565 10364 13629 10368
rect 13565 10308 13569 10364
rect 13569 10308 13625 10364
rect 13625 10308 13629 10364
rect 13565 10304 13629 10308
rect 13645 10364 13709 10368
rect 13645 10308 13649 10364
rect 13649 10308 13705 10364
rect 13705 10308 13709 10364
rect 13645 10304 13709 10308
rect 13725 10364 13789 10368
rect 13725 10308 13729 10364
rect 13729 10308 13785 10364
rect 13785 10308 13789 10364
rect 13725 10304 13789 10308
rect 13805 10364 13869 10368
rect 13805 10308 13809 10364
rect 13809 10308 13865 10364
rect 13865 10308 13869 10364
rect 13805 10304 13869 10308
rect 4105 9820 4169 9824
rect 4105 9764 4109 9820
rect 4109 9764 4165 9820
rect 4165 9764 4169 9820
rect 4105 9760 4169 9764
rect 4185 9820 4249 9824
rect 4185 9764 4189 9820
rect 4189 9764 4245 9820
rect 4245 9764 4249 9820
rect 4185 9760 4249 9764
rect 4265 9820 4329 9824
rect 4265 9764 4269 9820
rect 4269 9764 4325 9820
rect 4325 9764 4329 9820
rect 4265 9760 4329 9764
rect 4345 9820 4409 9824
rect 4345 9764 4349 9820
rect 4349 9764 4405 9820
rect 4405 9764 4409 9820
rect 4345 9760 4409 9764
rect 10411 9820 10475 9824
rect 10411 9764 10415 9820
rect 10415 9764 10471 9820
rect 10471 9764 10475 9820
rect 10411 9760 10475 9764
rect 10491 9820 10555 9824
rect 10491 9764 10495 9820
rect 10495 9764 10551 9820
rect 10551 9764 10555 9820
rect 10491 9760 10555 9764
rect 10571 9820 10635 9824
rect 10571 9764 10575 9820
rect 10575 9764 10631 9820
rect 10631 9764 10635 9820
rect 10571 9760 10635 9764
rect 10651 9820 10715 9824
rect 10651 9764 10655 9820
rect 10655 9764 10711 9820
rect 10711 9764 10715 9820
rect 10651 9760 10715 9764
rect 16718 9820 16782 9824
rect 16718 9764 16722 9820
rect 16722 9764 16778 9820
rect 16778 9764 16782 9820
rect 16718 9760 16782 9764
rect 16798 9820 16862 9824
rect 16798 9764 16802 9820
rect 16802 9764 16858 9820
rect 16858 9764 16862 9820
rect 16798 9760 16862 9764
rect 16878 9820 16942 9824
rect 16878 9764 16882 9820
rect 16882 9764 16938 9820
rect 16938 9764 16942 9820
rect 16878 9760 16942 9764
rect 16958 9820 17022 9824
rect 16958 9764 16962 9820
rect 16962 9764 17018 9820
rect 17018 9764 17022 9820
rect 16958 9760 17022 9764
rect 7258 9276 7322 9280
rect 7258 9220 7262 9276
rect 7262 9220 7318 9276
rect 7318 9220 7322 9276
rect 7258 9216 7322 9220
rect 7338 9276 7402 9280
rect 7338 9220 7342 9276
rect 7342 9220 7398 9276
rect 7398 9220 7402 9276
rect 7338 9216 7402 9220
rect 7418 9276 7482 9280
rect 7418 9220 7422 9276
rect 7422 9220 7478 9276
rect 7478 9220 7482 9276
rect 7418 9216 7482 9220
rect 7498 9276 7562 9280
rect 7498 9220 7502 9276
rect 7502 9220 7558 9276
rect 7558 9220 7562 9276
rect 7498 9216 7562 9220
rect 13565 9276 13629 9280
rect 13565 9220 13569 9276
rect 13569 9220 13625 9276
rect 13625 9220 13629 9276
rect 13565 9216 13629 9220
rect 13645 9276 13709 9280
rect 13645 9220 13649 9276
rect 13649 9220 13705 9276
rect 13705 9220 13709 9276
rect 13645 9216 13709 9220
rect 13725 9276 13789 9280
rect 13725 9220 13729 9276
rect 13729 9220 13785 9276
rect 13785 9220 13789 9276
rect 13725 9216 13789 9220
rect 13805 9276 13869 9280
rect 13805 9220 13809 9276
rect 13809 9220 13865 9276
rect 13865 9220 13869 9276
rect 13805 9216 13869 9220
rect 4105 8732 4169 8736
rect 4105 8676 4109 8732
rect 4109 8676 4165 8732
rect 4165 8676 4169 8732
rect 4105 8672 4169 8676
rect 4185 8732 4249 8736
rect 4185 8676 4189 8732
rect 4189 8676 4245 8732
rect 4245 8676 4249 8732
rect 4185 8672 4249 8676
rect 4265 8732 4329 8736
rect 4265 8676 4269 8732
rect 4269 8676 4325 8732
rect 4325 8676 4329 8732
rect 4265 8672 4329 8676
rect 4345 8732 4409 8736
rect 4345 8676 4349 8732
rect 4349 8676 4405 8732
rect 4405 8676 4409 8732
rect 4345 8672 4409 8676
rect 10411 8732 10475 8736
rect 10411 8676 10415 8732
rect 10415 8676 10471 8732
rect 10471 8676 10475 8732
rect 10411 8672 10475 8676
rect 10491 8732 10555 8736
rect 10491 8676 10495 8732
rect 10495 8676 10551 8732
rect 10551 8676 10555 8732
rect 10491 8672 10555 8676
rect 10571 8732 10635 8736
rect 10571 8676 10575 8732
rect 10575 8676 10631 8732
rect 10631 8676 10635 8732
rect 10571 8672 10635 8676
rect 10651 8732 10715 8736
rect 10651 8676 10655 8732
rect 10655 8676 10711 8732
rect 10711 8676 10715 8732
rect 10651 8672 10715 8676
rect 16718 8732 16782 8736
rect 16718 8676 16722 8732
rect 16722 8676 16778 8732
rect 16778 8676 16782 8732
rect 16718 8672 16782 8676
rect 16798 8732 16862 8736
rect 16798 8676 16802 8732
rect 16802 8676 16858 8732
rect 16858 8676 16862 8732
rect 16798 8672 16862 8676
rect 16878 8732 16942 8736
rect 16878 8676 16882 8732
rect 16882 8676 16938 8732
rect 16938 8676 16942 8732
rect 16878 8672 16942 8676
rect 16958 8732 17022 8736
rect 16958 8676 16962 8732
rect 16962 8676 17018 8732
rect 17018 8676 17022 8732
rect 16958 8672 17022 8676
rect 7258 8188 7322 8192
rect 7258 8132 7262 8188
rect 7262 8132 7318 8188
rect 7318 8132 7322 8188
rect 7258 8128 7322 8132
rect 7338 8188 7402 8192
rect 7338 8132 7342 8188
rect 7342 8132 7398 8188
rect 7398 8132 7402 8188
rect 7338 8128 7402 8132
rect 7418 8188 7482 8192
rect 7418 8132 7422 8188
rect 7422 8132 7478 8188
rect 7478 8132 7482 8188
rect 7418 8128 7482 8132
rect 7498 8188 7562 8192
rect 7498 8132 7502 8188
rect 7502 8132 7558 8188
rect 7558 8132 7562 8188
rect 7498 8128 7562 8132
rect 13565 8188 13629 8192
rect 13565 8132 13569 8188
rect 13569 8132 13625 8188
rect 13625 8132 13629 8188
rect 13565 8128 13629 8132
rect 13645 8188 13709 8192
rect 13645 8132 13649 8188
rect 13649 8132 13705 8188
rect 13705 8132 13709 8188
rect 13645 8128 13709 8132
rect 13725 8188 13789 8192
rect 13725 8132 13729 8188
rect 13729 8132 13785 8188
rect 13785 8132 13789 8188
rect 13725 8128 13789 8132
rect 13805 8188 13869 8192
rect 13805 8132 13809 8188
rect 13809 8132 13865 8188
rect 13865 8132 13869 8188
rect 13805 8128 13869 8132
rect 4105 7644 4169 7648
rect 4105 7588 4109 7644
rect 4109 7588 4165 7644
rect 4165 7588 4169 7644
rect 4105 7584 4169 7588
rect 4185 7644 4249 7648
rect 4185 7588 4189 7644
rect 4189 7588 4245 7644
rect 4245 7588 4249 7644
rect 4185 7584 4249 7588
rect 4265 7644 4329 7648
rect 4265 7588 4269 7644
rect 4269 7588 4325 7644
rect 4325 7588 4329 7644
rect 4265 7584 4329 7588
rect 4345 7644 4409 7648
rect 4345 7588 4349 7644
rect 4349 7588 4405 7644
rect 4405 7588 4409 7644
rect 4345 7584 4409 7588
rect 10411 7644 10475 7648
rect 10411 7588 10415 7644
rect 10415 7588 10471 7644
rect 10471 7588 10475 7644
rect 10411 7584 10475 7588
rect 10491 7644 10555 7648
rect 10491 7588 10495 7644
rect 10495 7588 10551 7644
rect 10551 7588 10555 7644
rect 10491 7584 10555 7588
rect 10571 7644 10635 7648
rect 10571 7588 10575 7644
rect 10575 7588 10631 7644
rect 10631 7588 10635 7644
rect 10571 7584 10635 7588
rect 10651 7644 10715 7648
rect 10651 7588 10655 7644
rect 10655 7588 10711 7644
rect 10711 7588 10715 7644
rect 10651 7584 10715 7588
rect 16718 7644 16782 7648
rect 16718 7588 16722 7644
rect 16722 7588 16778 7644
rect 16778 7588 16782 7644
rect 16718 7584 16782 7588
rect 16798 7644 16862 7648
rect 16798 7588 16802 7644
rect 16802 7588 16858 7644
rect 16858 7588 16862 7644
rect 16798 7584 16862 7588
rect 16878 7644 16942 7648
rect 16878 7588 16882 7644
rect 16882 7588 16938 7644
rect 16938 7588 16942 7644
rect 16878 7584 16942 7588
rect 16958 7644 17022 7648
rect 16958 7588 16962 7644
rect 16962 7588 17018 7644
rect 17018 7588 17022 7644
rect 16958 7584 17022 7588
rect 7258 7100 7322 7104
rect 7258 7044 7262 7100
rect 7262 7044 7318 7100
rect 7318 7044 7322 7100
rect 7258 7040 7322 7044
rect 7338 7100 7402 7104
rect 7338 7044 7342 7100
rect 7342 7044 7398 7100
rect 7398 7044 7402 7100
rect 7338 7040 7402 7044
rect 7418 7100 7482 7104
rect 7418 7044 7422 7100
rect 7422 7044 7478 7100
rect 7478 7044 7482 7100
rect 7418 7040 7482 7044
rect 7498 7100 7562 7104
rect 7498 7044 7502 7100
rect 7502 7044 7558 7100
rect 7558 7044 7562 7100
rect 7498 7040 7562 7044
rect 13565 7100 13629 7104
rect 13565 7044 13569 7100
rect 13569 7044 13625 7100
rect 13625 7044 13629 7100
rect 13565 7040 13629 7044
rect 13645 7100 13709 7104
rect 13645 7044 13649 7100
rect 13649 7044 13705 7100
rect 13705 7044 13709 7100
rect 13645 7040 13709 7044
rect 13725 7100 13789 7104
rect 13725 7044 13729 7100
rect 13729 7044 13785 7100
rect 13785 7044 13789 7100
rect 13725 7040 13789 7044
rect 13805 7100 13869 7104
rect 13805 7044 13809 7100
rect 13809 7044 13865 7100
rect 13865 7044 13869 7100
rect 13805 7040 13869 7044
rect 4105 6556 4169 6560
rect 4105 6500 4109 6556
rect 4109 6500 4165 6556
rect 4165 6500 4169 6556
rect 4105 6496 4169 6500
rect 4185 6556 4249 6560
rect 4185 6500 4189 6556
rect 4189 6500 4245 6556
rect 4245 6500 4249 6556
rect 4185 6496 4249 6500
rect 4265 6556 4329 6560
rect 4265 6500 4269 6556
rect 4269 6500 4325 6556
rect 4325 6500 4329 6556
rect 4265 6496 4329 6500
rect 4345 6556 4409 6560
rect 4345 6500 4349 6556
rect 4349 6500 4405 6556
rect 4405 6500 4409 6556
rect 4345 6496 4409 6500
rect 10411 6556 10475 6560
rect 10411 6500 10415 6556
rect 10415 6500 10471 6556
rect 10471 6500 10475 6556
rect 10411 6496 10475 6500
rect 10491 6556 10555 6560
rect 10491 6500 10495 6556
rect 10495 6500 10551 6556
rect 10551 6500 10555 6556
rect 10491 6496 10555 6500
rect 10571 6556 10635 6560
rect 10571 6500 10575 6556
rect 10575 6500 10631 6556
rect 10631 6500 10635 6556
rect 10571 6496 10635 6500
rect 10651 6556 10715 6560
rect 10651 6500 10655 6556
rect 10655 6500 10711 6556
rect 10711 6500 10715 6556
rect 10651 6496 10715 6500
rect 16718 6556 16782 6560
rect 16718 6500 16722 6556
rect 16722 6500 16778 6556
rect 16778 6500 16782 6556
rect 16718 6496 16782 6500
rect 16798 6556 16862 6560
rect 16798 6500 16802 6556
rect 16802 6500 16858 6556
rect 16858 6500 16862 6556
rect 16798 6496 16862 6500
rect 16878 6556 16942 6560
rect 16878 6500 16882 6556
rect 16882 6500 16938 6556
rect 16938 6500 16942 6556
rect 16878 6496 16942 6500
rect 16958 6556 17022 6560
rect 16958 6500 16962 6556
rect 16962 6500 17018 6556
rect 17018 6500 17022 6556
rect 16958 6496 17022 6500
rect 7258 6012 7322 6016
rect 7258 5956 7262 6012
rect 7262 5956 7318 6012
rect 7318 5956 7322 6012
rect 7258 5952 7322 5956
rect 7338 6012 7402 6016
rect 7338 5956 7342 6012
rect 7342 5956 7398 6012
rect 7398 5956 7402 6012
rect 7338 5952 7402 5956
rect 7418 6012 7482 6016
rect 7418 5956 7422 6012
rect 7422 5956 7478 6012
rect 7478 5956 7482 6012
rect 7418 5952 7482 5956
rect 7498 6012 7562 6016
rect 7498 5956 7502 6012
rect 7502 5956 7558 6012
rect 7558 5956 7562 6012
rect 7498 5952 7562 5956
rect 13565 6012 13629 6016
rect 13565 5956 13569 6012
rect 13569 5956 13625 6012
rect 13625 5956 13629 6012
rect 13565 5952 13629 5956
rect 13645 6012 13709 6016
rect 13645 5956 13649 6012
rect 13649 5956 13705 6012
rect 13705 5956 13709 6012
rect 13645 5952 13709 5956
rect 13725 6012 13789 6016
rect 13725 5956 13729 6012
rect 13729 5956 13785 6012
rect 13785 5956 13789 6012
rect 13725 5952 13789 5956
rect 13805 6012 13869 6016
rect 13805 5956 13809 6012
rect 13809 5956 13865 6012
rect 13865 5956 13869 6012
rect 13805 5952 13869 5956
rect 4105 5468 4169 5472
rect 4105 5412 4109 5468
rect 4109 5412 4165 5468
rect 4165 5412 4169 5468
rect 4105 5408 4169 5412
rect 4185 5468 4249 5472
rect 4185 5412 4189 5468
rect 4189 5412 4245 5468
rect 4245 5412 4249 5468
rect 4185 5408 4249 5412
rect 4265 5468 4329 5472
rect 4265 5412 4269 5468
rect 4269 5412 4325 5468
rect 4325 5412 4329 5468
rect 4265 5408 4329 5412
rect 4345 5468 4409 5472
rect 4345 5412 4349 5468
rect 4349 5412 4405 5468
rect 4405 5412 4409 5468
rect 4345 5408 4409 5412
rect 10411 5468 10475 5472
rect 10411 5412 10415 5468
rect 10415 5412 10471 5468
rect 10471 5412 10475 5468
rect 10411 5408 10475 5412
rect 10491 5468 10555 5472
rect 10491 5412 10495 5468
rect 10495 5412 10551 5468
rect 10551 5412 10555 5468
rect 10491 5408 10555 5412
rect 10571 5468 10635 5472
rect 10571 5412 10575 5468
rect 10575 5412 10631 5468
rect 10631 5412 10635 5468
rect 10571 5408 10635 5412
rect 10651 5468 10715 5472
rect 10651 5412 10655 5468
rect 10655 5412 10711 5468
rect 10711 5412 10715 5468
rect 10651 5408 10715 5412
rect 16718 5468 16782 5472
rect 16718 5412 16722 5468
rect 16722 5412 16778 5468
rect 16778 5412 16782 5468
rect 16718 5408 16782 5412
rect 16798 5468 16862 5472
rect 16798 5412 16802 5468
rect 16802 5412 16858 5468
rect 16858 5412 16862 5468
rect 16798 5408 16862 5412
rect 16878 5468 16942 5472
rect 16878 5412 16882 5468
rect 16882 5412 16938 5468
rect 16938 5412 16942 5468
rect 16878 5408 16942 5412
rect 16958 5468 17022 5472
rect 16958 5412 16962 5468
rect 16962 5412 17018 5468
rect 17018 5412 17022 5468
rect 16958 5408 17022 5412
rect 7258 4924 7322 4928
rect 7258 4868 7262 4924
rect 7262 4868 7318 4924
rect 7318 4868 7322 4924
rect 7258 4864 7322 4868
rect 7338 4924 7402 4928
rect 7338 4868 7342 4924
rect 7342 4868 7398 4924
rect 7398 4868 7402 4924
rect 7338 4864 7402 4868
rect 7418 4924 7482 4928
rect 7418 4868 7422 4924
rect 7422 4868 7478 4924
rect 7478 4868 7482 4924
rect 7418 4864 7482 4868
rect 7498 4924 7562 4928
rect 7498 4868 7502 4924
rect 7502 4868 7558 4924
rect 7558 4868 7562 4924
rect 7498 4864 7562 4868
rect 13565 4924 13629 4928
rect 13565 4868 13569 4924
rect 13569 4868 13625 4924
rect 13625 4868 13629 4924
rect 13565 4864 13629 4868
rect 13645 4924 13709 4928
rect 13645 4868 13649 4924
rect 13649 4868 13705 4924
rect 13705 4868 13709 4924
rect 13645 4864 13709 4868
rect 13725 4924 13789 4928
rect 13725 4868 13729 4924
rect 13729 4868 13785 4924
rect 13785 4868 13789 4924
rect 13725 4864 13789 4868
rect 13805 4924 13869 4928
rect 13805 4868 13809 4924
rect 13809 4868 13865 4924
rect 13865 4868 13869 4924
rect 13805 4864 13869 4868
rect 4105 4380 4169 4384
rect 4105 4324 4109 4380
rect 4109 4324 4165 4380
rect 4165 4324 4169 4380
rect 4105 4320 4169 4324
rect 4185 4380 4249 4384
rect 4185 4324 4189 4380
rect 4189 4324 4245 4380
rect 4245 4324 4249 4380
rect 4185 4320 4249 4324
rect 4265 4380 4329 4384
rect 4265 4324 4269 4380
rect 4269 4324 4325 4380
rect 4325 4324 4329 4380
rect 4265 4320 4329 4324
rect 4345 4380 4409 4384
rect 4345 4324 4349 4380
rect 4349 4324 4405 4380
rect 4405 4324 4409 4380
rect 4345 4320 4409 4324
rect 10411 4380 10475 4384
rect 10411 4324 10415 4380
rect 10415 4324 10471 4380
rect 10471 4324 10475 4380
rect 10411 4320 10475 4324
rect 10491 4380 10555 4384
rect 10491 4324 10495 4380
rect 10495 4324 10551 4380
rect 10551 4324 10555 4380
rect 10491 4320 10555 4324
rect 10571 4380 10635 4384
rect 10571 4324 10575 4380
rect 10575 4324 10631 4380
rect 10631 4324 10635 4380
rect 10571 4320 10635 4324
rect 10651 4380 10715 4384
rect 10651 4324 10655 4380
rect 10655 4324 10711 4380
rect 10711 4324 10715 4380
rect 10651 4320 10715 4324
rect 16718 4380 16782 4384
rect 16718 4324 16722 4380
rect 16722 4324 16778 4380
rect 16778 4324 16782 4380
rect 16718 4320 16782 4324
rect 16798 4380 16862 4384
rect 16798 4324 16802 4380
rect 16802 4324 16858 4380
rect 16858 4324 16862 4380
rect 16798 4320 16862 4324
rect 16878 4380 16942 4384
rect 16878 4324 16882 4380
rect 16882 4324 16938 4380
rect 16938 4324 16942 4380
rect 16878 4320 16942 4324
rect 16958 4380 17022 4384
rect 16958 4324 16962 4380
rect 16962 4324 17018 4380
rect 17018 4324 17022 4380
rect 16958 4320 17022 4324
rect 60 3980 124 4044
rect 7258 3836 7322 3840
rect 7258 3780 7262 3836
rect 7262 3780 7318 3836
rect 7318 3780 7322 3836
rect 7258 3776 7322 3780
rect 7338 3836 7402 3840
rect 7338 3780 7342 3836
rect 7342 3780 7398 3836
rect 7398 3780 7402 3836
rect 7338 3776 7402 3780
rect 7418 3836 7482 3840
rect 7418 3780 7422 3836
rect 7422 3780 7478 3836
rect 7478 3780 7482 3836
rect 7418 3776 7482 3780
rect 7498 3836 7562 3840
rect 7498 3780 7502 3836
rect 7502 3780 7558 3836
rect 7558 3780 7562 3836
rect 7498 3776 7562 3780
rect 13565 3836 13629 3840
rect 13565 3780 13569 3836
rect 13569 3780 13625 3836
rect 13625 3780 13629 3836
rect 13565 3776 13629 3780
rect 13645 3836 13709 3840
rect 13645 3780 13649 3836
rect 13649 3780 13705 3836
rect 13705 3780 13709 3836
rect 13645 3776 13709 3780
rect 13725 3836 13789 3840
rect 13725 3780 13729 3836
rect 13729 3780 13785 3836
rect 13785 3780 13789 3836
rect 13725 3776 13789 3780
rect 13805 3836 13869 3840
rect 13805 3780 13809 3836
rect 13809 3780 13865 3836
rect 13865 3780 13869 3836
rect 13805 3776 13869 3780
rect 4105 3292 4169 3296
rect 4105 3236 4109 3292
rect 4109 3236 4165 3292
rect 4165 3236 4169 3292
rect 4105 3232 4169 3236
rect 4185 3292 4249 3296
rect 4185 3236 4189 3292
rect 4189 3236 4245 3292
rect 4245 3236 4249 3292
rect 4185 3232 4249 3236
rect 4265 3292 4329 3296
rect 4265 3236 4269 3292
rect 4269 3236 4325 3292
rect 4325 3236 4329 3292
rect 4265 3232 4329 3236
rect 4345 3292 4409 3296
rect 4345 3236 4349 3292
rect 4349 3236 4405 3292
rect 4405 3236 4409 3292
rect 4345 3232 4409 3236
rect 10411 3292 10475 3296
rect 10411 3236 10415 3292
rect 10415 3236 10471 3292
rect 10471 3236 10475 3292
rect 10411 3232 10475 3236
rect 10491 3292 10555 3296
rect 10491 3236 10495 3292
rect 10495 3236 10551 3292
rect 10551 3236 10555 3292
rect 10491 3232 10555 3236
rect 10571 3292 10635 3296
rect 10571 3236 10575 3292
rect 10575 3236 10631 3292
rect 10631 3236 10635 3292
rect 10571 3232 10635 3236
rect 10651 3292 10715 3296
rect 10651 3236 10655 3292
rect 10655 3236 10711 3292
rect 10711 3236 10715 3292
rect 10651 3232 10715 3236
rect 16718 3292 16782 3296
rect 16718 3236 16722 3292
rect 16722 3236 16778 3292
rect 16778 3236 16782 3292
rect 16718 3232 16782 3236
rect 16798 3292 16862 3296
rect 16798 3236 16802 3292
rect 16802 3236 16858 3292
rect 16858 3236 16862 3292
rect 16798 3232 16862 3236
rect 16878 3292 16942 3296
rect 16878 3236 16882 3292
rect 16882 3236 16938 3292
rect 16938 3236 16942 3292
rect 16878 3232 16942 3236
rect 16958 3292 17022 3296
rect 16958 3236 16962 3292
rect 16962 3236 17018 3292
rect 17018 3236 17022 3292
rect 16958 3232 17022 3236
rect 60 2892 124 2956
rect 7258 2748 7322 2752
rect 7258 2692 7262 2748
rect 7262 2692 7318 2748
rect 7318 2692 7322 2748
rect 7258 2688 7322 2692
rect 7338 2748 7402 2752
rect 7338 2692 7342 2748
rect 7342 2692 7398 2748
rect 7398 2692 7402 2748
rect 7338 2688 7402 2692
rect 7418 2748 7482 2752
rect 7418 2692 7422 2748
rect 7422 2692 7478 2748
rect 7478 2692 7482 2748
rect 7418 2688 7482 2692
rect 7498 2748 7562 2752
rect 7498 2692 7502 2748
rect 7502 2692 7558 2748
rect 7558 2692 7562 2748
rect 7498 2688 7562 2692
rect 13565 2748 13629 2752
rect 13565 2692 13569 2748
rect 13569 2692 13625 2748
rect 13625 2692 13629 2748
rect 13565 2688 13629 2692
rect 13645 2748 13709 2752
rect 13645 2692 13649 2748
rect 13649 2692 13705 2748
rect 13705 2692 13709 2748
rect 13645 2688 13709 2692
rect 13725 2748 13789 2752
rect 13725 2692 13729 2748
rect 13729 2692 13785 2748
rect 13785 2692 13789 2748
rect 13725 2688 13789 2692
rect 13805 2748 13869 2752
rect 13805 2692 13809 2748
rect 13809 2692 13865 2748
rect 13865 2692 13869 2748
rect 13805 2688 13869 2692
rect 4105 2204 4169 2208
rect 4105 2148 4109 2204
rect 4109 2148 4165 2204
rect 4165 2148 4169 2204
rect 4105 2144 4169 2148
rect 4185 2204 4249 2208
rect 4185 2148 4189 2204
rect 4189 2148 4245 2204
rect 4245 2148 4249 2204
rect 4185 2144 4249 2148
rect 4265 2204 4329 2208
rect 4265 2148 4269 2204
rect 4269 2148 4325 2204
rect 4325 2148 4329 2204
rect 4265 2144 4329 2148
rect 4345 2204 4409 2208
rect 4345 2148 4349 2204
rect 4349 2148 4405 2204
rect 4405 2148 4409 2204
rect 4345 2144 4409 2148
rect 10411 2204 10475 2208
rect 10411 2148 10415 2204
rect 10415 2148 10471 2204
rect 10471 2148 10475 2204
rect 10411 2144 10475 2148
rect 10491 2204 10555 2208
rect 10491 2148 10495 2204
rect 10495 2148 10551 2204
rect 10551 2148 10555 2204
rect 10491 2144 10555 2148
rect 10571 2204 10635 2208
rect 10571 2148 10575 2204
rect 10575 2148 10631 2204
rect 10631 2148 10635 2204
rect 10571 2144 10635 2148
rect 10651 2204 10715 2208
rect 10651 2148 10655 2204
rect 10655 2148 10711 2204
rect 10711 2148 10715 2204
rect 10651 2144 10715 2148
rect 16718 2204 16782 2208
rect 16718 2148 16722 2204
rect 16722 2148 16778 2204
rect 16778 2148 16782 2204
rect 16718 2144 16782 2148
rect 16798 2204 16862 2208
rect 16798 2148 16802 2204
rect 16802 2148 16858 2204
rect 16858 2148 16862 2204
rect 16798 2144 16862 2148
rect 16878 2204 16942 2208
rect 16878 2148 16882 2204
rect 16882 2148 16938 2204
rect 16938 2148 16942 2204
rect 16878 2144 16942 2148
rect 16958 2204 17022 2208
rect 16958 2148 16962 2204
rect 16962 2148 17018 2204
rect 17018 2148 17022 2204
rect 16958 2144 17022 2148
<< metal4 >>
rect 4097 18528 4417 18544
rect 4097 18464 4105 18528
rect 4169 18464 4185 18528
rect 4249 18464 4265 18528
rect 4329 18464 4345 18528
rect 4409 18464 4417 18528
rect 4097 17440 4417 18464
rect 4097 17376 4105 17440
rect 4169 17376 4185 17440
rect 4249 17376 4265 17440
rect 4329 17376 4345 17440
rect 4409 17376 4417 17440
rect 4097 16352 4417 17376
rect 4097 16288 4105 16352
rect 4169 16288 4185 16352
rect 4249 16288 4265 16352
rect 4329 16288 4345 16352
rect 4409 16288 4417 16352
rect 4097 15264 4417 16288
rect 4097 15200 4105 15264
rect 4169 15200 4185 15264
rect 4249 15200 4265 15264
rect 4329 15200 4345 15264
rect 4409 15200 4417 15264
rect 4097 14176 4417 15200
rect 4097 14112 4105 14176
rect 4169 14112 4185 14176
rect 4249 14112 4265 14176
rect 4329 14112 4345 14176
rect 4409 14112 4417 14176
rect 4097 13088 4417 14112
rect 4097 13024 4105 13088
rect 4169 13024 4185 13088
rect 4249 13024 4265 13088
rect 4329 13024 4345 13088
rect 4409 13024 4417 13088
rect 4097 12000 4417 13024
rect 4097 11936 4105 12000
rect 4169 11936 4185 12000
rect 4249 11936 4265 12000
rect 4329 11936 4345 12000
rect 4409 11936 4417 12000
rect 4097 10912 4417 11936
rect 4097 10848 4105 10912
rect 4169 10848 4185 10912
rect 4249 10848 4265 10912
rect 4329 10848 4345 10912
rect 4409 10848 4417 10912
rect 4097 9824 4417 10848
rect 4097 9760 4105 9824
rect 4169 9760 4185 9824
rect 4249 9760 4265 9824
rect 4329 9760 4345 9824
rect 4409 9760 4417 9824
rect 4097 8736 4417 9760
rect 4097 8672 4105 8736
rect 4169 8672 4185 8736
rect 4249 8672 4265 8736
rect 4329 8672 4345 8736
rect 4409 8672 4417 8736
rect 4097 7648 4417 8672
rect 4097 7584 4105 7648
rect 4169 7584 4185 7648
rect 4249 7584 4265 7648
rect 4329 7584 4345 7648
rect 4409 7584 4417 7648
rect 4097 6560 4417 7584
rect 4097 6496 4105 6560
rect 4169 6496 4185 6560
rect 4249 6496 4265 6560
rect 4329 6496 4345 6560
rect 4409 6496 4417 6560
rect 4097 5472 4417 6496
rect 4097 5408 4105 5472
rect 4169 5408 4185 5472
rect 4249 5408 4265 5472
rect 4329 5408 4345 5472
rect 4409 5408 4417 5472
rect 4097 4384 4417 5408
rect 4097 4320 4105 4384
rect 4169 4320 4185 4384
rect 4249 4320 4265 4384
rect 4329 4320 4345 4384
rect 4409 4320 4417 4384
rect 59 4044 125 4045
rect 59 3980 60 4044
rect 124 3980 125 4044
rect 59 3979 125 3980
rect 62 2957 122 3979
rect 4097 3296 4417 4320
rect 4097 3232 4105 3296
rect 4169 3232 4185 3296
rect 4249 3232 4265 3296
rect 4329 3232 4345 3296
rect 4409 3232 4417 3296
rect 59 2956 125 2957
rect 59 2892 60 2956
rect 124 2892 125 2956
rect 59 2891 125 2892
rect 4097 2208 4417 3232
rect 4097 2144 4105 2208
rect 4169 2144 4185 2208
rect 4249 2144 4265 2208
rect 4329 2144 4345 2208
rect 4409 2144 4417 2208
rect 4097 2128 4417 2144
rect 7250 17984 7570 18544
rect 7250 17920 7258 17984
rect 7322 17920 7338 17984
rect 7402 17920 7418 17984
rect 7482 17920 7498 17984
rect 7562 17920 7570 17984
rect 7250 16896 7570 17920
rect 7250 16832 7258 16896
rect 7322 16832 7338 16896
rect 7402 16832 7418 16896
rect 7482 16832 7498 16896
rect 7562 16832 7570 16896
rect 7250 15808 7570 16832
rect 7250 15744 7258 15808
rect 7322 15744 7338 15808
rect 7402 15744 7418 15808
rect 7482 15744 7498 15808
rect 7562 15744 7570 15808
rect 7250 14720 7570 15744
rect 7250 14656 7258 14720
rect 7322 14656 7338 14720
rect 7402 14656 7418 14720
rect 7482 14656 7498 14720
rect 7562 14656 7570 14720
rect 7250 13632 7570 14656
rect 7250 13568 7258 13632
rect 7322 13568 7338 13632
rect 7402 13568 7418 13632
rect 7482 13568 7498 13632
rect 7562 13568 7570 13632
rect 7250 12544 7570 13568
rect 7250 12480 7258 12544
rect 7322 12480 7338 12544
rect 7402 12480 7418 12544
rect 7482 12480 7498 12544
rect 7562 12480 7570 12544
rect 7250 11456 7570 12480
rect 7250 11392 7258 11456
rect 7322 11392 7338 11456
rect 7402 11392 7418 11456
rect 7482 11392 7498 11456
rect 7562 11392 7570 11456
rect 7250 10368 7570 11392
rect 7250 10304 7258 10368
rect 7322 10304 7338 10368
rect 7402 10304 7418 10368
rect 7482 10304 7498 10368
rect 7562 10304 7570 10368
rect 7250 9280 7570 10304
rect 7250 9216 7258 9280
rect 7322 9216 7338 9280
rect 7402 9216 7418 9280
rect 7482 9216 7498 9280
rect 7562 9216 7570 9280
rect 7250 8192 7570 9216
rect 7250 8128 7258 8192
rect 7322 8128 7338 8192
rect 7402 8128 7418 8192
rect 7482 8128 7498 8192
rect 7562 8128 7570 8192
rect 7250 7104 7570 8128
rect 7250 7040 7258 7104
rect 7322 7040 7338 7104
rect 7402 7040 7418 7104
rect 7482 7040 7498 7104
rect 7562 7040 7570 7104
rect 7250 6016 7570 7040
rect 7250 5952 7258 6016
rect 7322 5952 7338 6016
rect 7402 5952 7418 6016
rect 7482 5952 7498 6016
rect 7562 5952 7570 6016
rect 7250 4928 7570 5952
rect 7250 4864 7258 4928
rect 7322 4864 7338 4928
rect 7402 4864 7418 4928
rect 7482 4864 7498 4928
rect 7562 4864 7570 4928
rect 7250 3840 7570 4864
rect 7250 3776 7258 3840
rect 7322 3776 7338 3840
rect 7402 3776 7418 3840
rect 7482 3776 7498 3840
rect 7562 3776 7570 3840
rect 7250 2752 7570 3776
rect 7250 2688 7258 2752
rect 7322 2688 7338 2752
rect 7402 2688 7418 2752
rect 7482 2688 7498 2752
rect 7562 2688 7570 2752
rect 7250 2128 7570 2688
rect 10403 18528 10723 18544
rect 10403 18464 10411 18528
rect 10475 18464 10491 18528
rect 10555 18464 10571 18528
rect 10635 18464 10651 18528
rect 10715 18464 10723 18528
rect 10403 17440 10723 18464
rect 10403 17376 10411 17440
rect 10475 17376 10491 17440
rect 10555 17376 10571 17440
rect 10635 17376 10651 17440
rect 10715 17376 10723 17440
rect 10403 16352 10723 17376
rect 10403 16288 10411 16352
rect 10475 16288 10491 16352
rect 10555 16288 10571 16352
rect 10635 16288 10651 16352
rect 10715 16288 10723 16352
rect 10403 15264 10723 16288
rect 10403 15200 10411 15264
rect 10475 15200 10491 15264
rect 10555 15200 10571 15264
rect 10635 15200 10651 15264
rect 10715 15200 10723 15264
rect 10403 14176 10723 15200
rect 10403 14112 10411 14176
rect 10475 14112 10491 14176
rect 10555 14112 10571 14176
rect 10635 14112 10651 14176
rect 10715 14112 10723 14176
rect 10403 13088 10723 14112
rect 10403 13024 10411 13088
rect 10475 13024 10491 13088
rect 10555 13024 10571 13088
rect 10635 13024 10651 13088
rect 10715 13024 10723 13088
rect 10403 12000 10723 13024
rect 10403 11936 10411 12000
rect 10475 11936 10491 12000
rect 10555 11936 10571 12000
rect 10635 11936 10651 12000
rect 10715 11936 10723 12000
rect 10403 10912 10723 11936
rect 10403 10848 10411 10912
rect 10475 10848 10491 10912
rect 10555 10848 10571 10912
rect 10635 10848 10651 10912
rect 10715 10848 10723 10912
rect 10403 9824 10723 10848
rect 10403 9760 10411 9824
rect 10475 9760 10491 9824
rect 10555 9760 10571 9824
rect 10635 9760 10651 9824
rect 10715 9760 10723 9824
rect 10403 8736 10723 9760
rect 10403 8672 10411 8736
rect 10475 8672 10491 8736
rect 10555 8672 10571 8736
rect 10635 8672 10651 8736
rect 10715 8672 10723 8736
rect 10403 7648 10723 8672
rect 10403 7584 10411 7648
rect 10475 7584 10491 7648
rect 10555 7584 10571 7648
rect 10635 7584 10651 7648
rect 10715 7584 10723 7648
rect 10403 6560 10723 7584
rect 10403 6496 10411 6560
rect 10475 6496 10491 6560
rect 10555 6496 10571 6560
rect 10635 6496 10651 6560
rect 10715 6496 10723 6560
rect 10403 5472 10723 6496
rect 10403 5408 10411 5472
rect 10475 5408 10491 5472
rect 10555 5408 10571 5472
rect 10635 5408 10651 5472
rect 10715 5408 10723 5472
rect 10403 4384 10723 5408
rect 10403 4320 10411 4384
rect 10475 4320 10491 4384
rect 10555 4320 10571 4384
rect 10635 4320 10651 4384
rect 10715 4320 10723 4384
rect 10403 3296 10723 4320
rect 10403 3232 10411 3296
rect 10475 3232 10491 3296
rect 10555 3232 10571 3296
rect 10635 3232 10651 3296
rect 10715 3232 10723 3296
rect 10403 2208 10723 3232
rect 10403 2144 10411 2208
rect 10475 2144 10491 2208
rect 10555 2144 10571 2208
rect 10635 2144 10651 2208
rect 10715 2144 10723 2208
rect 10403 2128 10723 2144
rect 13557 17984 13877 18544
rect 13557 17920 13565 17984
rect 13629 17920 13645 17984
rect 13709 17920 13725 17984
rect 13789 17920 13805 17984
rect 13869 17920 13877 17984
rect 13557 16896 13877 17920
rect 13557 16832 13565 16896
rect 13629 16832 13645 16896
rect 13709 16832 13725 16896
rect 13789 16832 13805 16896
rect 13869 16832 13877 16896
rect 13557 15808 13877 16832
rect 13557 15744 13565 15808
rect 13629 15744 13645 15808
rect 13709 15744 13725 15808
rect 13789 15744 13805 15808
rect 13869 15744 13877 15808
rect 13557 14720 13877 15744
rect 13557 14656 13565 14720
rect 13629 14656 13645 14720
rect 13709 14656 13725 14720
rect 13789 14656 13805 14720
rect 13869 14656 13877 14720
rect 13557 13632 13877 14656
rect 13557 13568 13565 13632
rect 13629 13568 13645 13632
rect 13709 13568 13725 13632
rect 13789 13568 13805 13632
rect 13869 13568 13877 13632
rect 13557 12544 13877 13568
rect 13557 12480 13565 12544
rect 13629 12480 13645 12544
rect 13709 12480 13725 12544
rect 13789 12480 13805 12544
rect 13869 12480 13877 12544
rect 13557 11456 13877 12480
rect 13557 11392 13565 11456
rect 13629 11392 13645 11456
rect 13709 11392 13725 11456
rect 13789 11392 13805 11456
rect 13869 11392 13877 11456
rect 13557 10368 13877 11392
rect 13557 10304 13565 10368
rect 13629 10304 13645 10368
rect 13709 10304 13725 10368
rect 13789 10304 13805 10368
rect 13869 10304 13877 10368
rect 13557 9280 13877 10304
rect 13557 9216 13565 9280
rect 13629 9216 13645 9280
rect 13709 9216 13725 9280
rect 13789 9216 13805 9280
rect 13869 9216 13877 9280
rect 13557 8192 13877 9216
rect 13557 8128 13565 8192
rect 13629 8128 13645 8192
rect 13709 8128 13725 8192
rect 13789 8128 13805 8192
rect 13869 8128 13877 8192
rect 13557 7104 13877 8128
rect 13557 7040 13565 7104
rect 13629 7040 13645 7104
rect 13709 7040 13725 7104
rect 13789 7040 13805 7104
rect 13869 7040 13877 7104
rect 13557 6016 13877 7040
rect 13557 5952 13565 6016
rect 13629 5952 13645 6016
rect 13709 5952 13725 6016
rect 13789 5952 13805 6016
rect 13869 5952 13877 6016
rect 13557 4928 13877 5952
rect 13557 4864 13565 4928
rect 13629 4864 13645 4928
rect 13709 4864 13725 4928
rect 13789 4864 13805 4928
rect 13869 4864 13877 4928
rect 13557 3840 13877 4864
rect 13557 3776 13565 3840
rect 13629 3776 13645 3840
rect 13709 3776 13725 3840
rect 13789 3776 13805 3840
rect 13869 3776 13877 3840
rect 13557 2752 13877 3776
rect 13557 2688 13565 2752
rect 13629 2688 13645 2752
rect 13709 2688 13725 2752
rect 13789 2688 13805 2752
rect 13869 2688 13877 2752
rect 13557 2128 13877 2688
rect 16710 18528 17030 18544
rect 16710 18464 16718 18528
rect 16782 18464 16798 18528
rect 16862 18464 16878 18528
rect 16942 18464 16958 18528
rect 17022 18464 17030 18528
rect 16710 17440 17030 18464
rect 16710 17376 16718 17440
rect 16782 17376 16798 17440
rect 16862 17376 16878 17440
rect 16942 17376 16958 17440
rect 17022 17376 17030 17440
rect 16710 16352 17030 17376
rect 16710 16288 16718 16352
rect 16782 16288 16798 16352
rect 16862 16288 16878 16352
rect 16942 16288 16958 16352
rect 17022 16288 17030 16352
rect 16710 15264 17030 16288
rect 16710 15200 16718 15264
rect 16782 15200 16798 15264
rect 16862 15200 16878 15264
rect 16942 15200 16958 15264
rect 17022 15200 17030 15264
rect 16710 14176 17030 15200
rect 16710 14112 16718 14176
rect 16782 14112 16798 14176
rect 16862 14112 16878 14176
rect 16942 14112 16958 14176
rect 17022 14112 17030 14176
rect 16710 13088 17030 14112
rect 16710 13024 16718 13088
rect 16782 13024 16798 13088
rect 16862 13024 16878 13088
rect 16942 13024 16958 13088
rect 17022 13024 17030 13088
rect 16710 12000 17030 13024
rect 16710 11936 16718 12000
rect 16782 11936 16798 12000
rect 16862 11936 16878 12000
rect 16942 11936 16958 12000
rect 17022 11936 17030 12000
rect 16710 10912 17030 11936
rect 16710 10848 16718 10912
rect 16782 10848 16798 10912
rect 16862 10848 16878 10912
rect 16942 10848 16958 10912
rect 17022 10848 17030 10912
rect 16710 9824 17030 10848
rect 16710 9760 16718 9824
rect 16782 9760 16798 9824
rect 16862 9760 16878 9824
rect 16942 9760 16958 9824
rect 17022 9760 17030 9824
rect 16710 8736 17030 9760
rect 16710 8672 16718 8736
rect 16782 8672 16798 8736
rect 16862 8672 16878 8736
rect 16942 8672 16958 8736
rect 17022 8672 17030 8736
rect 16710 7648 17030 8672
rect 16710 7584 16718 7648
rect 16782 7584 16798 7648
rect 16862 7584 16878 7648
rect 16942 7584 16958 7648
rect 17022 7584 17030 7648
rect 16710 6560 17030 7584
rect 16710 6496 16718 6560
rect 16782 6496 16798 6560
rect 16862 6496 16878 6560
rect 16942 6496 16958 6560
rect 17022 6496 17030 6560
rect 16710 5472 17030 6496
rect 16710 5408 16718 5472
rect 16782 5408 16798 5472
rect 16862 5408 16878 5472
rect 16942 5408 16958 5472
rect 17022 5408 17030 5472
rect 16710 4384 17030 5408
rect 16710 4320 16718 4384
rect 16782 4320 16798 4384
rect 16862 4320 16878 4384
rect 16942 4320 16958 4384
rect 17022 4320 17030 4384
rect 16710 3296 17030 4320
rect 16710 3232 16718 3296
rect 16782 3232 16798 3296
rect 16862 3232 16878 3296
rect 16942 3232 16958 3296
rect 17022 3232 17030 3296
rect 16710 2208 17030 3232
rect 16710 2144 16718 2208
rect 16782 2144 16798 2208
rect 16862 2144 16878 2208
rect 16942 2144 16958 2208
rect 17022 2144 17030 2208
rect 16710 2128 17030 2144
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_12 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_9
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_11 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_7
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_conb_1  _18_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _44_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_16
timestamp 1586364061
transform 1 0 2576 0 1 2720
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_60 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_33
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_37
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_41 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_49
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_44
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_48
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 590 592
use scs8hd_fill_1  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_76 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_88
timestamp 1586364061
transform 1 0 9200 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_6  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_92
timestamp 1586364061
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_104
timestamp 1586364061
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_108
timestamp 1586364061
transform 1 0 11040 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12880 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 13800 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_132
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_140
timestamp 1586364061
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_157
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 17756 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 17756 0 1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 774 592
use scs8hd_decap_8  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_9
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6164 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_2  FILLER_2_53
timestamp 1586364061
transform 1 0 5980 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_8  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_12  FILLER_2_123
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_163
timestamp 1586364061
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 17756 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_6
timestamp 1586364061
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_10
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_22
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_49
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_67
timestamp 1586364061
transform 1 0 7268 0 1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_79
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_87
timestamp 1586364061
transform 1 0 9108 0 1 3808
box -38 -48 130 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 10304 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_91
timestamp 1586364061
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_148
timestamp 1586364061
transform 1 0 14720 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_164
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 17756 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_99
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_4_110
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_124
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 17756 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_177
timestamp 1586364061
transform 1 0 17388 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_94
timestamp 1586364061
transform 1 0 9752 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_102
timestamp 1586364061
transform 1 0 10488 0 1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_144
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_152
timestamp 1586364061
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 17756 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_170
timestamp 1586364061
transform 1 0 16744 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_55
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_66
timestamp 1586364061
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_70
timestamp 1586364061
transform 1 0 7544 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_111
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 774 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_119
timestamp 1586364061
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_128
timestamp 1586364061
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_139
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_132
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_139
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_143
timestamp 1586364061
transform 1 0 14260 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_10.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_144
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_161
timestamp 1586364061
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_165
timestamp 1586364061
transform 1 0 16284 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 17756 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 17756 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_175
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_7_169
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_76
timestamp 1586364061
transform 1 0 8096 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_10.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_12  FILLER_8_128
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_10.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_6  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 17756 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_177
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 590 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_89
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_101
timestamp 1586364061
transform 1 0 10396 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13892 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_142
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_157
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 17756 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_170
timestamp 1586364061
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_174
timestamp 1586364061
transform 1 0 17112 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_4  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_39
timestamp 1586364061
transform 1 0 4692 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_10_51
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_55
timestamp 1586364061
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_65
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_77
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_6  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 866 592
use scs8hd_fill_1  FILLER_10_160
timestamp 1586364061
transform 1 0 15824 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 17756 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_98
timestamp 1586364061
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 14812 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_152
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 17756 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_177
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 130 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 1564 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_8
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_20
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_28
timestamp 1586364061
transform 1 0 3680 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_12  FILLER_12_65
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_77
timestamp 1586364061
transform 1 0 8188 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_12_89
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 17756 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_169
timestamp 1586364061
transform 1 0 16652 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_177
timestamp 1586364061
transform 1 0 17388 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_6
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_10
timestamp 1586364061
transform 1 0 2024 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_16
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_30
timestamp 1586364061
transform 1 0 3864 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_6  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_60
timestamp 1586364061
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_65
timestamp 1586364061
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_69
timestamp 1586364061
transform 1 0 7452 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_81
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_93
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 130 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 16284 0 1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 17756 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 17756 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_169
timestamp 1586364061
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_173
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_177
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_176
timestamp 1586364061
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_35
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _19_
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use scs8hd_decap_6  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 17756 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_15_170
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_83
timestamp 1586364061
transform 1 0 8740 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_91
timestamp 1586364061
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 11424
box -38 -48 866 592
use scs8hd_fill_1  FILLER_16_160
timestamp 1586364061
transform 1 0 15824 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 17756 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_6
timestamp 1586364061
transform 1 0 1656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_10
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_14
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 17756 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_177
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_14
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_26
timestamp 1586364061
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_30
timestamp 1586364061
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_6
timestamp 1586364061
transform 1 0 1656 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_14.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_8
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_21
timestamp 1586364061
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_18
timestamp 1586364061
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_34
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_30
timestamp 1586364061
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_35
timestamp 1586364061
transform 1 0 4324 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_59
timestamp 1586364061
transform 1 0 6532 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_71
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_83
timestamp 1586364061
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 130 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_163
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 17756 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 17756 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_173
timestamp 1586364061
transform 1 0 17020 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_177
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_20_175
timestamp 1586364061
transform 1 0 17204 0 -1 13600
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1656 0 1 13600
box -38 -48 866 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 5336 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_49
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 774 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 774 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_90
timestamp 1586364061
transform 1 0 9384 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_95
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_107
timestamp 1586364061
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_119
timestamp 1586364061
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 774 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 16284 0 1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_158
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_163
timestamp 1586364061
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 17756 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_169
timestamp 1586364061
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_173
timestamp 1586364061
transform 1 0 17020 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_177
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_22
timestamp 1586364061
transform 1 0 3128 0 -1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 5704 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_42
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 7912 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_66
timestamp 1586364061
transform 1 0 7176 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_77
timestamp 1586364061
transform 1 0 8188 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_22_89
timestamp 1586364061
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_96
timestamp 1586364061
transform 1 0 9936 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_120
timestamp 1586364061
transform 1 0 12144 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_132
timestamp 1586364061
transform 1 0 13248 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_6  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 14688
box -38 -48 866 592
use scs8hd_fill_1  FILLER_22_160
timestamp 1586364061
transform 1 0 15824 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 17756 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_22_170
timestamp 1586364061
transform 1 0 16744 0 -1 14688
box -38 -48 774 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_13
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_18
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_22
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_14.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3496 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_29
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_33
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_45
timestamp 1586364061
transform 1 0 5244 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_52
timestamp 1586364061
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_56
timestamp 1586364061
transform 1 0 6256 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_60
timestamp 1586364061
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_65
timestamp 1586364061
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_69
timestamp 1586364061
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 13892 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_12.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_142
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 590 592
use scs8hd_fill_2  FILLER_23_153
timestamp 1586364061
transform 1 0 15180 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_157
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 17756 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_170
timestamp 1586364061
transform 1 0 16744 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_8  FILLER_24_20
timestamp 1586364061
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_28
timestamp 1586364061
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 4968 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_40
timestamp 1586364061
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5980 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_1  FILLER_24_74
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_84
timestamp 1586364061
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_97
timestamp 1586364061
transform 1 0 10028 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_109
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_121
timestamp 1586364061
transform 1 0 12236 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_133
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_165
timestamp 1586364061
transform 1 0 16284 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 17756 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_177
timestamp 1586364061
transform 1 0 17388 0 -1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_7
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_19
timestamp 1586364061
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_23
timestamp 1586364061
transform 1 0 3220 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_29
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_42
timestamp 1586364061
transform 1 0 4968 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_53
timestamp 1586364061
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7544 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_81
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_85
timestamp 1586364061
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_89
timestamp 1586364061
transform 1 0 9292 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_101
timestamp 1586364061
transform 1 0 10396 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_113
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_121
timestamp 1586364061
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_150
timestamp 1586364061
transform 1 0 14904 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_153
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_166
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 17756 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_6
timestamp 1586364061
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_10
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_8  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_42
timestamp 1586364061
transform 1 0 4968 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_50
timestamp 1586364061
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_41
timestamp 1586364061
transform 1 0 4876 0 1 16864
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use scs8hd_decap_3  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_73
timestamp 1586364061
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_76
timestamp 1586364061
transform 1 0 8096 0 1 16864
box -38 -48 406 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_27_80
timestamp 1586364061
transform 1 0 8464 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_27_83
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_102
timestamp 1586364061
transform 1 0 10488 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_91
timestamp 1586364061
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_95
timestamp 1586364061
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_108
timestamp 1586364061
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_112
timestamp 1586364061
transform 1 0 11408 0 1 16864
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_126
timestamp 1586364061
transform 1 0 12696 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_120
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_127
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_134
timestamp 1586364061
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_140
timestamp 1586364061
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_6  FILLER_27_144
timestamp 1586364061
transform 1 0 14352 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_153
timestamp 1586364061
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_163
timestamp 1586364061
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_157
timestamp 1586364061
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 17756 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 17756 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_175
timestamp 1586364061
transform 1 0 17204 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_27_170
timestamp 1586364061
transform 1 0 16744 0 1 16864
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_18
timestamp 1586364061
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_30
timestamp 1586364061
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_35
timestamp 1586364061
transform 1 0 4324 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 17952
box -38 -48 866 592
use scs8hd_fill_1  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_57
timestamp 1586364061
transform 1 0 6348 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_72
timestamp 1586364061
transform 1 0 7728 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_84
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_101
timestamp 1586364061
transform 1 0 10396 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_4  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_139
timestamp 1586364061
transform 1 0 13892 0 -1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_163
timestamp 1586364061
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 17756 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_175
timestamp 1586364061
transform 1 0 17204 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 406 592
use scs8hd_decap_4  FILLER_29_32
timestamp 1586364061
transform 1 0 4048 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_36
timestamp 1586364061
transform 1 0 4416 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_40
timestamp 1586364061
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_44
timestamp 1586364061
transform 1 0 5152 0 1 17952
box -38 -48 590 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_53
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_57
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_61
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_66
timestamp 1586364061
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_70
timestamp 1586364061
transform 1 0 7544 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_76
timestamp 1586364061
transform 1 0 8096 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_80
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_84
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 9660 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_92
timestamp 1586364061
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_97
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_101
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 12512 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_125
timestamp 1586364061
transform 1 0 12604 0 1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13616 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_133
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_139
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_143
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_12.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_29_156
timestamp 1586364061
transform 1 0 15456 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_164
timestamp 1586364061
transform 1 0 16192 0 1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 17756 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_12.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_168
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_172
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 960 480 1080 6 address[0]
port 0 nsew default input
rlabel metal3 s 18439 552 18919 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 18439 1776 18919 1896 6 address[2]
port 2 nsew default input
rlabel metal3 s 18439 3000 18919 3120 6 address[3]
port 3 nsew default input
rlabel metal2 s 570 20583 626 21063 6 address[4]
port 4 nsew default input
rlabel metal3 s 18439 4224 18919 4344 6 address[5]
port 5 nsew default input
rlabel metal2 s 1766 20583 1822 21063 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal2 s 3054 20583 3110 21063 6 chanx_left_in[1]
port 7 nsew default input
rlabel metal3 s 0 2864 480 2984 6 chanx_left_in[2]
port 8 nsew default input
rlabel metal3 s 18439 5448 18919 5568 6 chanx_left_in[3]
port 9 nsew default input
rlabel metal3 s 18439 6672 18919 6792 6 chanx_left_in[4]
port 10 nsew default input
rlabel metal3 s 18439 7896 18919 8016 6 chanx_left_in[5]
port 11 nsew default input
rlabel metal2 s 2410 0 2466 480 6 chanx_left_in[6]
port 12 nsew default input
rlabel metal2 s 4342 20583 4398 21063 6 chanx_left_in[7]
port 13 nsew default input
rlabel metal2 s 3422 0 3478 480 6 chanx_left_in[8]
port 14 nsew default input
rlabel metal2 s 4434 0 4490 480 6 chanx_left_out[0]
port 15 nsew default tristate
rlabel metal2 s 5446 0 5502 480 6 chanx_left_out[1]
port 16 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[2]
port 17 nsew default tristate
rlabel metal2 s 6458 0 6514 480 6 chanx_left_out[3]
port 18 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chanx_left_out[4]
port 19 nsew default tristate
rlabel metal3 s 18439 9120 18919 9240 6 chanx_left_out[5]
port 20 nsew default tristate
rlabel metal2 s 5538 20583 5594 21063 6 chanx_left_out[6]
port 21 nsew default tristate
rlabel metal2 s 8390 0 8446 480 6 chanx_left_out[7]
port 22 nsew default tristate
rlabel metal2 s 9402 0 9458 480 6 chanx_left_out[8]
port 23 nsew default tristate
rlabel metal2 s 10414 0 10470 480 6 chany_top_in[0]
port 24 nsew default input
rlabel metal2 s 6826 20583 6882 21063 6 chany_top_in[1]
port 25 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_top_in[2]
port 26 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chany_top_in[3]
port 27 nsew default input
rlabel metal2 s 8114 20583 8170 21063 6 chany_top_in[4]
port 28 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chany_top_in[5]
port 29 nsew default input
rlabel metal3 s 18439 10344 18919 10464 6 chany_top_in[6]
port 30 nsew default input
rlabel metal3 s 18439 11704 18919 11824 6 chany_top_in[7]
port 31 nsew default input
rlabel metal2 s 9402 20583 9458 21063 6 chany_top_in[8]
port 32 nsew default input
rlabel metal3 s 18439 12928 18919 13048 6 chany_top_out[0]
port 33 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chany_top_out[1]
port 34 nsew default tristate
rlabel metal3 s 0 12384 480 12504 6 chany_top_out[2]
port 35 nsew default tristate
rlabel metal2 s 10598 20583 10654 21063 6 chany_top_out[3]
port 36 nsew default tristate
rlabel metal3 s 18439 14152 18919 14272 6 chany_top_out[4]
port 37 nsew default tristate
rlabel metal2 s 12438 0 12494 480 6 chany_top_out[5]
port 38 nsew default tristate
rlabel metal3 s 18439 15376 18919 15496 6 chany_top_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chany_top_out[7]
port 40 nsew default tristate
rlabel metal2 s 13358 0 13414 480 6 chany_top_out[8]
port 41 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 data_in
port 42 nsew default input
rlabel metal2 s 478 0 534 480 6 enable
port 43 nsew default input
rlabel metal3 s 18439 17824 18919 17944 6 left_bottom_grid_pin_11_
port 44 nsew default input
rlabel metal3 s 0 16192 480 16312 6 left_bottom_grid_pin_13_
port 45 nsew default input
rlabel metal3 s 18439 19048 18919 19168 6 left_bottom_grid_pin_15_
port 46 nsew default input
rlabel metal2 s 11886 20583 11942 21063 6 left_bottom_grid_pin_1_
port 47 nsew default input
rlabel metal2 s 14370 0 14426 480 6 left_bottom_grid_pin_3_
port 48 nsew default input
rlabel metal2 s 15382 0 15438 480 6 left_bottom_grid_pin_5_
port 49 nsew default input
rlabel metal2 s 13174 20583 13230 21063 6 left_bottom_grid_pin_7_
port 50 nsew default input
rlabel metal3 s 18439 16600 18919 16720 6 left_bottom_grid_pin_9_
port 51 nsew default input
rlabel metal3 s 0 18096 480 18216 6 left_top_grid_pin_10_
port 52 nsew default input
rlabel metal2 s 14462 20583 14518 21063 6 top_left_grid_pin_13_
port 53 nsew default input
rlabel metal2 s 18234 20583 18290 21063 6 top_right_grid_pin_11_
port 54 nsew default input
rlabel metal3 s 18439 20272 18919 20392 6 top_right_grid_pin_13_
port 55 nsew default input
rlabel metal2 s 18418 0 18474 480 6 top_right_grid_pin_15_
port 56 nsew default input
rlabel metal2 s 15658 20583 15714 21063 6 top_right_grid_pin_1_
port 57 nsew default input
rlabel metal2 s 16946 20583 17002 21063 6 top_right_grid_pin_3_
port 58 nsew default input
rlabel metal3 s 0 20000 480 20120 6 top_right_grid_pin_5_
port 59 nsew default input
rlabel metal2 s 16394 0 16450 480 6 top_right_grid_pin_7_
port 60 nsew default input
rlabel metal2 s 17406 0 17462 480 6 top_right_grid_pin_9_
port 61 nsew default input
rlabel metal4 s 4097 2128 4417 18544 6 vpwr
port 62 nsew default input
rlabel metal4 s 7250 2128 7570 18544 6 vgnd
port 63 nsew default input
<< end >>
