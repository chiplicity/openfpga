VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__8_
  CLASS BLOCK ;
  FOREIGN sb_0__8_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 111.600 85.930 114.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 2.400 57.760 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 19.080 114.000 19.680 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 42.200 114.000 42.800 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 44.920 114.000 45.520 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 46.960 114.000 47.560 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 49.680 114.000 50.280 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 51.720 114.000 52.320 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 53.760 114.000 54.360 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 56.480 114.000 57.080 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 58.520 114.000 59.120 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 61.240 114.000 61.840 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 63.280 114.000 63.880 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 21.120 114.000 21.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 23.840 114.000 24.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 25.880 114.000 26.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 28.600 114.000 29.200 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 30.640 114.000 31.240 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 33.360 114.000 33.960 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 35.400 114.000 36.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 37.440 114.000 38.040 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 40.160 114.000 40.760 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 66.000 114.000 66.600 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 89.120 114.000 89.720 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 91.160 114.000 91.760 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 93.880 114.000 94.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 95.920 114.000 96.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 98.640 114.000 99.240 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 100.680 114.000 101.280 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 102.720 114.000 103.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 105.440 114.000 106.040 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 107.480 114.000 108.080 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 110.200 114.000 110.800 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 68.040 114.000 68.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 70.080 114.000 70.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 72.800 114.000 73.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 74.840 114.000 75.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 77.560 114.000 78.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 79.600 114.000 80.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 82.320 114.000 82.920 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 84.360 114.000 84.960 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 86.400 114.000 87.000 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 111.600 28.890 114.000 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 2.760 114.000 3.360 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 4.800 114.000 5.400 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 7.520 114.000 8.120 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 9.560 114.000 10.160 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 12.280 114.000 12.880 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 14.320 114.000 14.920 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 17.040 114.000 17.640 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 112.240 114.000 112.840 ;
    END
  END right_top_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 4.210 4.800 112.630 100.880 ;
      LAYER met2 ;
        RECT 1.470 111.320 28.330 112.725 ;
        RECT 29.170 111.320 85.370 112.725 ;
        RECT 86.210 111.320 112.600 112.725 ;
        RECT 1.470 2.680 112.600 111.320 ;
        RECT 2.030 0.835 3.950 2.680 ;
        RECT 4.790 0.835 6.710 2.680 ;
        RECT 7.550 0.835 9.470 2.680 ;
        RECT 10.310 0.835 12.230 2.680 ;
        RECT 13.070 0.835 14.990 2.680 ;
        RECT 15.830 0.835 17.750 2.680 ;
        RECT 18.590 0.835 20.510 2.680 ;
        RECT 21.350 0.835 23.270 2.680 ;
        RECT 24.110 0.835 26.030 2.680 ;
        RECT 26.870 0.835 28.790 2.680 ;
        RECT 29.630 0.835 31.550 2.680 ;
        RECT 32.390 0.835 34.310 2.680 ;
        RECT 35.150 0.835 37.070 2.680 ;
        RECT 37.910 0.835 39.830 2.680 ;
        RECT 40.670 0.835 42.590 2.680 ;
        RECT 43.430 0.835 45.350 2.680 ;
        RECT 46.190 0.835 48.110 2.680 ;
        RECT 48.950 0.835 50.870 2.680 ;
        RECT 51.710 0.835 53.630 2.680 ;
        RECT 54.470 0.835 56.390 2.680 ;
        RECT 57.230 0.835 59.610 2.680 ;
        RECT 60.450 0.835 62.370 2.680 ;
        RECT 63.210 0.835 65.130 2.680 ;
        RECT 65.970 0.835 67.890 2.680 ;
        RECT 68.730 0.835 70.650 2.680 ;
        RECT 71.490 0.835 73.410 2.680 ;
        RECT 74.250 0.835 76.170 2.680 ;
        RECT 77.010 0.835 78.930 2.680 ;
        RECT 79.770 0.835 81.690 2.680 ;
        RECT 82.530 0.835 84.450 2.680 ;
        RECT 85.290 0.835 87.210 2.680 ;
        RECT 88.050 0.835 89.970 2.680 ;
        RECT 90.810 0.835 92.730 2.680 ;
        RECT 93.570 0.835 95.490 2.680 ;
        RECT 96.330 0.835 98.250 2.680 ;
        RECT 99.090 0.835 101.010 2.680 ;
        RECT 101.850 0.835 103.770 2.680 ;
        RECT 104.610 0.835 106.530 2.680 ;
        RECT 107.370 0.835 109.290 2.680 ;
        RECT 110.130 0.835 112.050 2.680 ;
      LAYER met3 ;
        RECT 1.445 111.840 111.200 112.705 ;
        RECT 1.445 111.200 111.600 111.840 ;
        RECT 1.445 109.800 111.200 111.200 ;
        RECT 1.445 108.480 111.600 109.800 ;
        RECT 1.445 107.080 111.200 108.480 ;
        RECT 1.445 106.440 111.600 107.080 ;
        RECT 1.445 105.040 111.200 106.440 ;
        RECT 1.445 103.720 111.600 105.040 ;
        RECT 1.445 102.320 111.200 103.720 ;
        RECT 1.445 101.680 111.600 102.320 ;
        RECT 1.445 100.280 111.200 101.680 ;
        RECT 1.445 99.640 111.600 100.280 ;
        RECT 1.445 98.240 111.200 99.640 ;
        RECT 1.445 96.920 111.600 98.240 ;
        RECT 1.445 95.520 111.200 96.920 ;
        RECT 1.445 94.880 111.600 95.520 ;
        RECT 1.445 93.480 111.200 94.880 ;
        RECT 1.445 92.160 111.600 93.480 ;
        RECT 1.445 90.760 111.200 92.160 ;
        RECT 1.445 90.120 111.600 90.760 ;
        RECT 1.445 88.720 111.200 90.120 ;
        RECT 1.445 87.400 111.600 88.720 ;
        RECT 1.445 86.000 111.200 87.400 ;
        RECT 1.445 85.360 111.600 86.000 ;
        RECT 1.445 83.960 111.200 85.360 ;
        RECT 1.445 83.320 111.600 83.960 ;
        RECT 1.445 81.920 111.200 83.320 ;
        RECT 1.445 80.600 111.600 81.920 ;
        RECT 1.445 79.200 111.200 80.600 ;
        RECT 1.445 78.560 111.600 79.200 ;
        RECT 1.445 77.160 111.200 78.560 ;
        RECT 1.445 75.840 111.600 77.160 ;
        RECT 1.445 74.440 111.200 75.840 ;
        RECT 1.445 73.800 111.600 74.440 ;
        RECT 1.445 72.400 111.200 73.800 ;
        RECT 1.445 71.080 111.600 72.400 ;
        RECT 1.445 69.680 111.200 71.080 ;
        RECT 1.445 69.040 111.600 69.680 ;
        RECT 1.445 67.640 111.200 69.040 ;
        RECT 1.445 67.000 111.600 67.640 ;
        RECT 1.445 65.600 111.200 67.000 ;
        RECT 1.445 64.280 111.600 65.600 ;
        RECT 1.445 62.880 111.200 64.280 ;
        RECT 1.445 62.240 111.600 62.880 ;
        RECT 1.445 60.840 111.200 62.240 ;
        RECT 1.445 59.520 111.600 60.840 ;
        RECT 1.445 58.160 111.200 59.520 ;
        RECT 2.800 58.120 111.200 58.160 ;
        RECT 2.800 57.480 111.600 58.120 ;
        RECT 2.800 56.760 111.200 57.480 ;
        RECT 1.445 56.080 111.200 56.760 ;
        RECT 1.445 54.760 111.600 56.080 ;
        RECT 1.445 53.360 111.200 54.760 ;
        RECT 1.445 52.720 111.600 53.360 ;
        RECT 1.445 51.320 111.200 52.720 ;
        RECT 1.445 50.680 111.600 51.320 ;
        RECT 1.445 49.280 111.200 50.680 ;
        RECT 1.445 47.960 111.600 49.280 ;
        RECT 1.445 46.560 111.200 47.960 ;
        RECT 1.445 45.920 111.600 46.560 ;
        RECT 1.445 44.520 111.200 45.920 ;
        RECT 1.445 43.200 111.600 44.520 ;
        RECT 1.445 41.800 111.200 43.200 ;
        RECT 1.445 41.160 111.600 41.800 ;
        RECT 1.445 39.760 111.200 41.160 ;
        RECT 1.445 38.440 111.600 39.760 ;
        RECT 1.445 37.040 111.200 38.440 ;
        RECT 1.445 36.400 111.600 37.040 ;
        RECT 1.445 35.000 111.200 36.400 ;
        RECT 1.445 34.360 111.600 35.000 ;
        RECT 1.445 32.960 111.200 34.360 ;
        RECT 1.445 31.640 111.600 32.960 ;
        RECT 1.445 30.240 111.200 31.640 ;
        RECT 1.445 29.600 111.600 30.240 ;
        RECT 1.445 28.200 111.200 29.600 ;
        RECT 1.445 26.880 111.600 28.200 ;
        RECT 1.445 25.480 111.200 26.880 ;
        RECT 1.445 24.840 111.600 25.480 ;
        RECT 1.445 23.440 111.200 24.840 ;
        RECT 1.445 22.120 111.600 23.440 ;
        RECT 1.445 20.720 111.200 22.120 ;
        RECT 1.445 20.080 111.600 20.720 ;
        RECT 1.445 18.680 111.200 20.080 ;
        RECT 1.445 18.040 111.600 18.680 ;
        RECT 1.445 16.640 111.200 18.040 ;
        RECT 1.445 15.320 111.600 16.640 ;
        RECT 1.445 13.920 111.200 15.320 ;
        RECT 1.445 13.280 111.600 13.920 ;
        RECT 1.445 11.880 111.200 13.280 ;
        RECT 1.445 10.560 111.600 11.880 ;
        RECT 1.445 9.160 111.200 10.560 ;
        RECT 1.445 8.520 111.600 9.160 ;
        RECT 1.445 7.120 111.200 8.520 ;
        RECT 1.445 5.800 111.600 7.120 ;
        RECT 1.445 4.400 111.200 5.800 ;
        RECT 1.445 3.760 111.600 4.400 ;
        RECT 1.445 2.360 111.200 3.760 ;
        RECT 1.445 1.720 111.600 2.360 ;
        RECT 1.445 0.855 111.200 1.720 ;
      LAYER met4 ;
        RECT 56.200 10.640 92.120 100.880 ;
  END
END sb_0__8_
END LIBRARY

