magic
tech EFS8A
magscale 1 2
timestamp 1604336873
<< viali >>
rect 23029 25449 23063 25483
rect 24777 25449 24811 25483
rect 19441 25381 19475 25415
rect 22845 25313 22879 25347
rect 24593 25313 24627 25347
rect 19441 25245 19475 25279
rect 19533 25245 19567 25279
rect 14289 25109 14323 25143
rect 18981 25109 19015 25143
rect 19349 24905 19383 24939
rect 20637 24905 20671 24939
rect 14841 24769 14875 24803
rect 18429 24769 18463 24803
rect 25145 24769 25179 24803
rect 14565 24701 14599 24735
rect 20269 24701 20303 24735
rect 22477 24701 22511 24735
rect 24593 24701 24627 24735
rect 14013 24633 14047 24667
rect 14271 24633 14305 24667
rect 19625 24633 19659 24667
rect 19901 24633 19935 24667
rect 14749 24565 14783 24599
rect 18705 24565 18739 24599
rect 19165 24565 19199 24599
rect 19809 24565 19843 24599
rect 22385 24565 22419 24599
rect 22661 24565 22695 24599
rect 23121 24565 23155 24599
rect 24409 24565 24443 24599
rect 24777 24565 24811 24599
rect 13829 24361 13863 24395
rect 14657 24361 14691 24395
rect 15485 24361 15519 24395
rect 21097 24361 21131 24395
rect 25421 24361 25455 24395
rect 19165 24293 19199 24327
rect 11417 24225 11451 24259
rect 13645 24225 13679 24259
rect 15301 24225 15335 24259
rect 20913 24225 20947 24259
rect 23020 24225 23054 24259
rect 25237 24225 25271 24259
rect 11161 24157 11195 24191
rect 19073 24157 19107 24191
rect 19257 24157 19291 24191
rect 22753 24157 22787 24191
rect 18705 24089 18739 24123
rect 10517 24021 10551 24055
rect 10885 24021 10919 24055
rect 12541 24021 12575 24055
rect 13461 24021 13495 24055
rect 14289 24021 14323 24055
rect 19717 24021 19751 24055
rect 20085 24021 20119 24055
rect 24133 24021 24167 24055
rect 10333 23817 10367 23851
rect 16865 23817 16899 23851
rect 22017 23817 22051 23851
rect 22753 23817 22787 23851
rect 23121 23817 23155 23851
rect 24777 23817 24811 23851
rect 10885 23749 10919 23783
rect 12541 23749 12575 23783
rect 11437 23681 11471 23715
rect 13001 23681 13035 23715
rect 13093 23681 13127 23715
rect 13461 23681 13495 23715
rect 25513 23681 25547 23715
rect 12173 23613 12207 23647
rect 14197 23613 14231 23647
rect 14464 23613 14498 23647
rect 16681 23613 16715 23647
rect 18613 23613 18647 23647
rect 19257 23613 19291 23647
rect 19349 23613 19383 23647
rect 19616 23613 19650 23647
rect 21833 23613 21867 23647
rect 24593 23613 24627 23647
rect 9781 23545 9815 23579
rect 10701 23545 10735 23579
rect 11161 23545 11195 23579
rect 13001 23545 13035 23579
rect 22477 23545 22511 23579
rect 11345 23477 11379 23511
rect 11805 23477 11839 23511
rect 14013 23477 14047 23511
rect 15577 23477 15611 23511
rect 16129 23477 16163 23511
rect 17233 23477 17267 23511
rect 18337 23477 18371 23511
rect 20729 23477 20763 23511
rect 21373 23477 21407 23511
rect 25237 23477 25271 23511
rect 11621 23273 11655 23307
rect 14105 23273 14139 23307
rect 18705 23273 18739 23307
rect 21097 23273 21131 23307
rect 24777 23273 24811 23307
rect 12970 23205 13004 23239
rect 19809 23205 19843 23239
rect 19901 23205 19935 23239
rect 23029 23205 23063 23239
rect 10508 23137 10542 23171
rect 16681 23137 16715 23171
rect 16948 23137 16982 23171
rect 19625 23137 19659 23171
rect 20913 23137 20947 23171
rect 22845 23137 22879 23171
rect 24593 23137 24627 23171
rect 10241 23069 10275 23103
rect 12725 23069 12759 23103
rect 15301 23069 15335 23103
rect 22385 23069 22419 23103
rect 23121 23069 23155 23103
rect 12541 22933 12575 22967
rect 16497 22933 16531 22967
rect 18061 22933 18095 22967
rect 19349 22933 19383 22967
rect 22569 22933 22603 22967
rect 23765 22933 23799 22967
rect 24133 22933 24167 22967
rect 10977 22729 11011 22763
rect 12725 22729 12759 22763
rect 13093 22729 13127 22763
rect 15945 22729 15979 22763
rect 18705 22729 18739 22763
rect 21557 22729 21591 22763
rect 23029 22729 23063 22763
rect 23489 22729 23523 22763
rect 25421 22729 25455 22763
rect 14289 22661 14323 22695
rect 16497 22661 16531 22695
rect 17509 22661 17543 22695
rect 22109 22661 22143 22695
rect 23765 22661 23799 22695
rect 14105 22593 14139 22627
rect 14749 22593 14783 22627
rect 14841 22593 14875 22627
rect 21833 22593 21867 22627
rect 24133 22593 24167 22627
rect 24317 22593 24351 22627
rect 13737 22525 13771 22559
rect 16773 22525 16807 22559
rect 19441 22525 19475 22559
rect 19533 22525 19567 22559
rect 24685 22525 24719 22559
rect 25237 22525 25271 22559
rect 14749 22457 14783 22491
rect 16221 22457 16255 22491
rect 17049 22457 17083 22491
rect 19800 22457 19834 22491
rect 22385 22457 22419 22491
rect 22569 22457 22603 22491
rect 22661 22457 22695 22491
rect 25881 22457 25915 22491
rect 10241 22389 10275 22423
rect 10517 22389 10551 22423
rect 16957 22389 16991 22423
rect 18981 22389 19015 22423
rect 20913 22389 20947 22423
rect 24225 22389 24259 22423
rect 10977 22185 11011 22219
rect 14657 22185 14691 22219
rect 17233 22185 17267 22219
rect 19349 22185 19383 22219
rect 19809 22185 19843 22219
rect 21097 22185 21131 22219
rect 23765 22185 23799 22219
rect 14197 22117 14231 22151
rect 18797 22117 18831 22151
rect 19717 22117 19751 22151
rect 22937 22117 22971 22151
rect 16497 22049 16531 22083
rect 17049 22049 17083 22083
rect 22753 22049 22787 22083
rect 23029 22049 23063 22083
rect 24205 22049 24239 22083
rect 10885 21981 10919 22015
rect 11069 21981 11103 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 17325 21981 17359 22015
rect 18705 21981 18739 22015
rect 18889 21981 18923 22015
rect 22109 21981 22143 22015
rect 23949 21981 23983 22015
rect 16773 21913 16807 21947
rect 18061 21913 18095 21947
rect 22477 21913 22511 21947
rect 10517 21845 10551 21879
rect 13737 21845 13771 21879
rect 18337 21845 18371 21879
rect 21741 21845 21775 21879
rect 25329 21845 25363 21879
rect 9873 21641 9907 21675
rect 13645 21641 13679 21675
rect 15761 21641 15795 21675
rect 17785 21641 17819 21675
rect 18613 21641 18647 21675
rect 21557 21641 21591 21675
rect 22109 21641 22143 21675
rect 10425 21573 10459 21607
rect 13001 21573 13035 21607
rect 16773 21573 16807 21607
rect 17049 21573 17083 21607
rect 19257 21573 19291 21607
rect 23121 21573 23155 21607
rect 10149 21505 10183 21539
rect 10977 21505 11011 21539
rect 11345 21505 11379 21539
rect 13369 21505 13403 21539
rect 19073 21505 19107 21539
rect 19809 21505 19843 21539
rect 22661 21505 22695 21539
rect 9505 21437 9539 21471
rect 10701 21437 10735 21471
rect 12081 21437 12115 21471
rect 14381 21437 14415 21471
rect 14648 21437 14682 21471
rect 19533 21437 19567 21471
rect 20177 21437 20211 21471
rect 23489 21437 23523 21471
rect 23673 21437 23707 21471
rect 10885 21369 10919 21403
rect 19717 21369 19751 21403
rect 21005 21369 21039 21403
rect 21925 21369 21959 21403
rect 22385 21369 22419 21403
rect 23918 21369 23952 21403
rect 11713 21301 11747 21335
rect 14197 21301 14231 21335
rect 17509 21301 17543 21335
rect 18061 21301 18095 21335
rect 22569 21301 22603 21335
rect 25053 21301 25087 21335
rect 11805 21097 11839 21131
rect 14013 21097 14047 21131
rect 14565 21097 14599 21131
rect 15853 21097 15887 21131
rect 16497 21097 16531 21131
rect 18889 21097 18923 21131
rect 19441 21097 19475 21131
rect 21741 21097 21775 21131
rect 24317 21097 24351 21131
rect 24777 21097 24811 21131
rect 10692 21029 10726 21063
rect 13829 21029 13863 21063
rect 21189 21029 21223 21063
rect 22109 21029 22143 21063
rect 22477 21029 22511 21063
rect 23213 21029 23247 21063
rect 23305 21029 23339 21063
rect 13001 20961 13035 20995
rect 17509 20961 17543 20995
rect 17776 20961 17810 20995
rect 20913 20961 20947 20995
rect 24593 20961 24627 20995
rect 10425 20893 10459 20927
rect 14105 20893 14139 20927
rect 16497 20893 16531 20927
rect 16589 20893 16623 20927
rect 23121 20893 23155 20927
rect 13369 20825 13403 20859
rect 22753 20825 22787 20859
rect 13553 20757 13587 20791
rect 16037 20757 16071 20791
rect 16957 20757 16991 20791
rect 20637 20757 20671 20791
rect 23949 20757 23983 20791
rect 13001 20553 13035 20587
rect 14841 20553 14875 20587
rect 15945 20553 15979 20587
rect 17509 20553 17543 20587
rect 17785 20553 17819 20587
rect 20637 20553 20671 20587
rect 21557 20553 21591 20587
rect 23397 20553 23431 20587
rect 25053 20553 25087 20587
rect 16497 20485 16531 20519
rect 16313 20417 16347 20451
rect 16957 20417 16991 20451
rect 18061 20417 18095 20451
rect 13461 20349 13495 20383
rect 13728 20349 13762 20383
rect 15577 20349 15611 20383
rect 18328 20349 18362 20383
rect 10517 20281 10551 20315
rect 16957 20281 16991 20315
rect 17049 20281 17083 20315
rect 20453 20281 20487 20315
rect 20913 20281 20947 20315
rect 21189 20281 21223 20315
rect 24317 20281 24351 20315
rect 10885 20213 10919 20247
rect 13277 20213 13311 20247
rect 19441 20213 19475 20247
rect 21097 20213 21131 20247
rect 22753 20213 22787 20247
rect 23029 20213 23063 20247
rect 24501 20213 24535 20247
rect 11805 20009 11839 20043
rect 12817 20009 12851 20043
rect 14289 20009 14323 20043
rect 18889 20009 18923 20043
rect 19809 20009 19843 20043
rect 20637 20009 20671 20043
rect 23121 20009 23155 20043
rect 24041 20009 24075 20043
rect 13461 19941 13495 19975
rect 13553 19941 13587 19975
rect 15568 19941 15602 19975
rect 18337 19941 18371 19975
rect 21986 19941 22020 19975
rect 24777 19941 24811 19975
rect 10692 19873 10726 19907
rect 13921 19873 13955 19907
rect 15301 19873 15335 19907
rect 17601 19873 17635 19907
rect 21741 19873 21775 19907
rect 24593 19873 24627 19907
rect 10425 19805 10459 19839
rect 13461 19805 13495 19839
rect 18245 19805 18279 19839
rect 18429 19805 18463 19839
rect 24869 19805 24903 19839
rect 17877 19737 17911 19771
rect 23765 19737 23799 19771
rect 13001 19669 13035 19703
rect 16681 19669 16715 19703
rect 24317 19669 24351 19703
rect 12909 19465 12943 19499
rect 15301 19465 15335 19499
rect 15669 19465 15703 19499
rect 16129 19465 16163 19499
rect 19441 19465 19475 19499
rect 23949 19465 23983 19499
rect 10333 19397 10367 19431
rect 9965 19261 9999 19295
rect 10867 19261 10901 19295
rect 13185 19261 13219 19295
rect 17141 19261 17175 19295
rect 17509 19261 17543 19295
rect 18429 19261 18463 19295
rect 19073 19261 19107 19295
rect 20545 19261 20579 19295
rect 20729 19261 20763 19295
rect 24140 19261 24174 19295
rect 10609 19193 10643 19227
rect 11161 19193 11195 19227
rect 11437 19193 11471 19227
rect 12265 19193 12299 19227
rect 13430 19193 13464 19227
rect 17785 19193 17819 19227
rect 18135 19193 18169 19227
rect 18705 19193 18739 19227
rect 20269 19193 20303 19227
rect 20996 19193 21030 19227
rect 24400 19193 24434 19227
rect 11345 19125 11379 19159
rect 11897 19125 11931 19159
rect 14565 19125 14599 19159
rect 18613 19125 18647 19159
rect 22109 19125 22143 19159
rect 22661 19125 22695 19159
rect 23489 19125 23523 19159
rect 25513 19125 25547 19159
rect 13737 18921 13771 18955
rect 21925 18921 21959 18955
rect 25145 18921 25179 18955
rect 13553 18853 13587 18887
rect 13829 18853 13863 18887
rect 16926 18853 16960 18887
rect 21465 18853 21499 18887
rect 10968 18785 11002 18819
rect 13001 18785 13035 18819
rect 24021 18785 24055 18819
rect 10701 18717 10735 18751
rect 15393 18717 15427 18751
rect 16681 18717 16715 18751
rect 21465 18717 21499 18751
rect 21557 18717 21591 18751
rect 23765 18717 23799 18751
rect 21005 18649 21039 18683
rect 10425 18581 10459 18615
rect 12081 18581 12115 18615
rect 13277 18581 13311 18615
rect 18061 18581 18095 18615
rect 18613 18581 18647 18615
rect 9873 18377 9907 18411
rect 12909 18377 12943 18411
rect 14013 18377 14047 18411
rect 15209 18377 15243 18411
rect 17049 18377 17083 18411
rect 21005 18377 21039 18411
rect 23489 18377 23523 18411
rect 24317 18377 24351 18411
rect 10793 18309 10827 18343
rect 13277 18309 13311 18343
rect 15393 18309 15427 18343
rect 16773 18309 16807 18343
rect 24501 18309 24535 18343
rect 11345 18241 11379 18275
rect 15761 18241 15795 18275
rect 24869 18241 24903 18275
rect 25053 18241 25087 18275
rect 25421 18173 25455 18207
rect 10241 18105 10275 18139
rect 11069 18105 11103 18139
rect 11253 18105 11287 18139
rect 14841 18105 14875 18139
rect 15945 18105 15979 18139
rect 24961 18105 24995 18139
rect 10609 18037 10643 18071
rect 11805 18037 11839 18071
rect 13553 18037 13587 18071
rect 15853 18037 15887 18071
rect 18705 18037 18739 18071
rect 21373 18037 21407 18071
rect 21649 18037 21683 18071
rect 23857 18037 23891 18071
rect 10793 17833 10827 17867
rect 11253 17833 11287 17867
rect 13369 17833 13403 17867
rect 15485 17833 15519 17867
rect 18153 17833 18187 17867
rect 24685 17833 24719 17867
rect 13829 17765 13863 17799
rect 14013 17765 14047 17799
rect 21465 17765 21499 17799
rect 23765 17765 23799 17799
rect 18593 17697 18627 17731
rect 23581 17697 23615 17731
rect 14105 17629 14139 17663
rect 18337 17629 18371 17663
rect 21373 17629 21407 17663
rect 21557 17629 21591 17663
rect 23857 17629 23891 17663
rect 24317 17629 24351 17663
rect 24777 17629 24811 17663
rect 13553 17493 13587 17527
rect 16405 17493 16439 17527
rect 19717 17493 19751 17527
rect 21005 17493 21039 17527
rect 23305 17493 23339 17527
rect 17509 17289 17543 17323
rect 19073 17289 19107 17323
rect 19533 17289 19567 17323
rect 21005 17289 21039 17323
rect 22845 17289 22879 17323
rect 16129 17221 16163 17255
rect 16405 17221 16439 17255
rect 18153 17221 18187 17255
rect 23857 17221 23891 17255
rect 16865 17153 16899 17187
rect 17877 17153 17911 17187
rect 18613 17153 18647 17187
rect 19625 17153 19659 17187
rect 21557 17153 21591 17187
rect 24225 17153 24259 17187
rect 13001 17085 13035 17119
rect 13268 17085 13302 17119
rect 23213 17085 23247 17119
rect 12265 17017 12299 17051
rect 16865 17017 16899 17051
rect 16957 17017 16991 17051
rect 18613 17017 18647 17051
rect 18705 17017 18739 17051
rect 19870 17017 19904 17051
rect 24409 17017 24443 17051
rect 24777 17017 24811 17051
rect 12817 16949 12851 16983
rect 14381 16949 14415 16983
rect 15025 16949 15059 16983
rect 15853 16949 15887 16983
rect 21925 16949 21959 16983
rect 22109 16949 22143 16983
rect 24317 16949 24351 16983
rect 12265 16745 12299 16779
rect 13277 16745 13311 16779
rect 13921 16745 13955 16779
rect 18153 16745 18187 16779
rect 19625 16745 19659 16779
rect 23857 16745 23891 16779
rect 25329 16745 25363 16779
rect 13737 16677 13771 16711
rect 14013 16677 14047 16711
rect 16006 16677 16040 16711
rect 18797 16677 18831 16711
rect 20729 16677 20763 16711
rect 21250 16677 21284 16711
rect 23305 16677 23339 16711
rect 24216 16677 24250 16711
rect 10885 16609 10919 16643
rect 11152 16609 11186 16643
rect 18613 16609 18647 16643
rect 23949 16609 23983 16643
rect 15761 16541 15795 16575
rect 18889 16541 18923 16575
rect 21012 16541 21046 16575
rect 17141 16473 17175 16507
rect 13461 16405 13495 16439
rect 18337 16405 18371 16439
rect 22385 16405 22419 16439
rect 11253 16201 11287 16235
rect 13093 16201 13127 16235
rect 15577 16201 15611 16235
rect 16589 16201 16623 16235
rect 18337 16201 18371 16235
rect 18981 16201 19015 16235
rect 21005 16201 21039 16235
rect 23121 16201 23155 16235
rect 23489 16201 23523 16235
rect 25421 16201 25455 16235
rect 25881 16201 25915 16235
rect 10885 16133 10919 16167
rect 21557 16133 21591 16167
rect 23765 16133 23799 16167
rect 24685 16133 24719 16167
rect 16865 16065 16899 16099
rect 18613 16065 18647 16099
rect 22017 16065 22051 16099
rect 24317 16065 24351 16099
rect 14197 15997 14231 16031
rect 20729 15997 20763 16031
rect 24041 15997 24075 16031
rect 25053 15997 25087 16031
rect 25237 15997 25271 16031
rect 13461 15929 13495 15963
rect 14442 15929 14476 15963
rect 22017 15929 22051 15963
rect 22109 15929 22143 15963
rect 24225 15929 24259 15963
rect 14105 15861 14139 15895
rect 16221 15861 16255 15895
rect 13461 15657 13495 15691
rect 14289 15657 14323 15691
rect 16773 15657 16807 15691
rect 21097 15657 21131 15691
rect 21925 15657 21959 15691
rect 23949 15657 23983 15691
rect 24501 15657 24535 15691
rect 25237 15657 25271 15691
rect 16865 15589 16899 15623
rect 18061 15589 18095 15623
rect 21557 15589 21591 15623
rect 17785 15521 17819 15555
rect 22836 15521 22870 15555
rect 25053 15521 25087 15555
rect 16773 15453 16807 15487
rect 19073 15453 19107 15487
rect 22569 15453 22603 15487
rect 16313 15317 16347 15351
rect 18613 15317 18647 15351
rect 20177 15317 20211 15351
rect 16405 15113 16439 15147
rect 16681 15113 16715 15147
rect 17509 15113 17543 15147
rect 18613 15113 18647 15147
rect 19901 15113 19935 15147
rect 21465 15113 21499 15147
rect 22569 15113 22603 15147
rect 22937 15113 22971 15147
rect 25053 15113 25087 15147
rect 13185 14977 13219 15011
rect 15853 14977 15887 15011
rect 18429 14977 18463 15011
rect 19073 14977 19107 15011
rect 20085 14977 20119 15011
rect 12909 14909 12943 14943
rect 13645 14909 13679 14943
rect 15577 14909 15611 14943
rect 19165 14841 19199 14875
rect 20352 14841 20386 14875
rect 15485 14773 15519 14807
rect 16865 14773 16899 14807
rect 17877 14773 17911 14807
rect 19073 14773 19107 14807
rect 16313 14569 16347 14603
rect 21465 14569 21499 14603
rect 24777 14569 24811 14603
rect 13553 14501 13587 14535
rect 14197 14501 14231 14535
rect 16773 14501 16807 14535
rect 16957 14501 16991 14535
rect 21281 14501 21315 14535
rect 12633 14433 12667 14467
rect 14013 14433 14047 14467
rect 18337 14433 18371 14467
rect 18604 14433 18638 14467
rect 24593 14433 24627 14467
rect 14289 14365 14323 14399
rect 17049 14365 17083 14399
rect 21557 14365 21591 14399
rect 13737 14297 13771 14331
rect 16497 14297 16531 14331
rect 21005 14297 21039 14331
rect 19717 14229 19751 14263
rect 12817 14025 12851 14059
rect 14289 14025 14323 14059
rect 14841 14025 14875 14059
rect 15209 14025 15243 14059
rect 17693 14025 17727 14059
rect 18337 14025 18371 14059
rect 19349 14025 19383 14059
rect 20913 14025 20947 14059
rect 21465 14025 21499 14059
rect 21833 14025 21867 14059
rect 24685 14025 24719 14059
rect 17325 13957 17359 13991
rect 18705 13957 18739 13991
rect 12909 13889 12943 13923
rect 15393 13889 15427 13923
rect 19533 13889 19567 13923
rect 19800 13821 19834 13855
rect 13176 13753 13210 13787
rect 15638 13753 15672 13787
rect 16773 13685 16807 13719
rect 13553 13481 13587 13515
rect 15485 13481 15519 13515
rect 16405 13481 16439 13515
rect 18245 13481 18279 13515
rect 19533 13481 19567 13515
rect 21189 13481 21223 13515
rect 14197 13413 14231 13447
rect 17110 13413 17144 13447
rect 13001 13345 13035 13379
rect 24593 13345 24627 13379
rect 14197 13277 14231 13311
rect 14289 13277 14323 13311
rect 16865 13277 16899 13311
rect 13737 13209 13771 13243
rect 24777 13209 24811 13243
rect 16497 12937 16531 12971
rect 17417 12937 17451 12971
rect 24685 12937 24719 12971
rect 13093 12801 13127 12835
rect 16313 12801 16347 12835
rect 17049 12801 17083 12835
rect 15945 12733 15979 12767
rect 13001 12665 13035 12699
rect 13360 12665 13394 12699
rect 16773 12665 16807 12699
rect 16957 12665 16991 12699
rect 14473 12597 14507 12631
rect 13093 12393 13127 12427
rect 13737 12393 13771 12427
rect 14473 12393 14507 12427
rect 16865 12393 16899 12427
rect 24777 12393 24811 12427
rect 14013 12325 14047 12359
rect 16405 12325 16439 12359
rect 24593 12257 24627 12291
rect 13277 11849 13311 11883
rect 24685 11849 24719 11883
rect 12725 11645 12759 11679
rect 12909 11509 12943 11543
rect 12081 11169 12115 11203
rect 12265 11033 12299 11067
rect 11805 10761 11839 10795
rect 12173 10761 12207 10795
rect 11253 10557 11287 10591
rect 11437 10421 11471 10455
rect 10701 10081 10735 10115
rect 10885 9945 10919 9979
rect 10977 9673 11011 9707
rect 10241 9605 10275 9639
rect 10057 9469 10091 9503
rect 10609 9469 10643 9503
rect 24593 9469 24627 9503
rect 25145 9469 25179 9503
rect 24777 9333 24811 9367
rect 24593 9061 24627 9095
rect 9689 8993 9723 9027
rect 24317 8993 24351 9027
rect 9873 8857 9907 8891
rect 9689 8585 9723 8619
rect 24961 8585 24995 8619
rect 25329 8517 25363 8551
rect 24593 8449 24627 8483
rect 23857 8381 23891 8415
rect 24133 8381 24167 8415
rect 25145 8381 25179 8415
rect 25697 8381 25731 8415
rect 19349 7905 19383 7939
rect 22937 7905 22971 7939
rect 23213 7905 23247 7939
rect 24317 7905 24351 7939
rect 19625 7837 19659 7871
rect 24501 7701 24535 7735
rect 19349 7497 19383 7531
rect 22937 7497 22971 7531
rect 24317 7497 24351 7531
rect 24593 7293 24627 7327
rect 25145 7293 25179 7327
rect 24777 7157 24811 7191
rect 23673 6817 23707 6851
rect 23949 6817 23983 6851
rect 24961 6817 24995 6851
rect 25145 6613 25179 6647
rect 23489 6409 23523 6443
rect 24777 6409 24811 6443
rect 14933 6205 14967 6239
rect 15669 6205 15703 6239
rect 23673 6205 23707 6239
rect 23949 6205 23983 6239
rect 24961 6205 24995 6239
rect 25513 6205 25547 6239
rect 15209 6137 15243 6171
rect 24409 6137 24443 6171
rect 25145 6069 25179 6103
rect 23673 5729 23707 5763
rect 24961 5729 24995 5763
rect 23857 5661 23891 5695
rect 25145 5525 25179 5559
rect 23489 5321 23523 5355
rect 24869 5321 24903 5355
rect 23673 5117 23707 5151
rect 24409 5117 24443 5151
rect 24961 5117 24995 5151
rect 23949 5049 23983 5083
rect 25513 5049 25547 5083
rect 25145 4981 25179 5015
rect 23489 4641 23523 4675
rect 24593 4641 24627 4675
rect 23673 4437 23707 4471
rect 24777 4437 24811 4471
rect 23857 4233 23891 4267
rect 24593 4029 24627 4063
rect 25145 4029 25179 4063
rect 24409 3893 24443 3927
rect 24777 3893 24811 3927
rect 23765 3621 23799 3655
rect 23489 3553 23523 3587
rect 24777 3553 24811 3587
rect 24961 3349 24995 3383
rect 23121 3145 23155 3179
rect 24869 3145 24903 3179
rect 23489 3077 23523 3111
rect 23949 3009 23983 3043
rect 25145 3009 25179 3043
rect 22293 2941 22327 2975
rect 23673 2941 23707 2975
rect 24409 2941 24443 2975
rect 24961 2941 24995 2975
rect 25697 2941 25731 2975
rect 22569 2873 22603 2907
rect 22845 2465 22879 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 23489 2397 23523 2431
rect 24225 2397 24259 2431
rect 23029 2261 23063 2295
rect 25513 2261 25547 2295
<< metal1 >>
rect 20346 26936 20352 26988
rect 20404 26976 20410 26988
rect 24762 26976 24768 26988
rect 20404 26948 24768 26976
rect 20404 26936 20410 26948
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 19978 26392 19984 26444
rect 20036 26432 20042 26444
rect 24762 26432 24768 26444
rect 20036 26404 24768 26432
rect 20036 26392 20042 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 21542 25440 21548 25492
rect 21600 25480 21606 25492
rect 23017 25483 23075 25489
rect 23017 25480 23029 25483
rect 21600 25452 23029 25480
rect 21600 25440 21606 25452
rect 23017 25449 23029 25452
rect 23063 25449 23075 25483
rect 23017 25443 23075 25449
rect 23566 25440 23572 25492
rect 23624 25480 23630 25492
rect 24765 25483 24823 25489
rect 24765 25480 24777 25483
rect 23624 25452 24777 25480
rect 23624 25440 23630 25452
rect 24765 25449 24777 25452
rect 24811 25449 24823 25483
rect 24765 25443 24823 25449
rect 18690 25372 18696 25424
rect 18748 25412 18754 25424
rect 19429 25415 19487 25421
rect 19429 25412 19441 25415
rect 18748 25384 19441 25412
rect 18748 25372 18754 25384
rect 19429 25381 19441 25384
rect 19475 25381 19487 25415
rect 19429 25375 19487 25381
rect 22833 25347 22891 25353
rect 22833 25313 22845 25347
rect 22879 25344 22891 25347
rect 23198 25344 23204 25356
rect 22879 25316 23204 25344
rect 22879 25313 22891 25316
rect 22833 25307 22891 25313
rect 23198 25304 23204 25316
rect 23256 25304 23262 25356
rect 24581 25347 24639 25353
rect 24581 25313 24593 25347
rect 24627 25344 24639 25347
rect 24762 25344 24768 25356
rect 24627 25316 24768 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 24762 25304 24768 25316
rect 24820 25304 24826 25356
rect 19426 25276 19432 25288
rect 19387 25248 19432 25276
rect 19426 25236 19432 25248
rect 19484 25236 19490 25288
rect 19521 25279 19579 25285
rect 19521 25245 19533 25279
rect 19567 25276 19579 25279
rect 19610 25276 19616 25288
rect 19567 25248 19616 25276
rect 19567 25245 19579 25248
rect 19521 25239 19579 25245
rect 19610 25236 19616 25248
rect 19668 25236 19674 25288
rect 14277 25143 14335 25149
rect 14277 25109 14289 25143
rect 14323 25140 14335 25143
rect 14826 25140 14832 25152
rect 14323 25112 14832 25140
rect 14323 25109 14335 25112
rect 14277 25103 14335 25109
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 18969 25143 19027 25149
rect 18969 25109 18981 25143
rect 19015 25140 19027 25143
rect 19334 25140 19340 25152
rect 19015 25112 19340 25140
rect 19015 25109 19027 25112
rect 18969 25103 19027 25109
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 19337 24939 19395 24945
rect 19337 24905 19349 24939
rect 19383 24936 19395 24939
rect 19426 24936 19432 24948
rect 19383 24908 19432 24936
rect 19383 24905 19395 24908
rect 19337 24899 19395 24905
rect 19426 24896 19432 24908
rect 19484 24936 19490 24948
rect 20625 24939 20683 24945
rect 20625 24936 20637 24939
rect 19484 24908 20637 24936
rect 19484 24896 19490 24908
rect 20625 24905 20637 24908
rect 20671 24905 20683 24939
rect 20625 24899 20683 24905
rect 23658 24896 23664 24948
rect 23716 24936 23722 24948
rect 24762 24936 24768 24948
rect 23716 24908 24768 24936
rect 23716 24896 23722 24908
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 19610 24868 19616 24880
rect 19260 24840 19616 24868
rect 9674 24760 9680 24812
rect 9732 24800 9738 24812
rect 10134 24800 10140 24812
rect 9732 24772 10140 24800
rect 9732 24760 9738 24772
rect 10134 24760 10140 24772
rect 10192 24760 10198 24812
rect 14826 24800 14832 24812
rect 14787 24772 14832 24800
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 18417 24803 18475 24809
rect 18417 24769 18429 24803
rect 18463 24800 18475 24803
rect 19260 24800 19288 24840
rect 19610 24828 19616 24840
rect 19668 24868 19674 24880
rect 20070 24868 20076 24880
rect 19668 24840 20076 24868
rect 19668 24828 19674 24840
rect 20070 24828 20076 24840
rect 20128 24828 20134 24880
rect 24670 24868 24676 24880
rect 20364 24840 24676 24868
rect 18463 24772 19288 24800
rect 18463 24769 18475 24772
rect 18417 24763 18475 24769
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 14553 24735 14611 24741
rect 14553 24732 14565 24735
rect 14424 24704 14565 24732
rect 14424 24692 14430 24704
rect 14553 24701 14565 24704
rect 14599 24701 14611 24735
rect 14553 24695 14611 24701
rect 18690 24692 18696 24744
rect 18748 24732 18754 24744
rect 20257 24735 20315 24741
rect 20257 24732 20269 24735
rect 18748 24704 20269 24732
rect 18748 24692 18754 24704
rect 20257 24701 20269 24704
rect 20303 24701 20315 24735
rect 20257 24695 20315 24701
rect 13998 24664 14004 24676
rect 13959 24636 14004 24664
rect 13998 24624 14004 24636
rect 14056 24624 14062 24676
rect 14259 24667 14317 24673
rect 14259 24633 14271 24667
rect 14305 24664 14317 24667
rect 14458 24664 14464 24676
rect 14305 24636 14464 24664
rect 14305 24633 14317 24636
rect 14259 24627 14317 24633
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 19613 24667 19671 24673
rect 19613 24664 19625 24667
rect 18708 24636 19625 24664
rect 14016 24596 14044 24624
rect 14737 24599 14795 24605
rect 14737 24596 14749 24599
rect 14016 24568 14749 24596
rect 14737 24565 14749 24568
rect 14783 24565 14795 24599
rect 14737 24559 14795 24565
rect 18506 24556 18512 24608
rect 18564 24596 18570 24608
rect 18708 24605 18736 24636
rect 19613 24633 19625 24636
rect 19659 24664 19671 24667
rect 19702 24664 19708 24676
rect 19659 24636 19708 24664
rect 19659 24633 19671 24636
rect 19613 24627 19671 24633
rect 19702 24624 19708 24636
rect 19760 24624 19766 24676
rect 19889 24667 19947 24673
rect 19889 24633 19901 24667
rect 19935 24664 19947 24667
rect 20162 24664 20168 24676
rect 19935 24636 20168 24664
rect 19935 24633 19947 24636
rect 19889 24627 19947 24633
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 18693 24599 18751 24605
rect 18693 24596 18705 24599
rect 18564 24568 18705 24596
rect 18564 24556 18570 24568
rect 18693 24565 18705 24568
rect 18739 24565 18751 24599
rect 19150 24596 19156 24608
rect 19063 24568 19156 24596
rect 18693 24559 18751 24565
rect 19150 24556 19156 24568
rect 19208 24596 19214 24608
rect 19797 24599 19855 24605
rect 19797 24596 19809 24599
rect 19208 24568 19809 24596
rect 19208 24556 19214 24568
rect 19797 24565 19809 24568
rect 19843 24596 19855 24599
rect 20364 24596 20392 24840
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 24780 24800 24808 24896
rect 25133 24803 25191 24809
rect 25133 24800 25145 24803
rect 24780 24772 25145 24800
rect 25133 24769 25145 24772
rect 25179 24769 25191 24803
rect 25133 24763 25191 24769
rect 22465 24735 22523 24741
rect 22465 24732 22477 24735
rect 22388 24704 22477 24732
rect 22388 24608 22416 24704
rect 22465 24701 22477 24704
rect 22511 24701 22523 24735
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 22465 24695 22523 24701
rect 24136 24704 24593 24732
rect 22370 24596 22376 24608
rect 19843 24568 20392 24596
rect 22331 24568 22376 24596
rect 19843 24565 19855 24568
rect 19797 24559 19855 24565
rect 22370 24556 22376 24568
rect 22428 24556 22434 24608
rect 22649 24599 22707 24605
rect 22649 24565 22661 24599
rect 22695 24596 22707 24599
rect 22922 24596 22928 24608
rect 22695 24568 22928 24596
rect 22695 24565 22707 24568
rect 22649 24559 22707 24565
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 23109 24599 23167 24605
rect 23109 24565 23121 24599
rect 23155 24596 23167 24599
rect 23198 24596 23204 24608
rect 23155 24568 23204 24596
rect 23155 24565 23167 24568
rect 23109 24559 23167 24565
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 24026 24556 24032 24608
rect 24084 24596 24090 24608
rect 24136 24596 24164 24704
rect 24581 24701 24593 24704
rect 24627 24701 24639 24735
rect 24581 24695 24639 24701
rect 24210 24624 24216 24676
rect 24268 24664 24274 24676
rect 24268 24636 24808 24664
rect 24268 24624 24274 24636
rect 24780 24605 24808 24636
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 24084 24568 24409 24596
rect 24084 24556 24090 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24397 24559 24455 24565
rect 24765 24599 24823 24605
rect 24765 24565 24777 24599
rect 24811 24565 24823 24599
rect 24765 24559 24823 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 13817 24395 13875 24401
rect 13817 24361 13829 24395
rect 13863 24392 13875 24395
rect 14274 24392 14280 24404
rect 13863 24364 14280 24392
rect 13863 24361 13875 24364
rect 13817 24355 13875 24361
rect 14274 24352 14280 24364
rect 14332 24352 14338 24404
rect 14645 24395 14703 24401
rect 14645 24361 14657 24395
rect 14691 24392 14703 24395
rect 14826 24392 14832 24404
rect 14691 24364 14832 24392
rect 14691 24361 14703 24364
rect 14645 24355 14703 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 15562 24392 15568 24404
rect 15519 24364 15568 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 20254 24352 20260 24404
rect 20312 24392 20318 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20312 24364 21097 24392
rect 20312 24352 20318 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 25406 24392 25412 24404
rect 25367 24364 25412 24392
rect 21085 24355 21143 24361
rect 25406 24352 25412 24364
rect 25464 24352 25470 24404
rect 18598 24284 18604 24336
rect 18656 24324 18662 24336
rect 19153 24327 19211 24333
rect 19153 24324 19165 24327
rect 18656 24296 19165 24324
rect 18656 24284 18662 24296
rect 19153 24293 19165 24296
rect 19199 24293 19211 24327
rect 19153 24287 19211 24293
rect 10318 24216 10324 24268
rect 10376 24256 10382 24268
rect 11238 24256 11244 24268
rect 10376 24228 11244 24256
rect 10376 24216 10382 24228
rect 11238 24216 11244 24228
rect 11296 24256 11302 24268
rect 11405 24259 11463 24265
rect 11405 24256 11417 24259
rect 11296 24228 11417 24256
rect 11296 24216 11302 24228
rect 11405 24225 11417 24228
rect 11451 24225 11463 24259
rect 13633 24259 13691 24265
rect 13633 24256 13645 24259
rect 11405 24219 11463 24225
rect 13464 24228 13645 24256
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11149 24191 11207 24197
rect 11149 24188 11161 24191
rect 11112 24160 11161 24188
rect 11112 24148 11118 24160
rect 11149 24157 11161 24160
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 10505 24055 10563 24061
rect 10505 24021 10517 24055
rect 10551 24052 10563 24055
rect 10778 24052 10784 24064
rect 10551 24024 10784 24052
rect 10551 24021 10563 24024
rect 10505 24015 10563 24021
rect 10778 24012 10784 24024
rect 10836 24012 10842 24064
rect 10873 24055 10931 24061
rect 10873 24021 10885 24055
rect 10919 24052 10931 24055
rect 11422 24052 11428 24064
rect 10919 24024 11428 24052
rect 10919 24021 10931 24024
rect 10873 24015 10931 24021
rect 11422 24012 11428 24024
rect 11480 24052 11486 24064
rect 12526 24052 12532 24064
rect 11480 24024 12532 24052
rect 11480 24012 11486 24024
rect 12526 24012 12532 24024
rect 12584 24012 12590 24064
rect 13170 24012 13176 24064
rect 13228 24052 13234 24064
rect 13464 24061 13492 24228
rect 13633 24225 13645 24228
rect 13679 24225 13691 24259
rect 13633 24219 13691 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 15838 24256 15844 24268
rect 15335 24228 15844 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 15838 24216 15844 24228
rect 15896 24216 15902 24268
rect 20901 24259 20959 24265
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 21358 24256 21364 24268
rect 20947 24228 21364 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21358 24216 21364 24228
rect 21416 24216 21422 24268
rect 23014 24265 23020 24268
rect 23008 24219 23020 24265
rect 23072 24256 23078 24268
rect 25222 24256 25228 24268
rect 23072 24228 23108 24256
rect 25183 24228 25228 24256
rect 23014 24216 23020 24219
rect 23072 24216 23078 24228
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 19058 24188 19064 24200
rect 19019 24160 19064 24188
rect 19058 24148 19064 24160
rect 19116 24148 19122 24200
rect 19245 24191 19303 24197
rect 19245 24157 19257 24191
rect 19291 24188 19303 24191
rect 22738 24188 22744 24200
rect 19291 24160 19748 24188
rect 22699 24160 22744 24188
rect 19291 24157 19303 24160
rect 19245 24151 19303 24157
rect 18690 24120 18696 24132
rect 18651 24092 18696 24120
rect 18690 24080 18696 24092
rect 18748 24080 18754 24132
rect 13449 24055 13507 24061
rect 13449 24052 13461 24055
rect 13228 24024 13461 24052
rect 13228 24012 13234 24024
rect 13449 24021 13461 24024
rect 13495 24021 13507 24055
rect 13449 24015 13507 24021
rect 14277 24055 14335 24061
rect 14277 24021 14289 24055
rect 14323 24052 14335 24055
rect 14366 24052 14372 24064
rect 14323 24024 14372 24052
rect 14323 24021 14335 24024
rect 14277 24015 14335 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 19610 24012 19616 24064
rect 19668 24052 19674 24064
rect 19720 24061 19748 24160
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 19705 24055 19763 24061
rect 19705 24052 19717 24055
rect 19668 24024 19717 24052
rect 19668 24012 19674 24024
rect 19705 24021 19717 24024
rect 19751 24052 19763 24055
rect 20073 24055 20131 24061
rect 20073 24052 20085 24055
rect 19751 24024 20085 24052
rect 19751 24021 19763 24024
rect 19705 24015 19763 24021
rect 20073 24021 20085 24024
rect 20119 24052 20131 24055
rect 20162 24052 20168 24064
rect 20119 24024 20168 24052
rect 20119 24021 20131 24024
rect 20073 24015 20131 24021
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 24118 24052 24124 24064
rect 24079 24024 24124 24052
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 10318 23848 10324 23860
rect 10279 23820 10324 23848
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 16850 23848 16856 23860
rect 11296 23820 13124 23848
rect 16811 23820 16856 23848
rect 11296 23808 11302 23820
rect 9858 23740 9864 23792
rect 9916 23780 9922 23792
rect 10873 23783 10931 23789
rect 10873 23780 10885 23783
rect 9916 23752 10885 23780
rect 9916 23740 9922 23752
rect 10873 23749 10885 23752
rect 10919 23749 10931 23783
rect 12529 23783 12587 23789
rect 12529 23780 12541 23783
rect 10873 23743 10931 23749
rect 11532 23752 12541 23780
rect 11422 23712 11428 23724
rect 11383 23684 11428 23712
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 11532 23644 11560 23752
rect 12529 23749 12541 23752
rect 12575 23749 12587 23783
rect 12529 23743 12587 23749
rect 12986 23712 12992 23724
rect 12947 23684 12992 23712
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 13096 23721 13124 23820
rect 16850 23808 16856 23820
rect 16908 23808 16914 23860
rect 20898 23808 20904 23860
rect 20956 23848 20962 23860
rect 22005 23851 22063 23857
rect 22005 23848 22017 23851
rect 20956 23820 22017 23848
rect 20956 23808 20962 23820
rect 22005 23817 22017 23820
rect 22051 23817 22063 23851
rect 22738 23848 22744 23860
rect 22699 23820 22744 23848
rect 22005 23811 22063 23817
rect 22738 23808 22744 23820
rect 22796 23808 22802 23860
rect 23014 23808 23020 23860
rect 23072 23848 23078 23860
rect 23109 23851 23167 23857
rect 23109 23848 23121 23851
rect 23072 23820 23121 23848
rect 23072 23808 23078 23820
rect 23109 23817 23121 23820
rect 23155 23848 23167 23851
rect 23382 23848 23388 23860
rect 23155 23820 23388 23848
rect 23155 23817 23167 23820
rect 23109 23811 23167 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 24670 23808 24676 23860
rect 24728 23848 24734 23860
rect 24765 23851 24823 23857
rect 24765 23848 24777 23851
rect 24728 23820 24777 23848
rect 24728 23808 24734 23820
rect 24765 23817 24777 23820
rect 24811 23817 24823 23851
rect 24765 23811 24823 23817
rect 17770 23740 17776 23792
rect 17828 23780 17834 23792
rect 17828 23752 19288 23780
rect 17828 23740 17834 23752
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23712 13139 23715
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 13127 23684 13461 23712
rect 13127 23681 13139 23684
rect 13081 23675 13139 23681
rect 13449 23681 13461 23684
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 18288 23684 19196 23712
rect 18288 23672 18294 23684
rect 19168 23656 19196 23684
rect 12158 23644 12164 23656
rect 11348 23616 11560 23644
rect 12119 23616 12164 23644
rect 9769 23579 9827 23585
rect 9769 23545 9781 23579
rect 9815 23576 9827 23579
rect 10689 23579 10747 23585
rect 10689 23576 10701 23579
rect 9815 23548 10701 23576
rect 9815 23545 9827 23548
rect 9769 23539 9827 23545
rect 10689 23545 10701 23548
rect 10735 23576 10747 23579
rect 11149 23579 11207 23585
rect 11149 23576 11161 23579
rect 10735 23548 11161 23576
rect 10735 23545 10747 23548
rect 10689 23539 10747 23545
rect 11149 23545 11161 23548
rect 11195 23545 11207 23579
rect 11149 23539 11207 23545
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 11348 23517 11376 23616
rect 12158 23604 12164 23616
rect 12216 23644 12222 23656
rect 14185 23647 14243 23653
rect 14185 23644 14197 23647
rect 12216 23616 13032 23644
rect 12216 23604 12222 23616
rect 13004 23585 13032 23616
rect 14016 23616 14197 23644
rect 12989 23579 13047 23585
rect 12989 23545 13001 23579
rect 13035 23545 13047 23579
rect 12989 23539 13047 23545
rect 11333 23511 11391 23517
rect 11333 23508 11345 23511
rect 10836 23480 11345 23508
rect 10836 23468 10842 23480
rect 11333 23477 11345 23480
rect 11379 23477 11391 23511
rect 11333 23471 11391 23477
rect 11422 23468 11428 23520
rect 11480 23508 11486 23520
rect 11793 23511 11851 23517
rect 11793 23508 11805 23511
rect 11480 23480 11805 23508
rect 11480 23468 11486 23480
rect 11793 23477 11805 23480
rect 11839 23508 11851 23511
rect 12434 23508 12440 23520
rect 11839 23480 12440 23508
rect 11839 23477 11851 23480
rect 11793 23471 11851 23477
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14016 23517 14044 23616
rect 14185 23613 14197 23616
rect 14231 23613 14243 23647
rect 14185 23607 14243 23613
rect 14274 23604 14280 23656
rect 14332 23644 14338 23656
rect 14452 23647 14510 23653
rect 14452 23644 14464 23647
rect 14332 23616 14464 23644
rect 14332 23604 14338 23616
rect 14452 23613 14464 23616
rect 14498 23644 14510 23647
rect 14826 23644 14832 23656
rect 14498 23616 14832 23644
rect 14498 23613 14510 23616
rect 14452 23607 14510 23613
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 16669 23647 16727 23653
rect 16669 23613 16681 23647
rect 16715 23644 16727 23647
rect 18598 23644 18604 23656
rect 16715 23616 17264 23644
rect 18559 23616 18604 23644
rect 16715 23613 16727 23616
rect 16669 23607 16727 23613
rect 17236 23520 17264 23616
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 19150 23604 19156 23656
rect 19208 23604 19214 23656
rect 19260 23653 19288 23752
rect 20530 23740 20536 23792
rect 20588 23780 20594 23792
rect 22756 23780 22784 23808
rect 20588 23752 22784 23780
rect 20588 23740 20594 23752
rect 24670 23672 24676 23724
rect 24728 23712 24734 23724
rect 25222 23712 25228 23724
rect 24728 23684 25228 23712
rect 24728 23672 24734 23684
rect 25222 23672 25228 23684
rect 25280 23712 25286 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 25280 23684 25513 23712
rect 25280 23672 25286 23684
rect 25501 23681 25513 23684
rect 25547 23681 25559 23715
rect 25501 23675 25559 23681
rect 19610 23653 19616 23656
rect 19245 23647 19303 23653
rect 19245 23613 19257 23647
rect 19291 23644 19303 23647
rect 19337 23647 19395 23653
rect 19337 23644 19349 23647
rect 19291 23616 19349 23644
rect 19291 23613 19303 23616
rect 19245 23607 19303 23613
rect 19337 23613 19349 23616
rect 19383 23613 19395 23647
rect 19604 23644 19616 23653
rect 19337 23607 19395 23613
rect 19444 23616 19616 23644
rect 18690 23536 18696 23588
rect 18748 23576 18754 23588
rect 19444 23576 19472 23616
rect 19604 23607 19616 23616
rect 19610 23604 19616 23607
rect 19668 23604 19674 23656
rect 21821 23647 21879 23653
rect 21821 23613 21833 23647
rect 21867 23613 21879 23647
rect 21821 23607 21879 23613
rect 24581 23647 24639 23653
rect 24581 23613 24593 23647
rect 24627 23644 24639 23647
rect 24627 23616 25268 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 18748 23548 19472 23576
rect 21836 23576 21864 23607
rect 22465 23579 22523 23585
rect 22465 23576 22477 23579
rect 21836 23548 22477 23576
rect 18748 23536 18754 23548
rect 22465 23545 22477 23548
rect 22511 23576 22523 23579
rect 23290 23576 23296 23588
rect 22511 23548 23296 23576
rect 22511 23545 22523 23548
rect 22465 23539 22523 23545
rect 23290 23536 23296 23548
rect 23348 23536 23354 23588
rect 25240 23520 25268 23616
rect 14001 23511 14059 23517
rect 14001 23508 14013 23511
rect 13872 23480 14013 23508
rect 13872 23468 13878 23480
rect 14001 23477 14013 23480
rect 14047 23477 14059 23511
rect 14001 23471 14059 23477
rect 14182 23468 14188 23520
rect 14240 23508 14246 23520
rect 14734 23508 14740 23520
rect 14240 23480 14740 23508
rect 14240 23468 14246 23480
rect 14734 23468 14740 23480
rect 14792 23468 14798 23520
rect 15286 23468 15292 23520
rect 15344 23508 15350 23520
rect 15565 23511 15623 23517
rect 15565 23508 15577 23511
rect 15344 23480 15577 23508
rect 15344 23468 15350 23480
rect 15565 23477 15577 23480
rect 15611 23477 15623 23511
rect 15565 23471 15623 23477
rect 15838 23468 15844 23520
rect 15896 23508 15902 23520
rect 16117 23511 16175 23517
rect 16117 23508 16129 23511
rect 15896 23480 16129 23508
rect 15896 23468 15902 23480
rect 16117 23477 16129 23480
rect 16163 23477 16175 23511
rect 17218 23508 17224 23520
rect 17179 23480 17224 23508
rect 16117 23471 16175 23477
rect 17218 23468 17224 23480
rect 17276 23468 17282 23520
rect 18325 23511 18383 23517
rect 18325 23477 18337 23511
rect 18371 23508 18383 23511
rect 19058 23508 19064 23520
rect 18371 23480 19064 23508
rect 18371 23477 18383 23480
rect 18325 23471 18383 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 20714 23508 20720 23520
rect 20675 23480 20720 23508
rect 20714 23468 20720 23480
rect 20772 23468 20778 23520
rect 21358 23508 21364 23520
rect 21319 23480 21364 23508
rect 21358 23468 21364 23480
rect 21416 23468 21422 23520
rect 25222 23508 25228 23520
rect 25183 23480 25228 23508
rect 25222 23468 25228 23480
rect 25280 23468 25286 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 10962 23264 10968 23316
rect 11020 23264 11026 23316
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 11296 23276 11621 23304
rect 11296 23264 11302 23276
rect 11609 23273 11621 23276
rect 11655 23273 11667 23307
rect 11609 23267 11667 23273
rect 14093 23307 14151 23313
rect 14093 23273 14105 23307
rect 14139 23304 14151 23307
rect 14274 23304 14280 23316
rect 14139 23276 14280 23304
rect 14139 23273 14151 23276
rect 14093 23267 14151 23273
rect 14274 23264 14280 23276
rect 14332 23264 14338 23316
rect 18690 23304 18696 23316
rect 18651 23276 18696 23304
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 20346 23304 20352 23316
rect 19812 23276 20352 23304
rect 10980 23236 11008 23264
rect 11422 23236 11428 23248
rect 10244 23208 11428 23236
rect 10134 23060 10140 23112
rect 10192 23100 10198 23112
rect 10244 23109 10272 23208
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 12526 23196 12532 23248
rect 12584 23236 12590 23248
rect 12958 23239 13016 23245
rect 12958 23236 12970 23239
rect 12584 23208 12970 23236
rect 12584 23196 12590 23208
rect 12958 23205 12970 23208
rect 13004 23236 13016 23239
rect 13078 23236 13084 23248
rect 13004 23208 13084 23236
rect 13004 23205 13016 23208
rect 12958 23199 13016 23205
rect 13078 23196 13084 23208
rect 13136 23196 13142 23248
rect 17770 23236 17776 23248
rect 16684 23208 17776 23236
rect 10496 23171 10554 23177
rect 10496 23137 10508 23171
rect 10542 23168 10554 23171
rect 10962 23168 10968 23180
rect 10542 23140 10968 23168
rect 10542 23137 10554 23140
rect 10496 23131 10554 23137
rect 10962 23128 10968 23140
rect 11020 23128 11026 23180
rect 13722 23168 13728 23180
rect 12728 23140 13728 23168
rect 10229 23103 10287 23109
rect 10229 23100 10241 23103
rect 10192 23072 10241 23100
rect 10192 23060 10198 23072
rect 10229 23069 10241 23072
rect 10275 23069 10287 23103
rect 10229 23063 10287 23069
rect 12434 23060 12440 23112
rect 12492 23100 12498 23112
rect 12728 23109 12756 23140
rect 13722 23128 13728 23140
rect 13780 23128 13786 23180
rect 16684 23177 16712 23208
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 18966 23196 18972 23248
rect 19024 23236 19030 23248
rect 19812 23245 19840 23276
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 21085 23307 21143 23313
rect 21085 23273 21097 23307
rect 21131 23304 21143 23307
rect 22002 23304 22008 23316
rect 21131 23276 22008 23304
rect 21131 23273 21143 23276
rect 21085 23267 21143 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 23474 23264 23480 23316
rect 23532 23304 23538 23316
rect 24765 23307 24823 23313
rect 24765 23304 24777 23307
rect 23532 23276 24777 23304
rect 23532 23264 23538 23276
rect 24765 23273 24777 23276
rect 24811 23273 24823 23307
rect 24765 23267 24823 23273
rect 19797 23239 19855 23245
rect 19797 23236 19809 23239
rect 19024 23208 19809 23236
rect 19024 23196 19030 23208
rect 19797 23205 19809 23208
rect 19843 23205 19855 23239
rect 19797 23199 19855 23205
rect 19886 23196 19892 23248
rect 19944 23236 19950 23248
rect 20070 23236 20076 23248
rect 19944 23208 20076 23236
rect 19944 23196 19950 23208
rect 20070 23196 20076 23208
rect 20128 23236 20134 23248
rect 20622 23236 20628 23248
rect 20128 23208 20628 23236
rect 20128 23196 20134 23208
rect 20622 23196 20628 23208
rect 20680 23196 20686 23248
rect 22922 23196 22928 23248
rect 22980 23236 22986 23248
rect 23017 23239 23075 23245
rect 23017 23236 23029 23239
rect 22980 23208 23029 23236
rect 22980 23196 22986 23208
rect 23017 23205 23029 23208
rect 23063 23236 23075 23239
rect 23566 23236 23572 23248
rect 23063 23208 23572 23236
rect 23063 23205 23075 23208
rect 23017 23199 23075 23205
rect 23566 23196 23572 23208
rect 23624 23196 23630 23248
rect 16942 23177 16948 23180
rect 16669 23171 16727 23177
rect 16669 23137 16681 23171
rect 16715 23137 16727 23171
rect 16936 23168 16948 23177
rect 16903 23140 16948 23168
rect 16669 23131 16727 23137
rect 16936 23131 16948 23140
rect 16942 23128 16948 23131
rect 17000 23128 17006 23180
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 19576 23140 19625 23168
rect 19576 23128 19582 23140
rect 19613 23137 19625 23140
rect 19659 23137 19671 23171
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 19613 23131 19671 23137
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22830 23168 22836 23180
rect 22791 23140 22836 23168
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 24581 23171 24639 23177
rect 24581 23168 24593 23171
rect 23900 23140 24593 23168
rect 23900 23128 23906 23140
rect 24581 23137 24593 23140
rect 24627 23137 24639 23171
rect 24581 23131 24639 23137
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12492 23072 12725 23100
rect 12492 23060 12498 23072
rect 12713 23069 12725 23072
rect 12759 23069 12771 23103
rect 12713 23063 12771 23069
rect 14734 23060 14740 23112
rect 14792 23100 14798 23112
rect 15289 23103 15347 23109
rect 15289 23100 15301 23103
rect 14792 23072 15301 23100
rect 14792 23060 14798 23072
rect 15289 23069 15301 23072
rect 15335 23069 15347 23103
rect 15289 23063 15347 23069
rect 22278 23060 22284 23112
rect 22336 23100 22342 23112
rect 22373 23103 22431 23109
rect 22373 23100 22385 23103
rect 22336 23072 22385 23100
rect 22336 23060 22342 23072
rect 22373 23069 22385 23072
rect 22419 23100 22431 23103
rect 23106 23100 23112 23112
rect 22419 23072 23112 23100
rect 22419 23069 22431 23072
rect 22373 23063 22431 23069
rect 23106 23060 23112 23072
rect 23164 23060 23170 23112
rect 12529 22967 12587 22973
rect 12529 22933 12541 22967
rect 12575 22964 12587 22967
rect 12986 22964 12992 22976
rect 12575 22936 12992 22964
rect 12575 22933 12587 22936
rect 12529 22927 12587 22933
rect 12986 22924 12992 22936
rect 13044 22964 13050 22976
rect 13722 22964 13728 22976
rect 13044 22936 13728 22964
rect 13044 22924 13050 22936
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 16485 22967 16543 22973
rect 16485 22933 16497 22967
rect 16531 22964 16543 22967
rect 17310 22964 17316 22976
rect 16531 22936 17316 22964
rect 16531 22933 16543 22936
rect 16485 22927 16543 22933
rect 17310 22924 17316 22936
rect 17368 22964 17374 22976
rect 18049 22967 18107 22973
rect 18049 22964 18061 22967
rect 17368 22936 18061 22964
rect 17368 22924 17374 22936
rect 18049 22933 18061 22936
rect 18095 22933 18107 22967
rect 19334 22964 19340 22976
rect 19295 22936 19340 22964
rect 18049 22927 18107 22933
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 22554 22964 22560 22976
rect 22515 22936 22560 22964
rect 22554 22924 22560 22936
rect 22612 22924 22618 22976
rect 23753 22967 23811 22973
rect 23753 22933 23765 22967
rect 23799 22964 23811 22967
rect 23934 22964 23940 22976
rect 23799 22936 23940 22964
rect 23799 22933 23811 22936
rect 23753 22927 23811 22933
rect 23934 22924 23940 22936
rect 23992 22924 23998 22976
rect 24118 22964 24124 22976
rect 24079 22936 24124 22964
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 10962 22760 10968 22772
rect 10923 22732 10968 22760
rect 10962 22720 10968 22732
rect 11020 22720 11026 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12713 22763 12771 22769
rect 12713 22760 12725 22763
rect 12492 22732 12725 22760
rect 12492 22720 12498 22732
rect 12713 22729 12725 22732
rect 12759 22729 12771 22763
rect 13078 22760 13084 22772
rect 13039 22732 13084 22760
rect 12713 22723 12771 22729
rect 13078 22720 13084 22732
rect 13136 22720 13142 22772
rect 15933 22763 15991 22769
rect 15933 22729 15945 22763
rect 15979 22760 15991 22763
rect 16942 22760 16948 22772
rect 15979 22732 16948 22760
rect 15979 22729 15991 22732
rect 15933 22723 15991 22729
rect 16942 22720 16948 22732
rect 17000 22760 17006 22772
rect 17954 22760 17960 22772
rect 17000 22732 17960 22760
rect 17000 22720 17006 22732
rect 17954 22720 17960 22732
rect 18012 22720 18018 22772
rect 18693 22763 18751 22769
rect 18693 22729 18705 22763
rect 18739 22760 18751 22763
rect 19886 22760 19892 22772
rect 18739 22732 19892 22760
rect 18739 22729 18751 22732
rect 18693 22723 18751 22729
rect 19886 22720 19892 22732
rect 19944 22720 19950 22772
rect 21545 22763 21603 22769
rect 21545 22729 21557 22763
rect 21591 22760 21603 22763
rect 22278 22760 22284 22772
rect 21591 22732 22284 22760
rect 21591 22729 21603 22732
rect 21545 22723 21603 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 22922 22720 22928 22772
rect 22980 22760 22986 22772
rect 23017 22763 23075 22769
rect 23017 22760 23029 22763
rect 22980 22732 23029 22760
rect 22980 22720 22986 22732
rect 23017 22729 23029 22732
rect 23063 22729 23075 22763
rect 23474 22760 23480 22772
rect 23435 22732 23480 22760
rect 23017 22723 23075 22729
rect 23474 22720 23480 22732
rect 23532 22720 23538 22772
rect 25409 22763 25467 22769
rect 23584 22732 24348 22760
rect 14277 22695 14335 22701
rect 14277 22661 14289 22695
rect 14323 22692 14335 22695
rect 14550 22692 14556 22704
rect 14323 22664 14556 22692
rect 14323 22661 14335 22664
rect 14277 22655 14335 22661
rect 14550 22652 14556 22664
rect 14608 22652 14614 22704
rect 16485 22695 16543 22701
rect 16485 22661 16497 22695
rect 16531 22692 16543 22695
rect 16574 22692 16580 22704
rect 16531 22664 16580 22692
rect 16531 22661 16543 22664
rect 16485 22655 16543 22661
rect 16574 22652 16580 22664
rect 16632 22652 16638 22704
rect 17494 22692 17500 22704
rect 17407 22664 17500 22692
rect 17494 22652 17500 22664
rect 17552 22692 17558 22704
rect 17770 22692 17776 22704
rect 17552 22664 17776 22692
rect 17552 22652 17558 22664
rect 17770 22652 17776 22664
rect 17828 22652 17834 22704
rect 22094 22652 22100 22704
rect 22152 22692 22158 22704
rect 22152 22664 22197 22692
rect 22152 22652 22158 22664
rect 23382 22652 23388 22704
rect 23440 22692 23446 22704
rect 23584 22692 23612 22732
rect 23750 22692 23756 22704
rect 23440 22664 23612 22692
rect 23711 22664 23756 22692
rect 23440 22652 23446 22664
rect 23750 22652 23756 22664
rect 23808 22652 23814 22704
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22624 14151 22627
rect 14734 22624 14740 22636
rect 14139 22596 14740 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 14734 22584 14740 22596
rect 14792 22584 14798 22636
rect 14829 22627 14887 22633
rect 14829 22593 14841 22627
rect 14875 22624 14887 22627
rect 15102 22624 15108 22636
rect 14875 22596 15108 22624
rect 14875 22593 14887 22596
rect 14829 22587 14887 22593
rect 13725 22559 13783 22565
rect 13725 22525 13737 22559
rect 13771 22556 13783 22559
rect 14642 22556 14648 22568
rect 13771 22528 14648 22556
rect 13771 22525 13783 22528
rect 13725 22519 13783 22525
rect 14642 22516 14648 22528
rect 14700 22556 14706 22568
rect 14844 22556 14872 22587
rect 15102 22584 15108 22596
rect 15160 22584 15166 22636
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 21818 22584 21824 22596
rect 21876 22624 21882 22636
rect 21876 22596 22600 22624
rect 21876 22584 21882 22596
rect 14700 22528 14872 22556
rect 16761 22559 16819 22565
rect 14700 22516 14706 22528
rect 16761 22525 16773 22559
rect 16807 22556 16819 22559
rect 16850 22556 16856 22568
rect 16807 22528 16856 22556
rect 16807 22525 16819 22528
rect 16761 22519 16819 22525
rect 16850 22516 16856 22528
rect 16908 22556 16914 22568
rect 19429 22559 19487 22565
rect 16908 22528 17908 22556
rect 16908 22516 16914 22528
rect 14458 22448 14464 22500
rect 14516 22488 14522 22500
rect 14737 22491 14795 22497
rect 14737 22488 14749 22491
rect 14516 22460 14749 22488
rect 14516 22448 14522 22460
rect 14737 22457 14749 22460
rect 14783 22457 14795 22491
rect 14737 22451 14795 22457
rect 16114 22448 16120 22500
rect 16172 22488 16178 22500
rect 16209 22491 16267 22497
rect 16209 22488 16221 22491
rect 16172 22460 16221 22488
rect 16172 22448 16178 22460
rect 16209 22457 16221 22460
rect 16255 22457 16267 22491
rect 16209 22451 16267 22457
rect 17037 22491 17095 22497
rect 17037 22457 17049 22491
rect 17083 22488 17095 22491
rect 17310 22488 17316 22500
rect 17083 22460 17316 22488
rect 17083 22457 17095 22460
rect 17037 22451 17095 22457
rect 10134 22380 10140 22432
rect 10192 22420 10198 22432
rect 10229 22423 10287 22429
rect 10229 22420 10241 22423
rect 10192 22392 10241 22420
rect 10192 22380 10198 22392
rect 10229 22389 10241 22392
rect 10275 22389 10287 22423
rect 10229 22383 10287 22389
rect 10505 22423 10563 22429
rect 10505 22389 10517 22423
rect 10551 22420 10563 22423
rect 10686 22420 10692 22432
rect 10551 22392 10692 22420
rect 10551 22389 10563 22392
rect 10505 22383 10563 22389
rect 10686 22380 10692 22392
rect 10744 22380 10750 22432
rect 16224 22420 16252 22451
rect 17310 22448 17316 22460
rect 17368 22448 17374 22500
rect 17880 22488 17908 22528
rect 19429 22525 19441 22559
rect 19475 22556 19487 22559
rect 19521 22559 19579 22565
rect 19521 22556 19533 22559
rect 19475 22528 19533 22556
rect 19475 22525 19487 22528
rect 19429 22519 19487 22525
rect 19521 22525 19533 22528
rect 19567 22556 19579 22559
rect 20530 22556 20536 22568
rect 19567 22528 20536 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 19788 22491 19846 22497
rect 17880 22460 19104 22488
rect 16945 22423 17003 22429
rect 16945 22420 16957 22423
rect 16224 22392 16957 22420
rect 16945 22389 16957 22392
rect 16991 22389 17003 22423
rect 18966 22420 18972 22432
rect 18927 22392 18972 22420
rect 16945 22383 17003 22389
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 19076 22420 19104 22460
rect 19788 22457 19800 22491
rect 19834 22488 19846 22491
rect 19886 22488 19892 22500
rect 19834 22460 19892 22488
rect 19834 22457 19846 22460
rect 19788 22451 19846 22457
rect 19886 22448 19892 22460
rect 19944 22448 19950 22500
rect 22373 22491 22431 22497
rect 22373 22488 22385 22491
rect 19996 22460 22385 22488
rect 19996 22420 20024 22460
rect 22373 22457 22385 22460
rect 22419 22488 22431 22491
rect 22462 22488 22468 22500
rect 22419 22460 22468 22488
rect 22419 22457 22431 22460
rect 22373 22451 22431 22457
rect 22462 22448 22468 22460
rect 22520 22448 22526 22500
rect 22572 22497 22600 22596
rect 23566 22584 23572 22636
rect 23624 22624 23630 22636
rect 24118 22624 24124 22636
rect 23624 22596 24124 22624
rect 23624 22584 23630 22596
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24320 22633 24348 22732
rect 25409 22729 25421 22763
rect 25455 22760 25467 22763
rect 25590 22760 25596 22772
rect 25455 22732 25596 22760
rect 25455 22729 25467 22732
rect 25409 22723 25467 22729
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22624 24363 22627
rect 24486 22624 24492 22636
rect 24351 22596 24492 22624
rect 24351 22593 24363 22596
rect 24305 22587 24363 22593
rect 24486 22584 24492 22596
rect 24544 22584 24550 22636
rect 23842 22516 23848 22568
rect 23900 22556 23906 22568
rect 24673 22559 24731 22565
rect 24673 22556 24685 22559
rect 23900 22528 24685 22556
rect 23900 22516 23906 22528
rect 24673 22525 24685 22528
rect 24719 22525 24731 22559
rect 24673 22519 24731 22525
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22525 25283 22559
rect 25225 22519 25283 22525
rect 22557 22491 22615 22497
rect 22557 22457 22569 22491
rect 22603 22457 22615 22491
rect 22557 22451 22615 22457
rect 22649 22491 22707 22497
rect 22649 22457 22661 22491
rect 22695 22488 22707 22491
rect 23106 22488 23112 22500
rect 22695 22460 23112 22488
rect 22695 22457 22707 22460
rect 22649 22451 22707 22457
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 23934 22448 23940 22500
rect 23992 22448 23998 22500
rect 25240 22488 25268 22519
rect 25866 22488 25872 22500
rect 25240 22460 25872 22488
rect 25866 22448 25872 22460
rect 25924 22448 25930 22500
rect 19076 22392 20024 22420
rect 20622 22380 20628 22432
rect 20680 22420 20686 22432
rect 20901 22423 20959 22429
rect 20901 22420 20913 22423
rect 20680 22392 20913 22420
rect 20680 22380 20686 22392
rect 20901 22389 20913 22392
rect 20947 22389 20959 22423
rect 20901 22383 20959 22389
rect 23474 22380 23480 22432
rect 23532 22420 23538 22432
rect 23952 22420 23980 22448
rect 24213 22423 24271 22429
rect 24213 22420 24225 22423
rect 23532 22392 24225 22420
rect 23532 22380 23538 22392
rect 24213 22389 24225 22392
rect 24259 22389 24271 22423
rect 24213 22383 24271 22389
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10965 22219 11023 22225
rect 10965 22216 10977 22219
rect 10008 22188 10977 22216
rect 10008 22176 10014 22188
rect 10965 22185 10977 22188
rect 11011 22185 11023 22219
rect 10965 22179 11023 22185
rect 14458 22176 14464 22228
rect 14516 22216 14522 22228
rect 14645 22219 14703 22225
rect 14645 22216 14657 22219
rect 14516 22188 14657 22216
rect 14516 22176 14522 22188
rect 14645 22185 14657 22188
rect 14691 22185 14703 22219
rect 14645 22179 14703 22185
rect 17221 22219 17279 22225
rect 17221 22185 17233 22219
rect 17267 22216 17279 22219
rect 17402 22216 17408 22228
rect 17267 22188 17408 22216
rect 17267 22185 17279 22188
rect 17221 22179 17279 22185
rect 17402 22176 17408 22188
rect 17460 22176 17466 22228
rect 19337 22219 19395 22225
rect 19337 22185 19349 22219
rect 19383 22216 19395 22219
rect 19518 22216 19524 22228
rect 19383 22188 19524 22216
rect 19383 22185 19395 22188
rect 19337 22179 19395 22185
rect 19518 22176 19524 22188
rect 19576 22216 19582 22228
rect 19797 22219 19855 22225
rect 19797 22216 19809 22219
rect 19576 22188 19809 22216
rect 19576 22176 19582 22188
rect 19797 22185 19809 22188
rect 19843 22185 19855 22219
rect 19797 22179 19855 22185
rect 20898 22176 20904 22228
rect 20956 22216 20962 22228
rect 21085 22219 21143 22225
rect 21085 22216 21097 22219
rect 20956 22188 21097 22216
rect 20956 22176 20962 22188
rect 21085 22185 21097 22188
rect 21131 22185 21143 22219
rect 21085 22179 21143 22185
rect 23014 22176 23020 22228
rect 23072 22216 23078 22228
rect 23072 22188 23336 22216
rect 23072 22176 23078 22188
rect 23308 22160 23336 22188
rect 23658 22176 23664 22228
rect 23716 22216 23722 22228
rect 23753 22219 23811 22225
rect 23753 22216 23765 22219
rect 23716 22188 23765 22216
rect 23716 22176 23722 22188
rect 23753 22185 23765 22188
rect 23799 22216 23811 22219
rect 24486 22216 24492 22228
rect 23799 22188 24492 22216
rect 23799 22185 23811 22188
rect 23753 22179 23811 22185
rect 24486 22176 24492 22188
rect 24544 22176 24550 22228
rect 14185 22151 14243 22157
rect 14185 22148 14197 22151
rect 13740 22120 14197 22148
rect 13630 22040 13636 22092
rect 13688 22080 13694 22092
rect 13740 22080 13768 22120
rect 14185 22117 14197 22120
rect 14231 22117 14243 22151
rect 16850 22148 16856 22160
rect 14185 22111 14243 22117
rect 16592 22120 16856 22148
rect 13688 22052 13768 22080
rect 16485 22083 16543 22089
rect 13688 22040 13694 22052
rect 16485 22049 16497 22083
rect 16531 22080 16543 22083
rect 16592 22080 16620 22120
rect 16850 22108 16856 22120
rect 16908 22108 16914 22160
rect 18785 22151 18843 22157
rect 18785 22148 18797 22151
rect 17880 22120 18797 22148
rect 17034 22080 17040 22092
rect 16531 22052 16620 22080
rect 16995 22052 17040 22080
rect 16531 22049 16543 22052
rect 16485 22043 16543 22049
rect 17034 22040 17040 22052
rect 17092 22040 17098 22092
rect 17770 22040 17776 22092
rect 17828 22080 17834 22092
rect 17880 22080 17908 22120
rect 18785 22117 18797 22120
rect 18831 22117 18843 22151
rect 18785 22111 18843 22117
rect 19705 22151 19763 22157
rect 19705 22117 19717 22151
rect 19751 22148 19763 22151
rect 19978 22148 19984 22160
rect 19751 22120 19984 22148
rect 19751 22117 19763 22120
rect 19705 22111 19763 22117
rect 19978 22108 19984 22120
rect 20036 22108 20042 22160
rect 22094 22108 22100 22160
rect 22152 22148 22158 22160
rect 22925 22151 22983 22157
rect 22925 22148 22937 22151
rect 22152 22120 22937 22148
rect 22152 22108 22158 22120
rect 22925 22117 22937 22120
rect 22971 22117 22983 22151
rect 22925 22111 22983 22117
rect 23290 22108 23296 22160
rect 23348 22108 23354 22160
rect 23952 22120 24164 22148
rect 17828 22052 17908 22080
rect 17828 22040 17834 22052
rect 22462 22040 22468 22092
rect 22520 22040 22526 22092
rect 22554 22040 22560 22092
rect 22612 22080 22618 22092
rect 22741 22083 22799 22089
rect 22741 22080 22753 22083
rect 22612 22052 22753 22080
rect 22612 22040 22618 22052
rect 22741 22049 22753 22052
rect 22787 22049 22799 22083
rect 23014 22080 23020 22092
rect 22927 22052 23020 22080
rect 22741 22043 22799 22049
rect 23014 22040 23020 22052
rect 23072 22080 23078 22092
rect 23952 22080 23980 22120
rect 23072 22052 23980 22080
rect 24136 22080 24164 22120
rect 24210 22089 24216 22092
rect 24193 22083 24216 22089
rect 24193 22080 24205 22083
rect 24136 22052 24205 22080
rect 23072 22040 23078 22052
rect 24193 22049 24205 22052
rect 24268 22080 24274 22092
rect 24268 22052 24341 22080
rect 24193 22043 24216 22049
rect 24210 22040 24216 22043
rect 24268 22040 24274 22052
rect 10870 22012 10876 22024
rect 10831 21984 10876 22012
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 14090 22012 14096 22024
rect 14051 21984 14096 22012
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 14274 22012 14280 22024
rect 14235 21984 14280 22012
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 17310 22012 17316 22024
rect 17271 21984 17316 22012
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 18693 22015 18751 22021
rect 18693 21981 18705 22015
rect 18739 21981 18751 22015
rect 18874 22012 18880 22024
rect 18835 21984 18880 22012
rect 18693 21975 18751 21981
rect 16761 21947 16819 21953
rect 16761 21913 16773 21947
rect 16807 21944 16819 21947
rect 18049 21947 18107 21953
rect 18049 21944 18061 21947
rect 16807 21916 18061 21944
rect 16807 21913 16819 21916
rect 16761 21907 16819 21913
rect 18049 21913 18061 21916
rect 18095 21944 18107 21947
rect 18708 21944 18736 21975
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 22097 22015 22155 22021
rect 22097 21981 22109 22015
rect 22143 22012 22155 22015
rect 22480 22012 22508 22040
rect 22830 22012 22836 22024
rect 22143 21984 22836 22012
rect 22143 21981 22155 21984
rect 22097 21975 22155 21981
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 22922 21972 22928 22024
rect 22980 22012 22986 22024
rect 23937 22015 23995 22021
rect 23937 22012 23949 22015
rect 22980 21984 23949 22012
rect 22980 21972 22986 21984
rect 23937 21981 23949 21984
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 18095 21916 18736 21944
rect 22465 21947 22523 21953
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 22465 21913 22477 21947
rect 22511 21944 22523 21947
rect 23474 21944 23480 21956
rect 22511 21916 23480 21944
rect 22511 21913 22523 21916
rect 22465 21907 22523 21913
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 23658 21904 23664 21956
rect 23716 21944 23722 21956
rect 23716 21916 23980 21944
rect 23716 21904 23722 21916
rect 10505 21879 10563 21885
rect 10505 21845 10517 21879
rect 10551 21876 10563 21879
rect 10870 21876 10876 21888
rect 10551 21848 10876 21876
rect 10551 21845 10563 21848
rect 10505 21839 10563 21845
rect 10870 21836 10876 21848
rect 10928 21836 10934 21888
rect 13722 21876 13728 21888
rect 13683 21848 13728 21876
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 18322 21876 18328 21888
rect 18283 21848 18328 21876
rect 18322 21836 18328 21848
rect 18380 21836 18386 21888
rect 21726 21876 21732 21888
rect 21687 21848 21732 21876
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 23952 21876 23980 21916
rect 25317 21879 25375 21885
rect 25317 21876 25329 21879
rect 23952 21848 25329 21876
rect 25317 21845 25329 21848
rect 25363 21845 25375 21879
rect 25317 21839 25375 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 10778 21672 10784 21684
rect 9907 21644 10784 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 13630 21672 13636 21684
rect 13591 21644 13636 21672
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 15562 21672 15568 21684
rect 14292 21644 15568 21672
rect 14292 21616 14320 21644
rect 15562 21632 15568 21644
rect 15620 21672 15626 21684
rect 15749 21675 15807 21681
rect 15749 21672 15761 21675
rect 15620 21644 15761 21672
rect 15620 21632 15626 21644
rect 15749 21641 15761 21644
rect 15795 21641 15807 21675
rect 15749 21635 15807 21641
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 17770 21672 17776 21684
rect 16632 21644 17776 21672
rect 16632 21632 16638 21644
rect 17770 21632 17776 21644
rect 17828 21632 17834 21684
rect 18601 21675 18659 21681
rect 18601 21641 18613 21675
rect 18647 21672 18659 21675
rect 18874 21672 18880 21684
rect 18647 21644 18880 21672
rect 18647 21641 18659 21644
rect 18601 21635 18659 21641
rect 18874 21632 18880 21644
rect 18932 21632 18938 21684
rect 21545 21675 21603 21681
rect 21545 21641 21557 21675
rect 21591 21672 21603 21675
rect 22002 21672 22008 21684
rect 21591 21644 22008 21672
rect 21591 21641 21603 21644
rect 21545 21635 21603 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 22097 21675 22155 21681
rect 22097 21641 22109 21675
rect 22143 21672 22155 21675
rect 23566 21672 23572 21684
rect 22143 21644 23572 21672
rect 22143 21641 22155 21644
rect 22097 21635 22155 21641
rect 23566 21632 23572 21644
rect 23624 21632 23630 21684
rect 10042 21564 10048 21616
rect 10100 21604 10106 21616
rect 10413 21607 10471 21613
rect 10413 21604 10425 21607
rect 10100 21576 10425 21604
rect 10100 21564 10106 21576
rect 10413 21573 10425 21576
rect 10459 21573 10471 21607
rect 10413 21567 10471 21573
rect 12989 21607 13047 21613
rect 12989 21573 13001 21607
rect 13035 21604 13047 21607
rect 14274 21604 14280 21616
rect 13035 21576 14280 21604
rect 13035 21573 13047 21576
rect 12989 21567 13047 21573
rect 14274 21564 14280 21576
rect 14332 21564 14338 21616
rect 16758 21604 16764 21616
rect 16719 21576 16764 21604
rect 16758 21564 16764 21576
rect 16816 21564 16822 21616
rect 17034 21604 17040 21616
rect 16995 21576 17040 21604
rect 17034 21564 17040 21576
rect 17092 21564 17098 21616
rect 19242 21604 19248 21616
rect 19203 21576 19248 21604
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 23106 21604 23112 21616
rect 23067 21576 23112 21604
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10137 21539 10195 21545
rect 10137 21536 10149 21539
rect 10008 21508 10149 21536
rect 10008 21496 10014 21508
rect 10137 21505 10149 21508
rect 10183 21505 10195 21539
rect 10962 21536 10968 21548
rect 10923 21508 10968 21536
rect 10137 21499 10195 21505
rect 10962 21496 10968 21508
rect 11020 21536 11026 21548
rect 11333 21539 11391 21545
rect 11333 21536 11345 21539
rect 11020 21508 11345 21536
rect 11020 21496 11026 21508
rect 11333 21505 11345 21508
rect 11379 21505 11391 21539
rect 11333 21499 11391 21505
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21536 13415 21539
rect 13814 21536 13820 21548
rect 13403 21508 13820 21536
rect 13403 21505 13415 21508
rect 13357 21499 13415 21505
rect 13814 21496 13820 21508
rect 13872 21536 13878 21548
rect 14090 21536 14096 21548
rect 13872 21508 14096 21536
rect 13872 21496 13878 21508
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18012 21508 19073 21536
rect 18012 21496 18018 21508
rect 19061 21505 19073 21508
rect 19107 21536 19119 21539
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19107 21508 19809 21536
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 19797 21505 19809 21508
rect 19843 21536 19855 21539
rect 20622 21536 20628 21548
rect 19843 21508 20628 21536
rect 19843 21505 19855 21508
rect 19797 21499 19855 21505
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 22462 21496 22468 21548
rect 22520 21536 22526 21548
rect 22649 21539 22707 21545
rect 22649 21536 22661 21539
rect 22520 21508 22661 21536
rect 22520 21496 22526 21508
rect 22649 21505 22661 21508
rect 22695 21536 22707 21539
rect 23014 21536 23020 21548
rect 22695 21508 23020 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 23014 21496 23020 21508
rect 23072 21496 23078 21548
rect 23124 21508 23520 21536
rect 9493 21471 9551 21477
rect 9493 21437 9505 21471
rect 9539 21468 9551 21471
rect 10686 21468 10692 21480
rect 9539 21440 10692 21468
rect 9539 21437 9551 21440
rect 9493 21431 9551 21437
rect 10686 21428 10692 21440
rect 10744 21428 10750 21480
rect 14642 21477 14648 21480
rect 12069 21471 12127 21477
rect 12069 21468 12081 21471
rect 10888 21440 12081 21468
rect 10888 21412 10916 21440
rect 12069 21437 12081 21440
rect 12115 21437 12127 21471
rect 14369 21471 14427 21477
rect 14369 21468 14381 21471
rect 12069 21431 12127 21437
rect 14200 21440 14381 21468
rect 10870 21400 10876 21412
rect 10831 21372 10876 21400
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 11698 21332 11704 21344
rect 11659 21304 11704 21332
rect 11698 21292 11704 21304
rect 11756 21292 11762 21344
rect 13998 21292 14004 21344
rect 14056 21332 14062 21344
rect 14200 21341 14228 21440
rect 14369 21437 14381 21440
rect 14415 21437 14427 21471
rect 14636 21468 14648 21477
rect 14603 21440 14648 21468
rect 14369 21431 14427 21437
rect 14636 21431 14648 21440
rect 14642 21428 14648 21431
rect 14700 21428 14706 21480
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 19521 21471 19579 21477
rect 19521 21468 19533 21471
rect 19392 21440 19533 21468
rect 19392 21428 19398 21440
rect 19521 21437 19533 21440
rect 19567 21468 19579 21471
rect 20165 21471 20223 21477
rect 20165 21468 20177 21471
rect 19567 21440 20177 21468
rect 19567 21437 19579 21440
rect 19521 21431 19579 21437
rect 20165 21437 20177 21440
rect 20211 21437 20223 21471
rect 20165 21431 20223 21437
rect 22922 21428 22928 21480
rect 22980 21468 22986 21480
rect 23124 21468 23152 21508
rect 22980 21440 23152 21468
rect 22980 21428 22986 21440
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 23382 21468 23388 21480
rect 23256 21440 23388 21468
rect 23256 21428 23262 21440
rect 23382 21428 23388 21440
rect 23440 21428 23446 21480
rect 23492 21477 23520 21508
rect 23477 21471 23535 21477
rect 23477 21437 23489 21471
rect 23523 21468 23535 21471
rect 23658 21468 23664 21480
rect 23523 21440 23664 21468
rect 23523 21437 23535 21440
rect 23477 21431 23535 21437
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 19426 21360 19432 21412
rect 19484 21400 19490 21412
rect 19705 21403 19763 21409
rect 19705 21400 19717 21403
rect 19484 21372 19717 21400
rect 19484 21360 19490 21372
rect 19705 21369 19717 21372
rect 19751 21369 19763 21403
rect 19705 21363 19763 21369
rect 20993 21403 21051 21409
rect 20993 21369 21005 21403
rect 21039 21400 21051 21403
rect 21913 21403 21971 21409
rect 21913 21400 21925 21403
rect 21039 21372 21925 21400
rect 21039 21369 21051 21372
rect 20993 21363 21051 21369
rect 21913 21369 21925 21372
rect 21959 21400 21971 21403
rect 22373 21403 22431 21409
rect 22373 21400 22385 21403
rect 21959 21372 22385 21400
rect 21959 21369 21971 21372
rect 21913 21363 21971 21369
rect 22373 21369 22385 21372
rect 22419 21369 22431 21403
rect 22373 21363 22431 21369
rect 23106 21360 23112 21412
rect 23164 21400 23170 21412
rect 23906 21403 23964 21409
rect 23906 21400 23918 21403
rect 23164 21372 23918 21400
rect 23164 21360 23170 21372
rect 23906 21369 23918 21372
rect 23952 21369 23964 21403
rect 23906 21363 23964 21369
rect 14185 21335 14243 21341
rect 14185 21332 14197 21335
rect 14056 21304 14197 21332
rect 14056 21292 14062 21304
rect 14185 21301 14197 21304
rect 14231 21301 14243 21335
rect 14185 21295 14243 21301
rect 17310 21292 17316 21344
rect 17368 21332 17374 21344
rect 17497 21335 17555 21341
rect 17497 21332 17509 21335
rect 17368 21304 17509 21332
rect 17368 21292 17374 21304
rect 17497 21301 17509 21304
rect 17543 21332 17555 21335
rect 17770 21332 17776 21344
rect 17543 21304 17776 21332
rect 17543 21301 17555 21304
rect 17497 21295 17555 21301
rect 17770 21292 17776 21304
rect 17828 21292 17834 21344
rect 17954 21292 17960 21344
rect 18012 21332 18018 21344
rect 18049 21335 18107 21341
rect 18049 21332 18061 21335
rect 18012 21304 18061 21332
rect 18012 21292 18018 21304
rect 18049 21301 18061 21304
rect 18095 21301 18107 21335
rect 18049 21295 18107 21301
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22557 21335 22615 21341
rect 22557 21332 22569 21335
rect 21784 21304 22569 21332
rect 21784 21292 21790 21304
rect 22557 21301 22569 21304
rect 22603 21332 22615 21335
rect 22738 21332 22744 21344
rect 22603 21304 22744 21332
rect 22603 21301 22615 21304
rect 22557 21295 22615 21301
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 25041 21335 25099 21341
rect 25041 21332 25053 21335
rect 24268 21304 25053 21332
rect 24268 21292 24274 21304
rect 25041 21301 25053 21304
rect 25087 21301 25099 21335
rect 25041 21295 25099 21301
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 10962 21088 10968 21140
rect 11020 21128 11026 21140
rect 11793 21131 11851 21137
rect 11793 21128 11805 21131
rect 11020 21100 11805 21128
rect 11020 21088 11026 21100
rect 11793 21097 11805 21100
rect 11839 21097 11851 21131
rect 11793 21091 11851 21097
rect 13630 21088 13636 21140
rect 13688 21128 13694 21140
rect 13906 21128 13912 21140
rect 13688 21100 13912 21128
rect 13688 21088 13694 21100
rect 13906 21088 13912 21100
rect 13964 21128 13970 21140
rect 14001 21131 14059 21137
rect 14001 21128 14013 21131
rect 13964 21100 14013 21128
rect 13964 21088 13970 21100
rect 14001 21097 14013 21100
rect 14047 21097 14059 21131
rect 14001 21091 14059 21097
rect 14553 21131 14611 21137
rect 14553 21097 14565 21131
rect 14599 21128 14611 21131
rect 14642 21128 14648 21140
rect 14599 21100 14648 21128
rect 14599 21097 14611 21100
rect 14553 21091 14611 21097
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 15841 21131 15899 21137
rect 15841 21097 15853 21131
rect 15887 21128 15899 21131
rect 16482 21128 16488 21140
rect 15887 21100 16488 21128
rect 15887 21097 15899 21100
rect 15841 21091 15899 21097
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 18874 21128 18880 21140
rect 18835 21100 18880 21128
rect 18874 21088 18880 21100
rect 18932 21088 18938 21140
rect 19426 21128 19432 21140
rect 19387 21100 19432 21128
rect 19426 21088 19432 21100
rect 19484 21088 19490 21140
rect 20898 21088 20904 21140
rect 20956 21088 20962 21140
rect 21729 21131 21787 21137
rect 21729 21097 21741 21131
rect 21775 21128 21787 21131
rect 22554 21128 22560 21140
rect 21775 21100 22560 21128
rect 21775 21097 21787 21100
rect 21729 21091 21787 21097
rect 22554 21088 22560 21100
rect 22612 21088 22618 21140
rect 23106 21088 23112 21140
rect 23164 21128 23170 21140
rect 23164 21100 23336 21128
rect 23164 21088 23170 21100
rect 10680 21063 10738 21069
rect 10680 21029 10692 21063
rect 10726 21060 10738 21063
rect 10870 21060 10876 21072
rect 10726 21032 10876 21060
rect 10726 21029 10738 21032
rect 10680 21023 10738 21029
rect 10870 21020 10876 21032
rect 10928 21060 10934 21072
rect 11054 21060 11060 21072
rect 10928 21032 11060 21060
rect 10928 21020 10934 21032
rect 11054 21020 11060 21032
rect 11112 21060 11118 21072
rect 11698 21060 11704 21072
rect 11112 21032 11704 21060
rect 11112 21020 11118 21032
rect 11698 21020 11704 21032
rect 11756 21020 11762 21072
rect 13814 21060 13820 21072
rect 13775 21032 13820 21060
rect 13814 21020 13820 21032
rect 13872 21020 13878 21072
rect 20916 21060 20944 21088
rect 21177 21063 21235 21069
rect 21177 21060 21189 21063
rect 20916 21032 21189 21060
rect 21177 21029 21189 21032
rect 21223 21029 21235 21063
rect 21177 21023 21235 21029
rect 22097 21063 22155 21069
rect 22097 21029 22109 21063
rect 22143 21060 22155 21063
rect 22462 21060 22468 21072
rect 22143 21032 22468 21060
rect 22143 21029 22155 21032
rect 22097 21023 22155 21029
rect 22462 21020 22468 21032
rect 22520 21020 22526 21072
rect 23014 21020 23020 21072
rect 23072 21060 23078 21072
rect 23198 21060 23204 21072
rect 23072 21032 23204 21060
rect 23072 21020 23078 21032
rect 23198 21020 23204 21032
rect 23256 21020 23262 21072
rect 23308 21069 23336 21100
rect 24210 21088 24216 21140
rect 24268 21128 24274 21140
rect 24305 21131 24363 21137
rect 24305 21128 24317 21131
rect 24268 21100 24317 21128
rect 24268 21088 24274 21100
rect 24305 21097 24317 21100
rect 24351 21097 24363 21131
rect 24762 21128 24768 21140
rect 24723 21100 24768 21128
rect 24305 21091 24363 21097
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 23293 21063 23351 21069
rect 23293 21029 23305 21063
rect 23339 21029 23351 21063
rect 23293 21023 23351 21029
rect 12989 20995 13047 21001
rect 12989 20961 13001 20995
rect 13035 20992 13047 20995
rect 17494 20992 17500 21004
rect 13035 20964 14136 20992
rect 17455 20964 17500 20992
rect 13035 20961 13047 20964
rect 12989 20955 13047 20961
rect 14108 20936 14136 20964
rect 17494 20952 17500 20964
rect 17552 20952 17558 21004
rect 17770 21001 17776 21004
rect 17764 20992 17776 21001
rect 17731 20964 17776 20992
rect 17764 20955 17776 20964
rect 17770 20952 17776 20955
rect 17828 20952 17834 21004
rect 20898 20992 20904 21004
rect 20859 20964 20904 20992
rect 20898 20952 20904 20964
rect 20956 20952 20962 21004
rect 24581 20995 24639 21001
rect 24581 20961 24593 20995
rect 24627 20992 24639 20995
rect 25038 20992 25044 21004
rect 24627 20964 25044 20992
rect 24627 20961 24639 20964
rect 24581 20955 24639 20961
rect 25038 20952 25044 20964
rect 25096 20952 25102 21004
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10410 20924 10416 20936
rect 10192 20896 10416 20924
rect 10192 20884 10198 20896
rect 10410 20884 10416 20896
rect 10468 20884 10474 20936
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 16482 20924 16488 20936
rect 16443 20896 16488 20924
rect 16482 20884 16488 20896
rect 16540 20884 16546 20936
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 16632 20896 16677 20924
rect 16632 20884 16638 20896
rect 22646 20884 22652 20936
rect 22704 20924 22710 20936
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 22704 20896 23121 20924
rect 22704 20884 22710 20896
rect 23109 20893 23121 20896
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 13357 20859 13415 20865
rect 13357 20825 13369 20859
rect 13403 20856 13415 20859
rect 13722 20856 13728 20868
rect 13403 20828 13728 20856
rect 13403 20825 13415 20828
rect 13357 20819 13415 20825
rect 13722 20816 13728 20828
rect 13780 20816 13786 20868
rect 22738 20856 22744 20868
rect 22699 20828 22744 20856
rect 22738 20816 22744 20828
rect 22796 20816 22802 20868
rect 13538 20788 13544 20800
rect 13499 20760 13544 20788
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 16022 20788 16028 20800
rect 15983 20760 16028 20788
rect 16022 20748 16028 20760
rect 16080 20748 16086 20800
rect 16942 20788 16948 20800
rect 16903 20760 16948 20788
rect 16942 20748 16948 20760
rect 17000 20748 17006 20800
rect 20625 20791 20683 20797
rect 20625 20757 20637 20791
rect 20671 20788 20683 20791
rect 20714 20788 20720 20800
rect 20671 20760 20720 20788
rect 20671 20757 20683 20760
rect 20625 20751 20683 20757
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 23658 20748 23664 20800
rect 23716 20788 23722 20800
rect 23937 20791 23995 20797
rect 23937 20788 23949 20791
rect 23716 20760 23949 20788
rect 23716 20748 23722 20760
rect 23937 20757 23949 20760
rect 23983 20757 23995 20791
rect 23937 20751 23995 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13630 20584 13636 20596
rect 13035 20556 13636 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14829 20587 14887 20593
rect 14829 20584 14841 20587
rect 14148 20556 14841 20584
rect 14148 20544 14154 20556
rect 14829 20553 14841 20556
rect 14875 20553 14887 20587
rect 14829 20547 14887 20553
rect 15933 20587 15991 20593
rect 15933 20553 15945 20587
rect 15979 20584 15991 20587
rect 16574 20584 16580 20596
rect 15979 20556 16580 20584
rect 15979 20553 15991 20556
rect 15933 20547 15991 20553
rect 16574 20544 16580 20556
rect 16632 20544 16638 20596
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 17494 20544 17500 20556
rect 17552 20584 17558 20596
rect 17773 20587 17831 20593
rect 17773 20584 17785 20587
rect 17552 20556 17785 20584
rect 17552 20544 17558 20556
rect 17773 20553 17785 20556
rect 17819 20553 17831 20587
rect 17773 20547 17831 20553
rect 20625 20587 20683 20593
rect 20625 20553 20637 20587
rect 20671 20584 20683 20587
rect 20898 20584 20904 20596
rect 20671 20556 20904 20584
rect 20671 20553 20683 20556
rect 20625 20547 20683 20553
rect 16482 20516 16488 20528
rect 16443 20488 16488 20516
rect 16482 20476 16488 20488
rect 16540 20476 16546 20528
rect 17788 20516 17816 20547
rect 20898 20544 20904 20556
rect 20956 20584 20962 20596
rect 21545 20587 21603 20593
rect 21545 20584 21557 20587
rect 20956 20556 21557 20584
rect 20956 20544 20962 20556
rect 21545 20553 21557 20556
rect 21591 20553 21603 20587
rect 21545 20547 21603 20553
rect 23106 20544 23112 20596
rect 23164 20584 23170 20596
rect 23385 20587 23443 20593
rect 23385 20584 23397 20587
rect 23164 20556 23397 20584
rect 23164 20544 23170 20556
rect 23385 20553 23397 20556
rect 23431 20553 23443 20587
rect 25038 20584 25044 20596
rect 24999 20556 25044 20584
rect 23385 20547 23443 20553
rect 25038 20544 25044 20556
rect 25096 20544 25102 20596
rect 17788 20488 18092 20516
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20448 16359 20451
rect 16945 20451 17003 20457
rect 16945 20448 16957 20451
rect 16347 20420 16957 20448
rect 16347 20417 16359 20420
rect 16301 20411 16359 20417
rect 16945 20417 16957 20420
rect 16991 20448 17003 20451
rect 17954 20448 17960 20460
rect 16991 20420 17960 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 18064 20457 18092 20488
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 13722 20389 13728 20392
rect 13449 20383 13507 20389
rect 13449 20380 13461 20383
rect 13280 20352 13461 20380
rect 10410 20272 10416 20324
rect 10468 20312 10474 20324
rect 10505 20315 10563 20321
rect 10505 20312 10517 20315
rect 10468 20284 10517 20312
rect 10468 20272 10474 20284
rect 10505 20281 10517 20284
rect 10551 20312 10563 20315
rect 10778 20312 10784 20324
rect 10551 20284 10784 20312
rect 10551 20281 10563 20284
rect 10505 20275 10563 20281
rect 10778 20272 10784 20284
rect 10836 20272 10842 20324
rect 10870 20244 10876 20256
rect 10831 20216 10876 20244
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 12802 20204 12808 20256
rect 12860 20244 12866 20256
rect 13280 20253 13308 20352
rect 13449 20349 13461 20352
rect 13495 20349 13507 20383
rect 13716 20380 13728 20389
rect 13683 20352 13728 20380
rect 13449 20343 13507 20349
rect 13716 20343 13728 20352
rect 13722 20340 13728 20343
rect 13780 20340 13786 20392
rect 15565 20383 15623 20389
rect 15565 20349 15577 20383
rect 15611 20380 15623 20383
rect 18316 20383 18374 20389
rect 18316 20380 18328 20383
rect 15611 20352 17080 20380
rect 15611 20349 15623 20352
rect 15565 20343 15623 20349
rect 16942 20312 16948 20324
rect 16903 20284 16948 20312
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 17052 20321 17080 20352
rect 18156 20352 18328 20380
rect 17037 20315 17095 20321
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 18156 20312 18184 20352
rect 18316 20349 18328 20352
rect 18362 20380 18374 20383
rect 18874 20380 18880 20392
rect 18362 20352 18880 20380
rect 18362 20349 18374 20352
rect 18316 20343 18374 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 20438 20312 20444 20324
rect 17083 20284 18184 20312
rect 20351 20284 20444 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 20438 20272 20444 20284
rect 20496 20312 20502 20324
rect 20901 20315 20959 20321
rect 20901 20312 20913 20315
rect 20496 20284 20913 20312
rect 20496 20272 20502 20284
rect 20901 20281 20913 20284
rect 20947 20281 20959 20315
rect 21174 20312 21180 20324
rect 21135 20284 21180 20312
rect 20901 20275 20959 20281
rect 21174 20272 21180 20284
rect 21232 20272 21238 20324
rect 24305 20315 24363 20321
rect 24305 20281 24317 20315
rect 24351 20312 24363 20315
rect 25130 20312 25136 20324
rect 24351 20284 25136 20312
rect 24351 20281 24363 20284
rect 24305 20275 24363 20281
rect 25130 20272 25136 20284
rect 25188 20272 25194 20324
rect 13265 20247 13323 20253
rect 13265 20244 13277 20247
rect 12860 20216 13277 20244
rect 12860 20204 12866 20216
rect 13265 20213 13277 20216
rect 13311 20213 13323 20247
rect 19426 20244 19432 20256
rect 19387 20216 19432 20244
rect 13265 20207 13323 20213
rect 19426 20204 19432 20216
rect 19484 20204 19490 20256
rect 20714 20204 20720 20256
rect 20772 20244 20778 20256
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 20772 20216 21097 20244
rect 20772 20204 20778 20216
rect 21085 20213 21097 20216
rect 21131 20213 21143 20247
rect 22738 20244 22744 20256
rect 22699 20216 22744 20244
rect 21085 20207 21143 20213
rect 22738 20204 22744 20216
rect 22796 20204 22802 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 24489 20247 24547 20253
rect 24489 20213 24501 20247
rect 24535 20244 24547 20247
rect 24762 20244 24768 20256
rect 24535 20216 24768 20244
rect 24535 20213 24547 20216
rect 24489 20207 24547 20213
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 10870 20000 10876 20052
rect 10928 20040 10934 20052
rect 11793 20043 11851 20049
rect 11793 20040 11805 20043
rect 10928 20012 11805 20040
rect 10928 20000 10934 20012
rect 11793 20009 11805 20012
rect 11839 20009 11851 20043
rect 11793 20003 11851 20009
rect 12805 20043 12863 20049
rect 12805 20009 12817 20043
rect 12851 20040 12863 20043
rect 13354 20040 13360 20052
rect 12851 20012 13360 20040
rect 12851 20009 12863 20012
rect 12805 20003 12863 20009
rect 13354 20000 13360 20012
rect 13412 20040 13418 20052
rect 13412 20012 13584 20040
rect 13412 20000 13418 20012
rect 12894 19932 12900 19984
rect 12952 19972 12958 19984
rect 13556 19981 13584 20012
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 13872 20012 14289 20040
rect 13872 20000 13878 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 14277 20003 14335 20009
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 19797 20043 19855 20049
rect 19797 20009 19809 20043
rect 19843 20040 19855 20043
rect 20438 20040 20444 20052
rect 19843 20012 20444 20040
rect 19843 20009 19855 20012
rect 19797 20003 19855 20009
rect 20438 20000 20444 20012
rect 20496 20000 20502 20052
rect 20625 20043 20683 20049
rect 20625 20009 20637 20043
rect 20671 20040 20683 20043
rect 21174 20040 21180 20052
rect 20671 20012 21180 20040
rect 20671 20009 20683 20012
rect 20625 20003 20683 20009
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 23106 20040 23112 20052
rect 23067 20012 23112 20040
rect 23106 20000 23112 20012
rect 23164 20000 23170 20052
rect 24026 20040 24032 20052
rect 23987 20012 24032 20040
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 13449 19975 13507 19981
rect 13449 19972 13461 19975
rect 12952 19944 13461 19972
rect 12952 19932 12958 19944
rect 13449 19941 13461 19944
rect 13495 19941 13507 19975
rect 13449 19935 13507 19941
rect 13541 19975 13599 19981
rect 13541 19941 13553 19975
rect 13587 19972 13599 19975
rect 14090 19972 14096 19984
rect 13587 19944 14096 19972
rect 13587 19941 13599 19944
rect 13541 19935 13599 19941
rect 14090 19932 14096 19944
rect 14148 19932 14154 19984
rect 15562 19981 15568 19984
rect 15556 19972 15568 19981
rect 15523 19944 15568 19972
rect 15556 19935 15568 19944
rect 15562 19932 15568 19935
rect 15620 19932 15626 19984
rect 18322 19972 18328 19984
rect 18283 19944 18328 19972
rect 18322 19932 18328 19944
rect 18380 19932 18386 19984
rect 21192 19972 21220 20000
rect 22002 19981 22008 19984
rect 21974 19975 22008 19981
rect 21974 19972 21986 19975
rect 21192 19944 21986 19972
rect 21974 19941 21986 19944
rect 22060 19972 22066 19984
rect 22060 19944 22122 19972
rect 21974 19935 22008 19941
rect 22002 19932 22008 19935
rect 22060 19932 22066 19944
rect 23934 19932 23940 19984
rect 23992 19972 23998 19984
rect 24765 19975 24823 19981
rect 24765 19972 24777 19975
rect 23992 19944 24777 19972
rect 23992 19932 23998 19944
rect 24765 19941 24777 19944
rect 24811 19941 24823 19975
rect 24765 19935 24823 19941
rect 10686 19913 10692 19916
rect 10680 19904 10692 19913
rect 10647 19876 10692 19904
rect 10680 19867 10692 19876
rect 10686 19864 10692 19867
rect 10744 19864 10750 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13909 19907 13967 19913
rect 13909 19904 13921 19907
rect 12860 19876 13921 19904
rect 12860 19864 12866 19876
rect 13909 19873 13921 19876
rect 13955 19904 13967 19907
rect 13998 19904 14004 19916
rect 13955 19876 14004 19904
rect 13955 19873 13967 19876
rect 13909 19867 13967 19873
rect 13998 19864 14004 19876
rect 14056 19904 14062 19916
rect 15286 19904 15292 19916
rect 14056 19876 15292 19904
rect 14056 19864 14062 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 17589 19907 17647 19913
rect 17589 19873 17601 19907
rect 17635 19904 17647 19907
rect 17770 19904 17776 19916
rect 17635 19876 17776 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 17770 19864 17776 19876
rect 17828 19904 17834 19916
rect 17828 19876 18460 19904
rect 17828 19864 17834 19876
rect 18432 19848 18460 19876
rect 20530 19864 20536 19916
rect 20588 19904 20594 19916
rect 21729 19907 21787 19913
rect 21729 19904 21741 19907
rect 20588 19876 21741 19904
rect 20588 19864 20594 19876
rect 21729 19873 21741 19876
rect 21775 19904 21787 19907
rect 21818 19904 21824 19916
rect 21775 19876 21824 19904
rect 21775 19873 21787 19876
rect 21729 19867 21787 19873
rect 21818 19864 21824 19876
rect 21876 19864 21882 19916
rect 24026 19864 24032 19916
rect 24084 19904 24090 19916
rect 24581 19907 24639 19913
rect 24581 19904 24593 19907
rect 24084 19876 24593 19904
rect 24084 19864 24090 19876
rect 24581 19873 24593 19876
rect 24627 19873 24639 19907
rect 24581 19867 24639 19873
rect 10410 19836 10416 19848
rect 10371 19808 10416 19836
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 13446 19836 13452 19848
rect 13407 19808 13452 19836
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19805 18291 19839
rect 18414 19836 18420 19848
rect 18375 19808 18420 19836
rect 18233 19799 18291 19805
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 17000 19740 17877 19768
rect 17000 19728 17006 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 18248 19768 18276 19799
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 24857 19839 24915 19845
rect 24857 19805 24869 19839
rect 24903 19836 24915 19839
rect 25130 19836 25136 19848
rect 24903 19808 25136 19836
rect 24903 19805 24915 19808
rect 24857 19799 24915 19805
rect 18782 19768 18788 19780
rect 18248 19740 18788 19768
rect 17865 19731 17923 19737
rect 18782 19728 18788 19740
rect 18840 19728 18846 19780
rect 23753 19771 23811 19777
rect 23753 19737 23765 19771
rect 23799 19768 23811 19771
rect 24872 19768 24900 19799
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 23799 19740 24900 19768
rect 23799 19737 23811 19740
rect 23753 19731 23811 19737
rect 12986 19700 12992 19712
rect 12947 19672 12992 19700
rect 12986 19660 12992 19672
rect 13044 19660 13050 19712
rect 16666 19700 16672 19712
rect 16627 19672 16672 19700
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 24305 19703 24363 19709
rect 24305 19669 24317 19703
rect 24351 19700 24363 19703
rect 24946 19700 24952 19712
rect 24351 19672 24952 19700
rect 24351 19669 24363 19672
rect 24305 19663 24363 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 12894 19496 12900 19508
rect 12855 19468 12900 19496
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 15286 19496 15292 19508
rect 15247 19468 15292 19496
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 15620 19468 15669 19496
rect 15620 19456 15626 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 16482 19496 16488 19508
rect 16163 19468 16488 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 18414 19456 18420 19508
rect 18472 19496 18478 19508
rect 19429 19499 19487 19505
rect 19429 19496 19441 19499
rect 18472 19468 19441 19496
rect 18472 19456 18478 19468
rect 19429 19465 19441 19468
rect 19475 19465 19487 19499
rect 19429 19459 19487 19465
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22094 19496 22100 19508
rect 22060 19468 22100 19496
rect 22060 19456 22066 19468
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 23934 19496 23940 19508
rect 23895 19468 23940 19496
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 10321 19431 10379 19437
rect 10321 19397 10333 19431
rect 10367 19428 10379 19431
rect 10410 19428 10416 19440
rect 10367 19400 10416 19428
rect 10367 19397 10379 19400
rect 10321 19391 10379 19397
rect 10410 19388 10416 19400
rect 10468 19428 10474 19440
rect 10778 19428 10784 19440
rect 10468 19400 10784 19428
rect 10468 19388 10474 19400
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 15304 19428 15332 19456
rect 16574 19428 16580 19440
rect 15304 19400 16580 19428
rect 16574 19388 16580 19400
rect 16632 19428 16638 19440
rect 17494 19428 17500 19440
rect 16632 19400 17500 19428
rect 16632 19388 16638 19400
rect 17494 19388 17500 19400
rect 17552 19388 17558 19440
rect 18322 19428 18328 19440
rect 17696 19400 18328 19428
rect 17696 19360 17724 19400
rect 18322 19388 18328 19400
rect 18380 19388 18386 19440
rect 18782 19360 18788 19372
rect 17420 19332 17724 19360
rect 17880 19332 18788 19360
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 10855 19295 10913 19301
rect 9999 19264 10824 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 10134 19184 10140 19236
rect 10192 19224 10198 19236
rect 10597 19227 10655 19233
rect 10597 19224 10609 19227
rect 10192 19196 10609 19224
rect 10192 19184 10198 19196
rect 10597 19193 10609 19196
rect 10643 19193 10655 19227
rect 10796 19224 10824 19264
rect 10855 19261 10867 19295
rect 10901 19292 10913 19295
rect 11238 19292 11244 19304
rect 10901 19264 11244 19292
rect 10901 19261 10913 19264
rect 10855 19255 10913 19261
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 12802 19252 12808 19304
rect 12860 19292 12866 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12860 19264 13185 19292
rect 12860 19252 12866 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 17129 19295 17187 19301
rect 17129 19261 17141 19295
rect 17175 19292 17187 19295
rect 17420 19292 17448 19332
rect 17175 19264 17448 19292
rect 17497 19295 17555 19301
rect 17175 19261 17187 19264
rect 17129 19255 17187 19261
rect 17497 19261 17509 19295
rect 17543 19292 17555 19295
rect 17880 19292 17908 19332
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 17543 19264 17908 19292
rect 17543 19261 17555 19264
rect 17497 19255 17555 19261
rect 18322 19252 18328 19304
rect 18380 19292 18386 19304
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 18380 19264 18429 19292
rect 18380 19252 18386 19264
rect 18417 19261 18429 19264
rect 18463 19292 18475 19295
rect 19058 19292 19064 19304
rect 18463 19264 19064 19292
rect 18463 19261 18475 19264
rect 18417 19255 18475 19261
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 20530 19252 20536 19264
rect 20588 19292 20594 19304
rect 20717 19295 20775 19301
rect 20717 19292 20729 19295
rect 20588 19264 20729 19292
rect 20588 19252 20594 19264
rect 20717 19261 20729 19264
rect 20763 19261 20775 19295
rect 20717 19255 20775 19261
rect 24128 19295 24186 19301
rect 24128 19261 24140 19295
rect 24174 19292 24186 19295
rect 24174 19264 24256 19292
rect 24174 19261 24186 19264
rect 24128 19255 24186 19261
rect 11146 19224 11152 19236
rect 10796 19196 11152 19224
rect 10597 19187 10655 19193
rect 10612 19156 10640 19187
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11425 19227 11483 19233
rect 11425 19193 11437 19227
rect 11471 19193 11483 19227
rect 11425 19187 11483 19193
rect 12253 19227 12311 19233
rect 12253 19193 12265 19227
rect 12299 19224 12311 19227
rect 13354 19224 13360 19236
rect 12299 19196 13360 19224
rect 12299 19193 12311 19196
rect 12253 19187 12311 19193
rect 11333 19159 11391 19165
rect 11333 19156 11345 19159
rect 10612 19128 11345 19156
rect 11333 19125 11345 19128
rect 11379 19125 11391 19159
rect 11440 19156 11468 19187
rect 13354 19184 13360 19196
rect 13412 19233 13418 19236
rect 13412 19227 13476 19233
rect 13412 19193 13430 19227
rect 13464 19193 13476 19227
rect 17770 19224 17776 19236
rect 17731 19196 17776 19224
rect 13412 19187 13476 19193
rect 13412 19184 13418 19187
rect 17770 19184 17776 19196
rect 17828 19184 17834 19236
rect 18138 19233 18144 19236
rect 18123 19227 18144 19233
rect 18123 19193 18135 19227
rect 18123 19187 18144 19193
rect 18138 19184 18144 19187
rect 18196 19184 18202 19236
rect 18690 19224 18696 19236
rect 18651 19196 18696 19224
rect 18690 19184 18696 19196
rect 18748 19184 18754 19236
rect 20257 19227 20315 19233
rect 20257 19193 20269 19227
rect 20303 19224 20315 19227
rect 20984 19227 21042 19233
rect 20984 19224 20996 19227
rect 20303 19196 20996 19224
rect 20303 19193 20315 19196
rect 20257 19187 20315 19193
rect 20984 19193 20996 19196
rect 21030 19224 21042 19227
rect 21634 19224 21640 19236
rect 21030 19196 21640 19224
rect 21030 19193 21042 19196
rect 20984 19187 21042 19193
rect 21634 19184 21640 19196
rect 21692 19184 21698 19236
rect 21818 19184 21824 19236
rect 21876 19224 21882 19236
rect 21876 19196 23520 19224
rect 21876 19184 21882 19196
rect 11882 19156 11888 19168
rect 11440 19128 11888 19156
rect 11333 19119 11391 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 13814 19116 13820 19168
rect 13872 19156 13878 19168
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 13872 19128 14565 19156
rect 13872 19116 13878 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 17788 19156 17816 19184
rect 18601 19159 18659 19165
rect 18601 19156 18613 19159
rect 17788 19128 18613 19156
rect 14553 19119 14611 19125
rect 18601 19125 18613 19128
rect 18647 19125 18659 19159
rect 18601 19119 18659 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 23492 19165 23520 19196
rect 22649 19159 22707 19165
rect 22649 19156 22661 19159
rect 22152 19128 22661 19156
rect 22152 19116 22158 19128
rect 22649 19125 22661 19128
rect 22695 19125 22707 19159
rect 22649 19119 22707 19125
rect 23477 19159 23535 19165
rect 23477 19125 23489 19159
rect 23523 19156 23535 19159
rect 23658 19156 23664 19168
rect 23523 19128 23664 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23658 19116 23664 19128
rect 23716 19156 23722 19168
rect 24228 19156 24256 19264
rect 25314 19252 25320 19304
rect 25372 19292 25378 19304
rect 26234 19292 26240 19304
rect 25372 19264 26240 19292
rect 25372 19252 25378 19264
rect 26234 19252 26240 19264
rect 26292 19252 26298 19304
rect 24388 19227 24446 19233
rect 24388 19193 24400 19227
rect 24434 19224 24446 19227
rect 25130 19224 25136 19236
rect 24434 19196 25136 19224
rect 24434 19193 24446 19196
rect 24388 19187 24446 19193
rect 25130 19184 25136 19196
rect 25188 19184 25194 19236
rect 25498 19156 25504 19168
rect 23716 19128 24256 19156
rect 25459 19128 25504 19156
rect 23716 19116 23722 19128
rect 25498 19116 25504 19128
rect 25556 19116 25562 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13044 18924 13737 18952
rect 13044 18912 13050 18924
rect 13725 18921 13737 18924
rect 13771 18952 13783 18955
rect 13998 18952 14004 18964
rect 13771 18924 14004 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 21818 18912 21824 18964
rect 21876 18952 21882 18964
rect 21913 18955 21971 18961
rect 21913 18952 21925 18955
rect 21876 18924 21925 18952
rect 21876 18912 21882 18924
rect 21913 18921 21925 18924
rect 21959 18921 21971 18955
rect 25130 18952 25136 18964
rect 25091 18924 25136 18952
rect 21913 18915 21971 18921
rect 25130 18912 25136 18924
rect 25188 18912 25194 18964
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 13538 18884 13544 18896
rect 11204 18856 13032 18884
rect 13499 18856 13544 18884
rect 11204 18844 11210 18856
rect 10778 18776 10784 18828
rect 10836 18776 10842 18828
rect 10956 18819 11014 18825
rect 10956 18785 10968 18819
rect 11002 18816 11014 18819
rect 11882 18816 11888 18828
rect 11002 18788 11888 18816
rect 11002 18785 11014 18788
rect 10956 18779 11014 18785
rect 11882 18776 11888 18788
rect 11940 18776 11946 18828
rect 13004 18825 13032 18856
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 13814 18884 13820 18896
rect 13775 18856 13820 18884
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 16666 18844 16672 18896
rect 16724 18884 16730 18896
rect 16914 18887 16972 18893
rect 16914 18884 16926 18887
rect 16724 18856 16926 18884
rect 16724 18844 16730 18856
rect 16914 18853 16926 18856
rect 16960 18853 16972 18887
rect 16914 18847 16972 18853
rect 21358 18844 21364 18896
rect 21416 18884 21422 18896
rect 21453 18887 21511 18893
rect 21453 18884 21465 18887
rect 21416 18856 21465 18884
rect 21416 18844 21422 18856
rect 21453 18853 21465 18856
rect 21499 18853 21511 18887
rect 21453 18847 21511 18853
rect 12989 18819 13047 18825
rect 12989 18785 13001 18819
rect 13035 18816 13047 18819
rect 13446 18816 13452 18828
rect 13035 18788 13452 18816
rect 13035 18785 13047 18788
rect 12989 18779 13047 18785
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 24009 18819 24067 18825
rect 24009 18816 24021 18819
rect 23532 18788 24021 18816
rect 23532 18776 23538 18788
rect 24009 18785 24021 18788
rect 24055 18785 24067 18819
rect 24009 18779 24067 18785
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 10652 18720 10701 18748
rect 10652 18708 10658 18720
rect 10689 18717 10701 18720
rect 10735 18748 10747 18751
rect 10796 18748 10824 18776
rect 10735 18720 10824 18748
rect 10735 18717 10747 18720
rect 10689 18711 10747 18717
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15381 18751 15439 18757
rect 15381 18748 15393 18751
rect 15344 18720 15393 18748
rect 15344 18708 15350 18720
rect 15381 18717 15393 18720
rect 15427 18717 15439 18751
rect 15381 18711 15439 18717
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16632 18720 16681 18748
rect 16632 18708 16638 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 21450 18748 21456 18760
rect 21411 18720 21456 18748
rect 16669 18711 16727 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18748 21603 18751
rect 21634 18748 21640 18760
rect 21591 18720 21640 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 23658 18708 23664 18760
rect 23716 18748 23722 18760
rect 23753 18751 23811 18757
rect 23753 18748 23765 18751
rect 23716 18720 23765 18748
rect 23716 18708 23722 18720
rect 23753 18717 23765 18720
rect 23799 18717 23811 18751
rect 23753 18711 23811 18717
rect 20714 18640 20720 18692
rect 20772 18680 20778 18692
rect 20993 18683 21051 18689
rect 20993 18680 21005 18683
rect 20772 18652 21005 18680
rect 20772 18640 20778 18652
rect 20993 18649 21005 18652
rect 21039 18649 21051 18683
rect 20993 18643 21051 18649
rect 10410 18612 10416 18624
rect 10371 18584 10416 18612
rect 10410 18572 10416 18584
rect 10468 18612 10474 18624
rect 10686 18612 10692 18624
rect 10468 18584 10692 18612
rect 10468 18572 10474 18584
rect 10686 18572 10692 18584
rect 10744 18612 10750 18624
rect 12069 18615 12127 18621
rect 12069 18612 12081 18615
rect 10744 18584 12081 18612
rect 10744 18572 10750 18584
rect 12069 18581 12081 18584
rect 12115 18581 12127 18615
rect 12069 18575 12127 18581
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 13722 18612 13728 18624
rect 13311 18584 13728 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 18046 18612 18052 18624
rect 18007 18584 18052 18612
rect 18046 18572 18052 18584
rect 18104 18612 18110 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18104 18584 18613 18612
rect 18104 18572 18110 18584
rect 18601 18581 18613 18584
rect 18647 18612 18659 18615
rect 18690 18612 18696 18624
rect 18647 18584 18696 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 9861 18411 9919 18417
rect 9861 18377 9873 18411
rect 9907 18408 9919 18411
rect 10410 18408 10416 18420
rect 9907 18380 10416 18408
rect 9907 18377 9919 18380
rect 9861 18371 9919 18377
rect 10410 18368 10416 18380
rect 10468 18408 10474 18420
rect 12897 18411 12955 18417
rect 10468 18380 11376 18408
rect 10468 18368 10474 18380
rect 10781 18343 10839 18349
rect 10781 18309 10793 18343
rect 10827 18340 10839 18343
rect 10962 18340 10968 18352
rect 10827 18312 10968 18340
rect 10827 18309 10839 18312
rect 10781 18303 10839 18309
rect 10962 18300 10968 18312
rect 11020 18300 11026 18352
rect 11348 18281 11376 18380
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 13538 18408 13544 18420
rect 12943 18380 13544 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 13998 18408 14004 18420
rect 13959 18380 14004 18408
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 15197 18411 15255 18417
rect 15197 18377 15209 18411
rect 15243 18408 15255 18411
rect 15286 18408 15292 18420
rect 15243 18380 15292 18408
rect 15243 18377 15255 18380
rect 15197 18371 15255 18377
rect 15286 18368 15292 18380
rect 15344 18408 15350 18420
rect 15344 18380 15516 18408
rect 15344 18368 15350 18380
rect 13265 18343 13323 18349
rect 13265 18309 13277 18343
rect 13311 18340 13323 18343
rect 13814 18340 13820 18352
rect 13311 18312 13820 18340
rect 13311 18309 13323 18312
rect 13265 18303 13323 18309
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 15378 18340 15384 18352
rect 15339 18312 15384 18340
rect 15378 18300 15384 18312
rect 15436 18300 15442 18352
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18241 11391 18275
rect 15488 18272 15516 18380
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 17037 18411 17095 18417
rect 17037 18408 17049 18411
rect 16724 18380 17049 18408
rect 16724 18368 16730 18380
rect 17037 18377 17049 18380
rect 17083 18377 17095 18411
rect 17037 18371 17095 18377
rect 20993 18411 21051 18417
rect 20993 18377 21005 18411
rect 21039 18408 21051 18411
rect 21450 18408 21456 18420
rect 21039 18380 21456 18408
rect 21039 18377 21051 18380
rect 20993 18371 21051 18377
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 23474 18408 23480 18420
rect 23435 18380 23480 18408
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 24305 18411 24363 18417
rect 24305 18377 24317 18411
rect 24351 18408 24363 18411
rect 24351 18380 25084 18408
rect 24351 18377 24363 18380
rect 24305 18371 24363 18377
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 16761 18343 16819 18349
rect 16761 18340 16773 18343
rect 16632 18312 16773 18340
rect 16632 18300 16638 18312
rect 16761 18309 16773 18312
rect 16807 18309 16819 18343
rect 16761 18303 16819 18309
rect 23658 18300 23664 18352
rect 23716 18340 23722 18352
rect 24489 18343 24547 18349
rect 24489 18340 24501 18343
rect 23716 18312 24501 18340
rect 23716 18300 23722 18312
rect 24489 18309 24501 18312
rect 24535 18309 24547 18343
rect 24489 18303 24547 18309
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15488 18244 15761 18272
rect 11333 18235 11391 18241
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 24854 18272 24860 18284
rect 24815 18244 24860 18272
rect 15749 18235 15807 18241
rect 24854 18232 24860 18244
rect 24912 18232 24918 18284
rect 25056 18281 25084 18380
rect 25041 18275 25099 18281
rect 25041 18241 25053 18275
rect 25087 18272 25099 18275
rect 25498 18272 25504 18284
rect 25087 18244 25504 18272
rect 25087 18241 25099 18244
rect 25041 18235 25099 18241
rect 25498 18232 25504 18244
rect 25556 18232 25562 18284
rect 16666 18204 16672 18216
rect 15948 18176 16672 18204
rect 10229 18139 10287 18145
rect 10229 18105 10241 18139
rect 10275 18136 10287 18139
rect 10778 18136 10784 18148
rect 10275 18108 10784 18136
rect 10275 18105 10287 18108
rect 10229 18099 10287 18105
rect 10778 18096 10784 18108
rect 10836 18136 10842 18148
rect 11057 18139 11115 18145
rect 11057 18136 11069 18139
rect 10836 18108 11069 18136
rect 10836 18096 10842 18108
rect 11057 18105 11069 18108
rect 11103 18105 11115 18139
rect 11238 18136 11244 18148
rect 11199 18108 11244 18136
rect 11057 18099 11115 18105
rect 11238 18096 11244 18108
rect 11296 18096 11302 18148
rect 15948 18145 15976 18176
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 25409 18207 25467 18213
rect 25409 18204 25421 18207
rect 24964 18176 25421 18204
rect 24964 18148 24992 18176
rect 25409 18173 25421 18176
rect 25455 18173 25467 18207
rect 25409 18167 25467 18173
rect 14829 18139 14887 18145
rect 14829 18105 14841 18139
rect 14875 18136 14887 18139
rect 15933 18139 15991 18145
rect 15933 18136 15945 18139
rect 14875 18108 15945 18136
rect 14875 18105 14887 18108
rect 14829 18099 14887 18105
rect 15933 18105 15945 18108
rect 15979 18105 15991 18139
rect 24946 18136 24952 18148
rect 24907 18108 24952 18136
rect 15933 18099 15991 18105
rect 24946 18096 24952 18108
rect 25004 18096 25010 18148
rect 10597 18071 10655 18077
rect 10597 18037 10609 18071
rect 10643 18068 10655 18071
rect 10686 18068 10692 18080
rect 10643 18040 10692 18068
rect 10643 18037 10655 18040
rect 10597 18031 10655 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11793 18071 11851 18077
rect 11793 18037 11805 18071
rect 11839 18068 11851 18071
rect 11882 18068 11888 18080
rect 11839 18040 11888 18068
rect 11839 18037 11851 18040
rect 11793 18031 11851 18037
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 13538 18068 13544 18080
rect 13499 18040 13544 18068
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15528 18040 15853 18068
rect 15528 18028 15534 18040
rect 15841 18037 15853 18040
rect 15887 18037 15899 18071
rect 15841 18031 15899 18037
rect 16298 18028 16304 18080
rect 16356 18068 16362 18080
rect 16574 18068 16580 18080
rect 16356 18040 16580 18068
rect 16356 18028 16362 18040
rect 16574 18028 16580 18040
rect 16632 18068 16638 18080
rect 17954 18068 17960 18080
rect 16632 18040 17960 18068
rect 16632 18028 16638 18040
rect 17954 18028 17960 18040
rect 18012 18028 18018 18080
rect 18690 18068 18696 18080
rect 18651 18040 18696 18068
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 21358 18068 21364 18080
rect 21319 18040 21364 18068
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 21634 18068 21640 18080
rect 21595 18040 21640 18068
rect 21634 18028 21640 18040
rect 21692 18028 21698 18080
rect 23382 18028 23388 18080
rect 23440 18068 23446 18080
rect 23566 18068 23572 18080
rect 23440 18040 23572 18068
rect 23440 18028 23446 18040
rect 23566 18028 23572 18040
rect 23624 18068 23630 18080
rect 23845 18071 23903 18077
rect 23845 18068 23857 18071
rect 23624 18040 23857 18068
rect 23624 18028 23630 18040
rect 23845 18037 23857 18040
rect 23891 18037 23903 18071
rect 23845 18031 23903 18037
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 10778 17864 10784 17876
rect 10739 17836 10784 17864
rect 10778 17824 10784 17836
rect 10836 17824 10842 17876
rect 11238 17864 11244 17876
rect 11199 17836 11244 17864
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 13538 17864 13544 17876
rect 13403 17836 13544 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 13538 17824 13544 17836
rect 13596 17864 13602 17876
rect 15470 17864 15476 17876
rect 13596 17836 13860 17864
rect 15431 17836 15476 17864
rect 13596 17824 13602 17836
rect 13832 17805 13860 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 18138 17864 18144 17876
rect 18099 17836 18144 17864
rect 18138 17824 18144 17836
rect 18196 17824 18202 17876
rect 24673 17867 24731 17873
rect 24673 17833 24685 17867
rect 24719 17864 24731 17867
rect 24762 17864 24768 17876
rect 24719 17836 24768 17864
rect 24719 17833 24731 17836
rect 24673 17827 24731 17833
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 13817 17799 13875 17805
rect 13817 17765 13829 17799
rect 13863 17765 13875 17799
rect 13817 17759 13875 17765
rect 14001 17799 14059 17805
rect 14001 17765 14013 17799
rect 14047 17796 14059 17799
rect 14458 17796 14464 17808
rect 14047 17768 14464 17796
rect 14047 17765 14059 17768
rect 14001 17759 14059 17765
rect 14458 17756 14464 17768
rect 14516 17756 14522 17808
rect 21450 17796 21456 17808
rect 21411 17768 21456 17796
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 23198 17756 23204 17808
rect 23256 17796 23262 17808
rect 23753 17799 23811 17805
rect 23753 17796 23765 17799
rect 23256 17768 23765 17796
rect 23256 17756 23262 17768
rect 23753 17765 23765 17768
rect 23799 17765 23811 17799
rect 23753 17759 23811 17765
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 18046 17728 18052 17740
rect 17552 17700 18052 17728
rect 17552 17688 17558 17700
rect 18046 17688 18052 17700
rect 18104 17728 18110 17740
rect 18581 17731 18639 17737
rect 18581 17728 18593 17731
rect 18104 17700 18593 17728
rect 18104 17688 18110 17700
rect 18581 17697 18593 17700
rect 18627 17697 18639 17731
rect 18581 17691 18639 17697
rect 22830 17688 22836 17740
rect 22888 17728 22894 17740
rect 23569 17731 23627 17737
rect 23569 17728 23581 17731
rect 22888 17700 23581 17728
rect 22888 17688 22894 17700
rect 23569 17697 23581 17700
rect 23615 17697 23627 17731
rect 23569 17691 23627 17697
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13872 17632 14105 17660
rect 13872 17620 13878 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18012 17632 18337 17660
rect 18012 17620 18018 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 21361 17663 21419 17669
rect 21361 17629 21373 17663
rect 21407 17629 21419 17663
rect 21542 17660 21548 17672
rect 21503 17632 21548 17660
rect 21361 17623 21419 17629
rect 21376 17592 21404 17623
rect 21542 17620 21548 17632
rect 21600 17620 21606 17672
rect 23842 17660 23848 17672
rect 23803 17632 23848 17660
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 24210 17620 24216 17672
rect 24268 17660 24274 17672
rect 24305 17663 24363 17669
rect 24305 17660 24317 17663
rect 24268 17632 24317 17660
rect 24268 17620 24274 17632
rect 24305 17629 24317 17632
rect 24351 17660 24363 17663
rect 24765 17663 24823 17669
rect 24765 17660 24777 17663
rect 24351 17632 24777 17660
rect 24351 17629 24363 17632
rect 24305 17623 24363 17629
rect 24765 17629 24777 17632
rect 24811 17629 24823 17663
rect 24765 17623 24823 17629
rect 21818 17592 21824 17604
rect 21376 17564 21824 17592
rect 21818 17552 21824 17564
rect 21876 17552 21882 17604
rect 13538 17524 13544 17536
rect 13499 17496 13544 17524
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 16393 17527 16451 17533
rect 16393 17493 16405 17527
rect 16439 17524 16451 17527
rect 16850 17524 16856 17536
rect 16439 17496 16856 17524
rect 16439 17493 16451 17496
rect 16393 17487 16451 17493
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 19702 17524 19708 17536
rect 19663 17496 19708 17524
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 20993 17527 21051 17533
rect 20993 17493 21005 17527
rect 21039 17524 21051 17527
rect 21910 17524 21916 17536
rect 21039 17496 21916 17524
rect 21039 17493 21051 17496
rect 20993 17487 21051 17493
rect 21910 17484 21916 17496
rect 21968 17484 21974 17536
rect 23293 17527 23351 17533
rect 23293 17493 23305 17527
rect 23339 17524 23351 17527
rect 23474 17524 23480 17536
rect 23339 17496 23480 17524
rect 23339 17493 23351 17496
rect 23293 17487 23351 17493
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 16298 17320 16304 17332
rect 15804 17292 16304 17320
rect 15804 17280 15810 17292
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 17494 17320 17500 17332
rect 17455 17292 17500 17320
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 18322 17320 18328 17332
rect 18012 17292 18328 17320
rect 18012 17280 18018 17292
rect 18322 17280 18328 17292
rect 18380 17320 18386 17332
rect 19061 17323 19119 17329
rect 19061 17320 19073 17323
rect 18380 17292 19073 17320
rect 18380 17280 18386 17292
rect 19061 17289 19073 17292
rect 19107 17289 19119 17323
rect 19061 17283 19119 17289
rect 19521 17323 19579 17329
rect 19521 17289 19533 17323
rect 19567 17320 19579 17323
rect 20530 17320 20536 17332
rect 19567 17292 20536 17320
rect 19567 17289 19579 17292
rect 19521 17283 19579 17289
rect 16114 17252 16120 17264
rect 16075 17224 16120 17252
rect 16114 17212 16120 17224
rect 16172 17212 16178 17264
rect 16393 17255 16451 17261
rect 16393 17221 16405 17255
rect 16439 17252 16451 17255
rect 16574 17252 16580 17264
rect 16439 17224 16580 17252
rect 16439 17221 16451 17224
rect 16393 17215 16451 17221
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 18138 17252 18144 17264
rect 18099 17224 18144 17252
rect 18138 17212 18144 17224
rect 18196 17212 18202 17264
rect 12802 17076 12808 17128
rect 12860 17116 12866 17128
rect 12989 17119 13047 17125
rect 12989 17116 13001 17119
rect 12860 17088 13001 17116
rect 12860 17076 12866 17088
rect 12989 17085 13001 17088
rect 13035 17085 13047 17119
rect 12989 17079 13047 17085
rect 13256 17119 13314 17125
rect 13256 17085 13268 17119
rect 13302 17116 13314 17119
rect 13814 17116 13820 17128
rect 13302 17088 13820 17116
rect 13302 17085 13314 17088
rect 13256 17079 13314 17085
rect 13372 17060 13400 17088
rect 13814 17076 13820 17088
rect 13872 17076 13878 17128
rect 16132 17116 16160 17212
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18601 17187 18659 17193
rect 18601 17184 18613 17187
rect 17911 17156 18613 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18601 17153 18613 17156
rect 18647 17184 18659 17187
rect 18690 17184 18696 17196
rect 18647 17156 18696 17184
rect 18647 17153 18659 17156
rect 18601 17147 18659 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 19628 17193 19656 17292
rect 20530 17280 20536 17292
rect 20588 17280 20594 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 21082 17320 21088 17332
rect 21039 17292 21088 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 21082 17280 21088 17292
rect 21140 17320 21146 17332
rect 21542 17320 21548 17332
rect 21140 17292 21548 17320
rect 21140 17280 21146 17292
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 22830 17320 22836 17332
rect 22791 17292 22836 17320
rect 22830 17280 22836 17292
rect 22888 17280 22894 17332
rect 23845 17255 23903 17261
rect 23845 17221 23857 17255
rect 23891 17252 23903 17255
rect 24026 17252 24032 17264
rect 23891 17224 24032 17252
rect 23891 17221 23903 17224
rect 23845 17215 23903 17221
rect 24026 17212 24032 17224
rect 24084 17212 24090 17264
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 21450 17144 21456 17196
rect 21508 17184 21514 17196
rect 21545 17187 21603 17193
rect 21545 17184 21557 17187
rect 21508 17156 21557 17184
rect 21508 17144 21514 17156
rect 21545 17153 21557 17156
rect 21591 17153 21603 17187
rect 24210 17184 24216 17196
rect 24171 17156 24216 17184
rect 21545 17147 21603 17153
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 23198 17116 23204 17128
rect 16132 17088 16896 17116
rect 23159 17088 23204 17116
rect 12253 17051 12311 17057
rect 12253 17017 12265 17051
rect 12299 17048 12311 17051
rect 13354 17048 13360 17060
rect 12299 17020 13360 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 13354 17008 13360 17020
rect 13412 17008 13418 17060
rect 16868 17057 16896 17088
rect 23198 17076 23204 17088
rect 23256 17076 23262 17128
rect 16853 17051 16911 17057
rect 16853 17017 16865 17051
rect 16899 17017 16911 17051
rect 16853 17011 16911 17017
rect 16942 17008 16948 17060
rect 17000 17048 17006 17060
rect 17000 17020 17045 17048
rect 17000 17008 17006 17020
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18601 17051 18659 17057
rect 18601 17048 18613 17051
rect 18288 17020 18613 17048
rect 18288 17008 18294 17020
rect 18601 17017 18613 17020
rect 18647 17017 18659 17051
rect 18601 17011 18659 17017
rect 18690 17008 18696 17060
rect 18748 17048 18754 17060
rect 19702 17048 19708 17060
rect 18748 17020 19708 17048
rect 18748 17008 18754 17020
rect 19702 17008 19708 17020
rect 19760 17048 19766 17060
rect 19858 17051 19916 17057
rect 19858 17048 19870 17051
rect 19760 17020 19870 17048
rect 19760 17008 19766 17020
rect 19858 17017 19870 17020
rect 19904 17017 19916 17051
rect 19858 17011 19916 17017
rect 23842 17008 23848 17060
rect 23900 17048 23906 17060
rect 24394 17048 24400 17060
rect 23900 17020 24400 17048
rect 23900 17008 23906 17020
rect 24394 17008 24400 17020
rect 24452 17048 24458 17060
rect 24765 17051 24823 17057
rect 24765 17048 24777 17051
rect 24452 17020 24777 17048
rect 24452 17008 24458 17020
rect 24765 17017 24777 17020
rect 24811 17017 24823 17051
rect 24765 17011 24823 17017
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 14366 16980 14372 16992
rect 14327 16952 14372 16980
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 14458 16940 14464 16992
rect 14516 16980 14522 16992
rect 15010 16980 15016 16992
rect 14516 16952 15016 16980
rect 14516 16940 14522 16952
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 15930 16980 15936 16992
rect 15887 16952 15936 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 15930 16940 15936 16952
rect 15988 16980 15994 16992
rect 16960 16980 16988 17008
rect 15988 16952 16988 16980
rect 15988 16940 15994 16952
rect 21818 16940 21824 16992
rect 21876 16980 21882 16992
rect 21913 16983 21971 16989
rect 21913 16980 21925 16983
rect 21876 16952 21925 16980
rect 21876 16940 21882 16952
rect 21913 16949 21925 16952
rect 21959 16949 21971 16983
rect 21913 16943 21971 16949
rect 22002 16940 22008 16992
rect 22060 16980 22066 16992
rect 22097 16983 22155 16989
rect 22097 16980 22109 16983
rect 22060 16952 22109 16980
rect 22060 16940 22066 16952
rect 22097 16949 22109 16952
rect 22143 16949 22155 16983
rect 22097 16943 22155 16949
rect 24118 16940 24124 16992
rect 24176 16980 24182 16992
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 24176 16952 24317 16980
rect 24176 16940 24182 16952
rect 24305 16949 24317 16952
rect 24351 16949 24363 16983
rect 24305 16943 24363 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12253 16779 12311 16785
rect 12253 16776 12265 16779
rect 11940 16748 12265 16776
rect 11940 16736 11946 16748
rect 12253 16745 12265 16748
rect 12299 16745 12311 16779
rect 12253 16739 12311 16745
rect 13265 16779 13323 16785
rect 13265 16745 13277 16779
rect 13311 16776 13323 16779
rect 13354 16776 13360 16788
rect 13311 16748 13360 16776
rect 13311 16745 13323 16748
rect 13265 16739 13323 16745
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 13909 16779 13967 16785
rect 13909 16776 13921 16779
rect 13872 16748 13921 16776
rect 13872 16736 13878 16748
rect 13909 16745 13921 16748
rect 13955 16745 13967 16779
rect 13909 16739 13967 16745
rect 18141 16779 18199 16785
rect 18141 16745 18153 16779
rect 18187 16776 18199 16779
rect 18690 16776 18696 16788
rect 18187 16748 18696 16776
rect 18187 16745 18199 16748
rect 18141 16739 18199 16745
rect 18690 16736 18696 16748
rect 18748 16776 18754 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 18748 16748 19625 16776
rect 18748 16736 18754 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 23845 16779 23903 16785
rect 23845 16745 23857 16779
rect 23891 16776 23903 16779
rect 24118 16776 24124 16788
rect 23891 16748 24124 16776
rect 23891 16745 23903 16748
rect 23845 16739 23903 16745
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 24854 16736 24860 16788
rect 24912 16776 24918 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 24912 16748 25329 16776
rect 24912 16736 24918 16748
rect 25317 16745 25329 16748
rect 25363 16745 25375 16779
rect 25317 16739 25375 16745
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 13725 16711 13783 16717
rect 13725 16708 13737 16711
rect 13596 16680 13737 16708
rect 13596 16668 13602 16680
rect 13725 16677 13737 16680
rect 13771 16677 13783 16711
rect 13725 16671 13783 16677
rect 14001 16711 14059 16717
rect 14001 16677 14013 16711
rect 14047 16708 14059 16711
rect 14366 16708 14372 16720
rect 14047 16680 14372 16708
rect 14047 16677 14059 16680
rect 14001 16671 14059 16677
rect 14366 16668 14372 16680
rect 14424 16668 14430 16720
rect 15930 16668 15936 16720
rect 15988 16717 15994 16720
rect 15988 16711 16052 16717
rect 15988 16677 16006 16711
rect 16040 16677 16052 16711
rect 18782 16708 18788 16720
rect 18743 16680 18788 16708
rect 15988 16671 16052 16677
rect 15988 16668 15994 16671
rect 18782 16668 18788 16680
rect 18840 16668 18846 16720
rect 20717 16711 20775 16717
rect 20717 16677 20729 16711
rect 20763 16708 20775 16711
rect 21082 16708 21088 16720
rect 20763 16680 21088 16708
rect 20763 16677 20775 16680
rect 20717 16671 20775 16677
rect 21082 16668 21088 16680
rect 21140 16708 21146 16720
rect 21238 16711 21296 16717
rect 21238 16708 21250 16711
rect 21140 16680 21250 16708
rect 21140 16668 21146 16680
rect 21238 16677 21250 16680
rect 21284 16677 21296 16711
rect 21238 16671 21296 16677
rect 23106 16668 23112 16720
rect 23164 16708 23170 16720
rect 23293 16711 23351 16717
rect 23293 16708 23305 16711
rect 23164 16680 23305 16708
rect 23164 16668 23170 16680
rect 23293 16677 23305 16680
rect 23339 16708 23351 16711
rect 24204 16711 24262 16717
rect 24204 16708 24216 16711
rect 23339 16680 24216 16708
rect 23339 16677 23351 16680
rect 23293 16671 23351 16677
rect 24204 16677 24216 16680
rect 24250 16708 24262 16711
rect 24394 16708 24400 16720
rect 24250 16680 24400 16708
rect 24250 16677 24262 16680
rect 24204 16671 24262 16677
rect 24394 16668 24400 16680
rect 24452 16668 24458 16720
rect 10686 16600 10692 16652
rect 10744 16640 10750 16652
rect 11146 16649 11152 16652
rect 10873 16643 10931 16649
rect 10873 16640 10885 16643
rect 10744 16612 10885 16640
rect 10744 16600 10750 16612
rect 10873 16609 10885 16612
rect 10919 16609 10931 16643
rect 10873 16603 10931 16609
rect 11140 16603 11152 16649
rect 11204 16640 11210 16652
rect 18598 16640 18604 16652
rect 11204 16612 11240 16640
rect 18559 16612 18604 16640
rect 11146 16600 11152 16603
rect 11204 16600 11210 16612
rect 18598 16600 18604 16612
rect 18656 16600 18662 16652
rect 23382 16600 23388 16652
rect 23440 16640 23446 16652
rect 23937 16643 23995 16649
rect 23937 16640 23949 16643
rect 23440 16612 23949 16640
rect 23440 16600 23446 16612
rect 23937 16609 23949 16612
rect 23983 16640 23995 16643
rect 24670 16640 24676 16652
rect 23983 16612 24676 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24670 16600 24676 16612
rect 24728 16600 24734 16652
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 18874 16572 18880 16584
rect 17000 16544 18880 16572
rect 17000 16532 17006 16544
rect 18874 16532 18880 16544
rect 18932 16532 18938 16584
rect 21000 16575 21058 16581
rect 21000 16572 21012 16575
rect 20916 16544 21012 16572
rect 17126 16504 17132 16516
rect 17087 16476 17132 16504
rect 17126 16464 17132 16476
rect 17184 16464 17190 16516
rect 13446 16436 13452 16448
rect 13407 16408 13452 16436
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 16758 16396 16764 16448
rect 16816 16436 16822 16448
rect 18325 16439 18383 16445
rect 18325 16436 18337 16439
rect 16816 16408 18337 16436
rect 16816 16396 16822 16408
rect 18325 16405 18337 16408
rect 18371 16405 18383 16439
rect 18325 16399 18383 16405
rect 18414 16396 18420 16448
rect 18472 16436 18478 16448
rect 19150 16436 19156 16448
rect 18472 16408 19156 16436
rect 18472 16396 18478 16408
rect 19150 16396 19156 16408
rect 19208 16436 19214 16448
rect 20530 16436 20536 16448
rect 19208 16408 20536 16436
rect 19208 16396 19214 16408
rect 20530 16396 20536 16408
rect 20588 16436 20594 16448
rect 20916 16436 20944 16544
rect 21000 16541 21012 16544
rect 21046 16541 21058 16575
rect 21000 16535 21058 16541
rect 20990 16436 20996 16448
rect 20588 16408 20996 16436
rect 20588 16396 20594 16408
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 22370 16436 22376 16448
rect 22331 16408 22376 16436
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11241 16235 11299 16241
rect 11241 16232 11253 16235
rect 11204 16204 11253 16232
rect 11204 16192 11210 16204
rect 11241 16201 11253 16204
rect 11287 16201 11299 16235
rect 11241 16195 11299 16201
rect 13081 16235 13139 16241
rect 13081 16201 13093 16235
rect 13127 16232 13139 16235
rect 13722 16232 13728 16244
rect 13127 16204 13728 16232
rect 13127 16201 13139 16204
rect 13081 16195 13139 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15565 16235 15623 16241
rect 15565 16201 15577 16235
rect 15611 16232 15623 16235
rect 16577 16235 16635 16241
rect 16577 16232 16589 16235
rect 15611 16204 16589 16232
rect 15611 16201 15623 16204
rect 15565 16195 15623 16201
rect 16577 16201 16589 16204
rect 16623 16232 16635 16235
rect 16942 16232 16948 16244
rect 16623 16204 16948 16232
rect 16623 16201 16635 16204
rect 16577 16195 16635 16201
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 18325 16235 18383 16241
rect 18325 16201 18337 16235
rect 18371 16232 18383 16235
rect 18782 16232 18788 16244
rect 18371 16204 18788 16232
rect 18371 16201 18383 16204
rect 18325 16195 18383 16201
rect 18782 16192 18788 16204
rect 18840 16192 18846 16244
rect 18874 16192 18880 16244
rect 18932 16232 18938 16244
rect 18969 16235 19027 16241
rect 18969 16232 18981 16235
rect 18932 16204 18981 16232
rect 18932 16192 18938 16204
rect 18969 16201 18981 16204
rect 19015 16201 19027 16235
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 18969 16195 19027 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23477 16235 23535 16241
rect 23477 16201 23489 16235
rect 23523 16232 23535 16235
rect 23566 16232 23572 16244
rect 23523 16204 23572 16232
rect 23523 16201 23535 16204
rect 23477 16195 23535 16201
rect 23566 16192 23572 16204
rect 23624 16232 23630 16244
rect 24762 16232 24768 16244
rect 23624 16204 24768 16232
rect 23624 16192 23630 16204
rect 10686 16124 10692 16176
rect 10744 16164 10750 16176
rect 10873 16167 10931 16173
rect 10873 16164 10885 16167
rect 10744 16136 10885 16164
rect 10744 16124 10750 16136
rect 10873 16133 10885 16136
rect 10919 16133 10931 16167
rect 10873 16127 10931 16133
rect 21545 16167 21603 16173
rect 21545 16133 21557 16167
rect 21591 16164 21603 16167
rect 21818 16164 21824 16176
rect 21591 16136 21824 16164
rect 21591 16133 21603 16136
rect 21545 16127 21603 16133
rect 21818 16124 21824 16136
rect 21876 16124 21882 16176
rect 23753 16167 23811 16173
rect 23753 16133 23765 16167
rect 23799 16164 23811 16167
rect 23842 16164 23848 16176
rect 23799 16136 23848 16164
rect 23799 16133 23811 16136
rect 23753 16127 23811 16133
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 18598 16096 18604 16108
rect 16899 16068 18604 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16056 22066 16108
rect 24320 16105 24348 16204
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25406 16232 25412 16244
rect 25367 16204 25412 16232
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 25866 16232 25872 16244
rect 25827 16204 25872 16232
rect 25866 16192 25872 16204
rect 25924 16192 25930 16244
rect 24670 16164 24676 16176
rect 24631 16136 24676 16164
rect 24670 16124 24676 16136
rect 24728 16124 24734 16176
rect 24305 16099 24363 16105
rect 24305 16065 24317 16099
rect 24351 16065 24363 16099
rect 24305 16059 24363 16065
rect 14185 16031 14243 16037
rect 14185 15997 14197 16031
rect 14231 16028 14243 16031
rect 20717 16031 20775 16037
rect 14231 16000 14596 16028
rect 14231 15997 14243 16000
rect 14185 15991 14243 15997
rect 13449 15963 13507 15969
rect 13449 15929 13461 15963
rect 13495 15960 13507 15963
rect 14366 15960 14372 15972
rect 13495 15932 14372 15960
rect 13495 15929 13507 15932
rect 13449 15923 13507 15929
rect 14366 15920 14372 15932
rect 14424 15969 14430 15972
rect 14424 15963 14488 15969
rect 14424 15929 14442 15963
rect 14476 15929 14488 15963
rect 14424 15923 14488 15929
rect 14424 15920 14430 15923
rect 14093 15895 14151 15901
rect 14093 15861 14105 15895
rect 14139 15892 14151 15895
rect 14568 15892 14596 16000
rect 20717 15997 20729 16031
rect 20763 16028 20775 16031
rect 24026 16028 24032 16040
rect 20763 16000 22140 16028
rect 23987 16000 24032 16028
rect 20763 15997 20775 16000
rect 20717 15991 20775 15997
rect 21910 15920 21916 15972
rect 21968 15960 21974 15972
rect 22112 15969 22140 16000
rect 24026 15988 24032 16000
rect 24084 16028 24090 16040
rect 25041 16031 25099 16037
rect 25041 16028 25053 16031
rect 24084 16000 25053 16028
rect 24084 15988 24090 16000
rect 25041 15997 25053 16000
rect 25087 15997 25099 16031
rect 25041 15991 25099 15997
rect 25225 16031 25283 16037
rect 25225 15997 25237 16031
rect 25271 16028 25283 16031
rect 25866 16028 25872 16040
rect 25271 16000 25872 16028
rect 25271 15997 25283 16000
rect 25225 15991 25283 15997
rect 25866 15988 25872 16000
rect 25924 15988 25930 16040
rect 22005 15963 22063 15969
rect 22005 15960 22017 15963
rect 21968 15932 22017 15960
rect 21968 15920 21974 15932
rect 22005 15929 22017 15932
rect 22051 15929 22063 15963
rect 22005 15923 22063 15929
rect 22097 15963 22155 15969
rect 22097 15929 22109 15963
rect 22143 15960 22155 15963
rect 22370 15960 22376 15972
rect 22143 15932 22376 15960
rect 22143 15929 22155 15932
rect 22097 15923 22155 15929
rect 22370 15920 22376 15932
rect 22428 15960 22434 15972
rect 22830 15960 22836 15972
rect 22428 15932 22836 15960
rect 22428 15920 22434 15932
rect 22830 15920 22836 15932
rect 22888 15920 22894 15972
rect 23474 15920 23480 15972
rect 23532 15960 23538 15972
rect 24210 15960 24216 15972
rect 23532 15932 24216 15960
rect 23532 15920 23538 15932
rect 24210 15920 24216 15932
rect 24268 15920 24274 15972
rect 15746 15892 15752 15904
rect 14139 15864 15752 15892
rect 14139 15861 14151 15864
rect 14093 15855 14151 15861
rect 15746 15852 15752 15864
rect 15804 15892 15810 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15804 15864 16221 15892
rect 15804 15852 15810 15864
rect 16209 15861 16221 15864
rect 16255 15892 16267 15895
rect 16298 15892 16304 15904
rect 16255 15864 16304 15892
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 13449 15691 13507 15697
rect 13449 15657 13461 15691
rect 13495 15688 13507 15691
rect 13538 15688 13544 15700
rect 13495 15660 13544 15688
rect 13495 15657 13507 15660
rect 13449 15651 13507 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 14277 15691 14335 15697
rect 14277 15657 14289 15691
rect 14323 15688 14335 15691
rect 14366 15688 14372 15700
rect 14323 15660 14372 15688
rect 14323 15657 14335 15660
rect 14277 15651 14335 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 16574 15648 16580 15700
rect 16632 15688 16638 15700
rect 16761 15691 16819 15697
rect 16761 15688 16773 15691
rect 16632 15660 16773 15688
rect 16632 15648 16638 15660
rect 16761 15657 16773 15660
rect 16807 15657 16819 15691
rect 21082 15688 21088 15700
rect 21043 15660 21088 15688
rect 16761 15651 16819 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 21910 15688 21916 15700
rect 21871 15660 21916 15688
rect 21910 15648 21916 15660
rect 21968 15648 21974 15700
rect 23106 15648 23112 15700
rect 23164 15688 23170 15700
rect 23937 15691 23995 15697
rect 23937 15688 23949 15691
rect 23164 15660 23949 15688
rect 23164 15648 23170 15660
rect 23937 15657 23949 15660
rect 23983 15657 23995 15691
rect 23937 15651 23995 15657
rect 24210 15648 24216 15700
rect 24268 15688 24274 15700
rect 24489 15691 24547 15697
rect 24489 15688 24501 15691
rect 24268 15660 24501 15688
rect 24268 15648 24274 15660
rect 24489 15657 24501 15660
rect 24535 15657 24547 15691
rect 25222 15688 25228 15700
rect 25183 15660 25228 15688
rect 24489 15651 24547 15657
rect 25222 15648 25228 15660
rect 25280 15648 25286 15700
rect 16482 15580 16488 15632
rect 16540 15620 16546 15632
rect 16853 15623 16911 15629
rect 16853 15620 16865 15623
rect 16540 15592 16865 15620
rect 16540 15580 16546 15592
rect 16853 15589 16865 15592
rect 16899 15620 16911 15623
rect 17126 15620 17132 15632
rect 16899 15592 17132 15620
rect 16899 15589 16911 15592
rect 16853 15583 16911 15589
rect 17126 15580 17132 15592
rect 17184 15580 17190 15632
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 17276 15592 18061 15620
rect 17276 15580 17282 15592
rect 18049 15589 18061 15592
rect 18095 15589 18107 15623
rect 18049 15583 18107 15589
rect 21545 15623 21603 15629
rect 21545 15589 21557 15623
rect 21591 15620 21603 15623
rect 22002 15620 22008 15632
rect 21591 15592 22008 15620
rect 21591 15589 21603 15592
rect 21545 15583 21603 15589
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 17770 15552 17776 15564
rect 17731 15524 17776 15552
rect 17770 15512 17776 15524
rect 17828 15512 17834 15564
rect 22830 15561 22836 15564
rect 22824 15552 22836 15561
rect 22791 15524 22836 15552
rect 22824 15515 22836 15524
rect 22830 15512 22836 15515
rect 22888 15512 22894 15564
rect 25038 15552 25044 15564
rect 24999 15524 25044 15552
rect 25038 15512 25044 15524
rect 25096 15512 25102 15564
rect 16390 15444 16396 15496
rect 16448 15484 16454 15496
rect 16758 15484 16764 15496
rect 16448 15456 16764 15484
rect 16448 15444 16454 15456
rect 16758 15444 16764 15456
rect 16816 15444 16822 15496
rect 19058 15484 19064 15496
rect 19019 15456 19064 15484
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 20990 15444 20996 15496
rect 21048 15484 21054 15496
rect 22554 15484 22560 15496
rect 21048 15456 22560 15484
rect 21048 15444 21054 15456
rect 22554 15444 22560 15456
rect 22612 15444 22618 15496
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16172 15320 16313 15348
rect 16172 15308 16178 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16301 15311 16359 15317
rect 18601 15351 18659 15357
rect 18601 15317 18613 15351
rect 18647 15348 18659 15351
rect 20162 15348 20168 15360
rect 18647 15320 20168 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 20162 15308 20168 15320
rect 20220 15308 20226 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16482 15144 16488 15156
rect 16439 15116 16488 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 16669 15147 16727 15153
rect 16669 15144 16681 15147
rect 16632 15116 16681 15144
rect 16632 15104 16638 15116
rect 16669 15113 16681 15116
rect 16715 15113 16727 15147
rect 16669 15107 16727 15113
rect 17497 15147 17555 15153
rect 17497 15113 17509 15147
rect 17543 15144 17555 15147
rect 17770 15144 17776 15156
rect 17543 15116 17776 15144
rect 17543 15113 17555 15116
rect 17497 15107 17555 15113
rect 17770 15104 17776 15116
rect 17828 15144 17834 15156
rect 18601 15147 18659 15153
rect 18601 15144 18613 15147
rect 17828 15116 18613 15144
rect 17828 15104 17834 15116
rect 18601 15113 18613 15116
rect 18647 15113 18659 15147
rect 18601 15107 18659 15113
rect 19150 15104 19156 15156
rect 19208 15144 19214 15156
rect 19889 15147 19947 15153
rect 19889 15144 19901 15147
rect 19208 15116 19901 15144
rect 19208 15104 19214 15116
rect 19889 15113 19901 15116
rect 19935 15113 19947 15147
rect 19889 15107 19947 15113
rect 21453 15147 21511 15153
rect 21453 15113 21465 15147
rect 21499 15144 21511 15147
rect 21634 15144 21640 15156
rect 21499 15116 21640 15144
rect 21499 15113 21511 15116
rect 21453 15107 21511 15113
rect 13170 15008 13176 15020
rect 13131 14980 13176 15008
rect 13170 14968 13176 14980
rect 13228 14968 13234 15020
rect 15838 15008 15844 15020
rect 15799 14980 15844 15008
rect 15838 14968 15844 14980
rect 15896 14968 15902 15020
rect 18417 15011 18475 15017
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 19058 15008 19064 15020
rect 18463 14980 19064 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 19058 14968 19064 14980
rect 19116 14968 19122 15020
rect 19904 15008 19932 15107
rect 21634 15104 21640 15116
rect 21692 15104 21698 15156
rect 22554 15144 22560 15156
rect 22515 15116 22560 15144
rect 22554 15104 22560 15116
rect 22612 15104 22618 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22888 15116 22937 15144
rect 22888 15104 22894 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 25038 15144 25044 15156
rect 24999 15116 25044 15144
rect 22925 15107 22983 15113
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19904 14980 20085 15008
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 12897 14943 12955 14949
rect 12897 14909 12909 14943
rect 12943 14940 12955 14943
rect 13633 14943 13691 14949
rect 13633 14940 13645 14943
rect 12943 14912 13645 14940
rect 12943 14909 12955 14912
rect 12897 14903 12955 14909
rect 13633 14909 13645 14912
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15488 14912 15577 14940
rect 15488 14816 15516 14912
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 19153 14875 19211 14881
rect 19153 14841 19165 14875
rect 19199 14872 19211 14875
rect 20162 14872 20168 14884
rect 19199 14844 20168 14872
rect 19199 14841 19211 14844
rect 19153 14835 19211 14841
rect 20162 14832 20168 14844
rect 20220 14872 20226 14884
rect 20340 14875 20398 14881
rect 20340 14872 20352 14875
rect 20220 14844 20352 14872
rect 20220 14832 20226 14844
rect 20340 14841 20352 14844
rect 20386 14872 20398 14875
rect 20898 14872 20904 14884
rect 20386 14844 20904 14872
rect 20386 14841 20398 14844
rect 20340 14835 20398 14841
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 15470 14804 15476 14816
rect 15431 14776 15476 14804
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 16850 14804 16856 14816
rect 16811 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 17865 14807 17923 14813
rect 17865 14773 17877 14807
rect 17911 14804 17923 14807
rect 19058 14804 19064 14816
rect 17911 14776 19064 14804
rect 17911 14773 17923 14776
rect 17865 14767 17923 14773
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 16301 14603 16359 14609
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 16390 14600 16396 14612
rect 16347 14572 16396 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21453 14603 21511 14609
rect 21453 14600 21465 14603
rect 21416 14572 21465 14600
rect 21416 14560 21422 14572
rect 21453 14569 21465 14572
rect 21499 14569 21511 14603
rect 24762 14600 24768 14612
rect 24723 14572 24768 14600
rect 21453 14563 21511 14569
rect 24762 14560 24768 14572
rect 24820 14560 24826 14612
rect 13541 14535 13599 14541
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 13630 14532 13636 14544
rect 13587 14504 13636 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 13630 14492 13636 14504
rect 13688 14532 13694 14544
rect 14185 14535 14243 14541
rect 14185 14532 14197 14535
rect 13688 14504 14197 14532
rect 13688 14492 13694 14504
rect 14185 14501 14197 14504
rect 14231 14501 14243 14535
rect 14185 14495 14243 14501
rect 16761 14535 16819 14541
rect 16761 14501 16773 14535
rect 16807 14532 16819 14535
rect 16850 14532 16856 14544
rect 16807 14504 16856 14532
rect 16807 14501 16819 14504
rect 16761 14495 16819 14501
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14464 12679 14467
rect 14001 14467 14059 14473
rect 14001 14464 14013 14467
rect 12667 14436 14013 14464
rect 12667 14433 12679 14436
rect 12621 14427 12679 14433
rect 14001 14433 14013 14436
rect 14047 14464 14059 14467
rect 14826 14464 14832 14476
rect 14047 14436 14832 14464
rect 14047 14433 14059 14436
rect 14001 14427 14059 14433
rect 14826 14424 14832 14436
rect 14884 14424 14890 14476
rect 16574 14424 16580 14476
rect 16632 14464 16638 14476
rect 16776 14464 16804 14495
rect 16850 14492 16856 14504
rect 16908 14492 16914 14544
rect 16942 14492 16948 14544
rect 17000 14532 17006 14544
rect 19150 14532 19156 14544
rect 17000 14504 17045 14532
rect 18340 14504 19156 14532
rect 17000 14492 17006 14504
rect 18340 14476 18368 14504
rect 19150 14492 19156 14504
rect 19208 14492 19214 14544
rect 21266 14532 21272 14544
rect 21227 14504 21272 14532
rect 21266 14492 21272 14504
rect 21324 14492 21330 14544
rect 18322 14464 18328 14476
rect 16632 14436 16804 14464
rect 18235 14436 18328 14464
rect 16632 14424 16638 14436
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 18598 14473 18604 14476
rect 18592 14464 18604 14473
rect 18559 14436 18604 14464
rect 18592 14427 18604 14436
rect 18598 14424 18604 14427
rect 18656 14424 18662 14476
rect 24578 14464 24584 14476
rect 24539 14436 24584 14464
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 14274 14396 14280 14408
rect 14235 14368 14280 14396
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14396 17095 14399
rect 17310 14396 17316 14408
rect 17083 14368 17316 14396
rect 17083 14365 17095 14368
rect 17037 14359 17095 14365
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 21542 14396 21548 14408
rect 21503 14368 21548 14396
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 13722 14328 13728 14340
rect 13683 14300 13728 14328
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 16485 14331 16543 14337
rect 16485 14328 16497 14331
rect 15528 14300 16497 14328
rect 15528 14288 15534 14300
rect 16485 14297 16497 14300
rect 16531 14297 16543 14331
rect 20990 14328 20996 14340
rect 20951 14300 20996 14328
rect 16485 14291 16543 14297
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 19794 14260 19800 14272
rect 19751 14232 19800 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 19794 14220 19800 14232
rect 19852 14260 19858 14272
rect 21542 14260 21548 14272
rect 19852 14232 21548 14260
rect 19852 14220 19858 14232
rect 21542 14220 21548 14232
rect 21600 14220 21606 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 12802 14056 12808 14068
rect 12763 14028 12808 14056
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14274 14056 14280 14068
rect 13872 14028 14280 14056
rect 13872 14016 13878 14028
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 14826 14056 14832 14068
rect 14787 14028 14832 14056
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 16298 14056 16304 14068
rect 15243 14028 16304 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 12820 13920 12848 14016
rect 14292 13988 14320 14016
rect 15286 13988 15292 14000
rect 14292 13960 15292 13988
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 15396 13929 15424 14028
rect 16298 14016 16304 14028
rect 16356 14056 16362 14068
rect 16850 14056 16856 14068
rect 16356 14028 16856 14056
rect 16356 14016 16362 14028
rect 16850 14016 16856 14028
rect 16908 14016 16914 14068
rect 16942 14016 16948 14068
rect 17000 14056 17006 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17000 14028 17693 14056
rect 17000 14016 17006 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 18322 14056 18328 14068
rect 18283 14028 18328 14056
rect 17681 14019 17739 14025
rect 18322 14016 18328 14028
rect 18380 14056 18386 14068
rect 19337 14059 19395 14065
rect 19337 14056 19349 14059
rect 18380 14028 19349 14056
rect 18380 14016 18386 14028
rect 19337 14025 19349 14028
rect 19383 14025 19395 14059
rect 20898 14056 20904 14068
rect 20859 14028 20904 14056
rect 19337 14019 19395 14025
rect 17310 13988 17316 14000
rect 17271 13960 17316 13988
rect 17310 13948 17316 13960
rect 17368 13988 17374 14000
rect 18230 13988 18236 14000
rect 17368 13960 18236 13988
rect 17368 13948 17374 13960
rect 18230 13948 18236 13960
rect 18288 13988 18294 14000
rect 18598 13988 18604 14000
rect 18288 13960 18604 13988
rect 18288 13948 18294 13960
rect 18598 13948 18604 13960
rect 18656 13988 18662 14000
rect 18693 13991 18751 13997
rect 18693 13988 18705 13991
rect 18656 13960 18705 13988
rect 18656 13948 18662 13960
rect 18693 13957 18705 13960
rect 18739 13957 18751 13991
rect 18693 13951 18751 13957
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12820 13892 12909 13920
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 19352 13920 19380 14019
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21266 14016 21272 14068
rect 21324 14056 21330 14068
rect 21453 14059 21511 14065
rect 21453 14056 21465 14059
rect 21324 14028 21465 14056
rect 21324 14016 21330 14028
rect 21453 14025 21465 14028
rect 21499 14025 21511 14059
rect 21453 14019 21511 14025
rect 21542 14016 21548 14068
rect 21600 14056 21606 14068
rect 21821 14059 21879 14065
rect 21821 14056 21833 14059
rect 21600 14028 21833 14056
rect 21600 14016 21606 14028
rect 21821 14025 21833 14028
rect 21867 14025 21879 14059
rect 24670 14056 24676 14068
rect 24631 14028 24676 14056
rect 21821 14019 21879 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 19352 13892 19533 13920
rect 15381 13883 15439 13889
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 16942 13852 16948 13864
rect 16500 13824 16948 13852
rect 16500 13796 16528 13824
rect 16942 13812 16948 13824
rect 17000 13812 17006 13864
rect 19610 13812 19616 13864
rect 19668 13852 19674 13864
rect 19794 13861 19800 13864
rect 19788 13852 19800 13861
rect 19668 13824 19800 13852
rect 19668 13812 19674 13824
rect 19788 13815 19800 13824
rect 19794 13812 19800 13815
rect 19852 13812 19858 13864
rect 13170 13793 13176 13796
rect 13164 13784 13176 13793
rect 13131 13756 13176 13784
rect 13164 13747 13176 13756
rect 13170 13744 13176 13747
rect 13228 13744 13234 13796
rect 15286 13744 15292 13796
rect 15344 13784 15350 13796
rect 15626 13787 15684 13793
rect 15626 13784 15638 13787
rect 15344 13756 15638 13784
rect 15344 13744 15350 13756
rect 15626 13753 15638 13756
rect 15672 13753 15684 13787
rect 15626 13747 15684 13753
rect 16482 13744 16488 13796
rect 16540 13744 16546 13796
rect 16758 13716 16764 13728
rect 16719 13688 16764 13716
rect 16758 13676 16764 13688
rect 16816 13676 16822 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 13541 13515 13599 13521
rect 13541 13481 13553 13515
rect 13587 13512 13599 13515
rect 13722 13512 13728 13524
rect 13587 13484 13728 13512
rect 13587 13481 13599 13484
rect 13541 13475 13599 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15473 13515 15531 13521
rect 15473 13512 15485 13515
rect 15344 13484 15485 13512
rect 15344 13472 15350 13484
rect 15473 13481 15485 13484
rect 15519 13481 15531 13515
rect 16390 13512 16396 13524
rect 16351 13484 16396 13512
rect 15473 13475 15531 13481
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19518 13512 19524 13524
rect 19479 13484 19524 13512
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 21174 13512 21180 13524
rect 21087 13484 21180 13512
rect 21174 13472 21180 13484
rect 21232 13512 21238 13524
rect 21358 13512 21364 13524
rect 21232 13484 21364 13512
rect 21232 13472 21238 13484
rect 21358 13472 21364 13484
rect 21416 13472 21422 13524
rect 13998 13404 14004 13456
rect 14056 13444 14062 13456
rect 14185 13447 14243 13453
rect 14185 13444 14197 13447
rect 14056 13416 14197 13444
rect 14056 13404 14062 13416
rect 14185 13413 14197 13416
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 16758 13404 16764 13456
rect 16816 13444 16822 13456
rect 17098 13447 17156 13453
rect 17098 13444 17110 13447
rect 16816 13416 17110 13444
rect 16816 13404 16822 13416
rect 17098 13413 17110 13416
rect 17144 13413 17156 13447
rect 17098 13407 17156 13413
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13170 13376 13176 13388
rect 13035 13348 13176 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 13170 13336 13176 13348
rect 13228 13376 13234 13388
rect 24578 13376 24584 13388
rect 13228 13348 14320 13376
rect 24539 13348 24584 13376
rect 13228 13336 13234 13348
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 14292 13317 14320 13348
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 16850 13308 16856 13320
rect 16811 13280 16856 13308
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 13630 13200 13636 13252
rect 13688 13240 13694 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 13688 13212 13737 13240
rect 13688 13200 13694 13212
rect 13725 13209 13737 13212
rect 13771 13209 13783 13243
rect 24762 13240 24768 13252
rect 24723 13212 24768 13240
rect 13725 13203 13783 13209
rect 24762 13200 24768 13212
rect 24820 13200 24826 13252
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 16482 12968 16488 12980
rect 16443 12940 16488 12968
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16850 12928 16856 12980
rect 16908 12968 16914 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 16908 12940 17417 12968
rect 16908 12928 16914 12940
rect 17405 12937 17417 12940
rect 17451 12937 17463 12971
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 17405 12931 17463 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12860 12804 13093 12832
rect 12860 12792 12866 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16666 12832 16672 12844
rect 16347 12804 16672 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16816 12804 17049 12832
rect 16816 12792 16822 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 16776 12764 16804 12792
rect 15979 12736 16804 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 13354 12705 13360 12708
rect 12989 12699 13047 12705
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 13348 12696 13360 12705
rect 13035 12668 13360 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 13348 12659 13360 12668
rect 13354 12656 13360 12659
rect 13412 12656 13418 12708
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 16724 12668 16773 12696
rect 16724 12656 16730 12668
rect 16761 12665 16773 12668
rect 16807 12696 16819 12699
rect 16850 12696 16856 12708
rect 16807 12668 16856 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 16942 12656 16948 12708
rect 17000 12696 17006 12708
rect 17000 12668 17045 12696
rect 17000 12656 17006 12668
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16960 12628 16988 12656
rect 16632 12600 16988 12628
rect 16632 12588 16638 12600
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12860 12396 13093 12424
rect 12860 12384 12866 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 13725 12427 13783 12433
rect 13725 12393 13737 12427
rect 13771 12424 13783 12427
rect 14182 12424 14188 12436
rect 13771 12396 14188 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 14458 12424 14464 12436
rect 14419 12396 14464 12424
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 16758 12384 16764 12436
rect 16816 12424 16822 12436
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 16816 12396 16865 12424
rect 16816 12384 16822 12396
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 16853 12387 16911 12393
rect 24765 12427 24823 12433
rect 24765 12393 24777 12427
rect 24811 12424 24823 12427
rect 25314 12424 25320 12436
rect 24811 12396 25320 12424
rect 24811 12393 24823 12396
rect 24765 12387 24823 12393
rect 25314 12384 25320 12396
rect 25372 12384 25378 12436
rect 13998 12356 14004 12368
rect 13959 12328 14004 12356
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 16393 12359 16451 12365
rect 16393 12356 16405 12359
rect 14056 12328 16405 12356
rect 14056 12316 14062 12328
rect 16393 12325 16405 12328
rect 16439 12356 16451 12359
rect 16482 12356 16488 12368
rect 16439 12328 16488 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 24578 12288 24584 12300
rect 24539 12260 24584 12288
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 13262 11880 13268 11892
rect 13223 11852 13268 11880
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 24670 11880 24676 11892
rect 24631 11852 24676 11880
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 12713 11679 12771 11685
rect 12713 11645 12725 11679
rect 12759 11676 12771 11679
rect 13262 11676 13268 11688
rect 12759 11648 13268 11676
rect 12759 11645 12771 11648
rect 12713 11639 12771 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 12066 11200 12072 11212
rect 12027 11172 12072 11200
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 12250 11064 12256 11076
rect 12211 11036 12256 11064
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11664 10764 11805 10792
rect 11664 10752 11670 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12124 10764 12173 10792
rect 12124 10752 12130 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10588 11299 10591
rect 11606 10588 11612 10600
rect 11287 10560 11612 10588
rect 11287 10557 11299 10560
rect 11241 10551 11299 10557
rect 11606 10548 11612 10560
rect 11664 10548 11670 10600
rect 11422 10452 11428 10464
rect 11383 10424 11428 10452
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 9858 10072 9864 10124
rect 9916 10112 9922 10124
rect 10689 10115 10747 10121
rect 10689 10112 10701 10115
rect 9916 10084 10701 10112
rect 9916 10072 9922 10084
rect 10689 10081 10701 10084
rect 10735 10112 10747 10115
rect 10962 10112 10968 10124
rect 10735 10084 10968 10112
rect 10735 10081 10747 10084
rect 10689 10075 10747 10081
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 10870 9976 10876 9988
rect 10831 9948 10876 9976
rect 10870 9936 10876 9948
rect 10928 9936 10934 9988
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 10962 9704 10968 9716
rect 10923 9676 10968 9704
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 10226 9636 10232 9648
rect 10187 9608 10232 9636
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9824 9472 10057 9500
rect 9824 9460 9830 9472
rect 10045 9469 10057 9472
rect 10091 9500 10103 9503
rect 10597 9503 10655 9509
rect 10597 9500 10609 9503
rect 10091 9472 10609 9500
rect 10091 9469 10103 9472
rect 10045 9463 10103 9469
rect 10597 9469 10609 9472
rect 10643 9469 10655 9503
rect 24578 9500 24584 9512
rect 24491 9472 24584 9500
rect 10597 9463 10655 9469
rect 24578 9460 24584 9472
rect 24636 9500 24642 9512
rect 25133 9503 25191 9509
rect 25133 9500 25145 9503
rect 24636 9472 25145 9500
rect 24636 9460 24642 9472
rect 25133 9469 25145 9472
rect 25179 9469 25191 9503
rect 25133 9463 25191 9469
rect 24762 9364 24768 9376
rect 24723 9336 24768 9364
rect 24762 9324 24768 9336
rect 24820 9324 24826 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 24578 9092 24584 9104
rect 24539 9064 24584 9092
rect 24578 9052 24584 9064
rect 24636 9052 24642 9104
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 23658 8984 23664 9036
rect 23716 9024 23722 9036
rect 24305 9027 24363 9033
rect 24305 9024 24317 9027
rect 23716 8996 24317 9024
rect 23716 8984 23722 8996
rect 24305 8993 24317 8996
rect 24351 9024 24363 9027
rect 24946 9024 24952 9036
rect 24351 8996 24952 9024
rect 24351 8993 24363 8996
rect 24305 8987 24363 8993
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 9858 8888 9864 8900
rect 9819 8860 9864 8888
rect 9858 8848 9864 8860
rect 9916 8848 9922 8900
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 9674 8616 9680 8628
rect 9635 8588 9680 8616
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 25314 8548 25320 8560
rect 25275 8520 25320 8548
rect 25314 8508 25320 8520
rect 25372 8508 25378 8560
rect 24581 8483 24639 8489
rect 24581 8480 24593 8483
rect 23860 8452 24593 8480
rect 23860 8424 23888 8452
rect 24581 8449 24593 8452
rect 24627 8449 24639 8483
rect 24581 8443 24639 8449
rect 23842 8412 23848 8424
rect 23803 8384 23848 8412
rect 23842 8372 23848 8384
rect 23900 8372 23906 8424
rect 24121 8415 24179 8421
rect 24121 8381 24133 8415
rect 24167 8412 24179 8415
rect 25133 8415 25191 8421
rect 25133 8412 25145 8415
rect 24167 8384 25145 8412
rect 24167 8381 24179 8384
rect 24121 8375 24179 8381
rect 25133 8381 25145 8384
rect 25179 8412 25191 8415
rect 25685 8415 25743 8421
rect 25685 8412 25697 8415
rect 25179 8384 25697 8412
rect 25179 8381 25191 8384
rect 25133 8375 25191 8381
rect 25685 8381 25697 8384
rect 25731 8381 25743 8415
rect 25685 8375 25743 8381
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 19334 7936 19340 7948
rect 19295 7908 19340 7936
rect 19334 7896 19340 7908
rect 19392 7896 19398 7948
rect 21818 7896 21824 7948
rect 21876 7936 21882 7948
rect 22922 7936 22928 7948
rect 21876 7908 22928 7936
rect 21876 7896 21882 7908
rect 22922 7896 22928 7908
rect 22980 7896 22986 7948
rect 23201 7939 23259 7945
rect 23201 7905 23213 7939
rect 23247 7936 23259 7939
rect 24210 7936 24216 7948
rect 23247 7908 24216 7936
rect 23247 7905 23259 7908
rect 23201 7899 23259 7905
rect 24210 7896 24216 7908
rect 24268 7936 24274 7948
rect 24305 7939 24363 7945
rect 24305 7936 24317 7939
rect 24268 7908 24317 7936
rect 24268 7896 24274 7908
rect 24305 7905 24317 7908
rect 24351 7905 24363 7939
rect 24305 7899 24363 7905
rect 19610 7868 19616 7880
rect 19571 7840 19616 7868
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 24489 7735 24547 7741
rect 24489 7701 24501 7735
rect 24535 7732 24547 7735
rect 24762 7732 24768 7744
rect 24535 7704 24768 7732
rect 24535 7701 24547 7704
rect 24489 7695 24547 7701
rect 24762 7692 24768 7704
rect 24820 7692 24826 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 19334 7528 19340 7540
rect 19295 7500 19340 7528
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 22922 7528 22928 7540
rect 22883 7500 22928 7528
rect 22922 7488 22928 7500
rect 22980 7488 22986 7540
rect 24210 7488 24216 7540
rect 24268 7528 24274 7540
rect 24305 7531 24363 7537
rect 24305 7528 24317 7531
rect 24268 7500 24317 7528
rect 24268 7488 24274 7500
rect 24305 7497 24317 7500
rect 24351 7497 24363 7531
rect 24305 7491 24363 7497
rect 24578 7324 24584 7336
rect 24539 7296 24584 7324
rect 24578 7284 24584 7296
rect 24636 7324 24642 7336
rect 25133 7327 25191 7333
rect 25133 7324 25145 7327
rect 24636 7296 25145 7324
rect 24636 7284 24642 7296
rect 25133 7293 25145 7296
rect 25179 7293 25191 7327
rect 25133 7287 25191 7293
rect 24670 7148 24676 7200
rect 24728 7188 24734 7200
rect 24765 7191 24823 7197
rect 24765 7188 24777 7191
rect 24728 7160 24777 7188
rect 24728 7148 24734 7160
rect 24765 7157 24777 7160
rect 24811 7157 24823 7191
rect 24765 7151 24823 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 23474 6808 23480 6860
rect 23532 6848 23538 6860
rect 23661 6851 23719 6857
rect 23661 6848 23673 6851
rect 23532 6820 23673 6848
rect 23532 6808 23538 6820
rect 23661 6817 23673 6820
rect 23707 6817 23719 6851
rect 23661 6811 23719 6817
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24762 6848 24768 6860
rect 23983 6820 24768 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24762 6808 24768 6820
rect 24820 6848 24826 6860
rect 24949 6851 25007 6857
rect 24949 6848 24961 6851
rect 24820 6820 24961 6848
rect 24820 6808 24826 6820
rect 24949 6817 24961 6820
rect 24995 6817 25007 6851
rect 24949 6811 25007 6817
rect 25130 6644 25136 6656
rect 25091 6616 25136 6644
rect 25130 6604 25136 6616
rect 25188 6604 25194 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 23474 6440 23480 6452
rect 23435 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 24762 6440 24768 6452
rect 24723 6412 24768 6440
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14608 6208 14933 6236
rect 14608 6196 14614 6208
rect 14921 6205 14933 6208
rect 14967 6236 14979 6239
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 14967 6208 15669 6236
rect 14967 6205 14979 6208
rect 14921 6199 14979 6205
rect 15657 6205 15669 6208
rect 15703 6205 15715 6239
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 15657 6199 15715 6205
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 23937 6239 23995 6245
rect 23937 6205 23949 6239
rect 23983 6236 23995 6239
rect 24949 6239 25007 6245
rect 24949 6236 24961 6239
rect 23983 6208 24961 6236
rect 23983 6205 23995 6208
rect 23937 6199 23995 6205
rect 24949 6205 24961 6208
rect 24995 6236 25007 6239
rect 25501 6239 25559 6245
rect 25501 6236 25513 6239
rect 24995 6208 25513 6236
rect 24995 6205 25007 6208
rect 24949 6199 25007 6205
rect 25501 6205 25513 6208
rect 25547 6205 25559 6239
rect 25501 6199 25559 6205
rect 15194 6168 15200 6180
rect 15155 6140 15200 6168
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 23676 6168 23704 6196
rect 24397 6171 24455 6177
rect 24397 6168 24409 6171
rect 23676 6140 24409 6168
rect 24397 6137 24409 6140
rect 24443 6137 24455 6171
rect 24397 6131 24455 6137
rect 25133 6103 25191 6109
rect 25133 6069 25145 6103
rect 25179 6100 25191 6103
rect 26142 6100 26148 6112
rect 25179 6072 26148 6100
rect 25179 6069 25191 6072
rect 25133 6063 25191 6069
rect 26142 6060 26148 6072
rect 26200 6060 26206 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 23658 5760 23664 5772
rect 23619 5732 23664 5760
rect 23658 5720 23664 5732
rect 23716 5720 23722 5772
rect 24946 5760 24952 5772
rect 24907 5732 24952 5760
rect 24946 5720 24952 5732
rect 25004 5720 25010 5772
rect 23842 5692 23848 5704
rect 23803 5664 23848 5692
rect 23842 5652 23848 5664
rect 23900 5652 23906 5704
rect 25130 5556 25136 5568
rect 25091 5528 25136 5556
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 23477 5355 23535 5361
rect 23477 5321 23489 5355
rect 23523 5352 23535 5355
rect 23658 5352 23664 5364
rect 23523 5324 23664 5352
rect 23523 5321 23535 5324
rect 23477 5315 23535 5321
rect 23658 5312 23664 5324
rect 23716 5312 23722 5364
rect 24857 5355 24915 5361
rect 24857 5321 24869 5355
rect 24903 5352 24915 5355
rect 24946 5352 24952 5364
rect 24903 5324 24952 5352
rect 24903 5321 24915 5324
rect 24857 5315 24915 5321
rect 24946 5312 24952 5324
rect 25004 5312 25010 5364
rect 23658 5148 23664 5160
rect 23619 5120 23664 5148
rect 23658 5108 23664 5120
rect 23716 5148 23722 5160
rect 24397 5151 24455 5157
rect 24397 5148 24409 5151
rect 23716 5120 24409 5148
rect 23716 5108 23722 5120
rect 24397 5117 24409 5120
rect 24443 5117 24455 5151
rect 24397 5111 24455 5117
rect 24949 5151 25007 5157
rect 24949 5117 24961 5151
rect 24995 5117 25007 5151
rect 24949 5111 25007 5117
rect 23937 5083 23995 5089
rect 23937 5049 23949 5083
rect 23983 5080 23995 5083
rect 24964 5080 24992 5111
rect 25501 5083 25559 5089
rect 25501 5080 25513 5083
rect 23983 5052 25513 5080
rect 23983 5049 23995 5052
rect 23937 5043 23995 5049
rect 25501 5049 25513 5052
rect 25547 5049 25559 5083
rect 25501 5043 25559 5049
rect 25130 5012 25136 5024
rect 25091 4984 25136 5012
rect 25130 4972 25136 4984
rect 25188 4972 25194 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 23477 4675 23535 4681
rect 23477 4641 23489 4675
rect 23523 4672 23535 4675
rect 23842 4672 23848 4684
rect 23523 4644 23848 4672
rect 23523 4641 23535 4644
rect 23477 4635 23535 4641
rect 23842 4632 23848 4644
rect 23900 4632 23906 4684
rect 24210 4632 24216 4684
rect 24268 4672 24274 4684
rect 24581 4675 24639 4681
rect 24581 4672 24593 4675
rect 24268 4644 24593 4672
rect 24268 4632 24274 4644
rect 24581 4641 24593 4644
rect 24627 4641 24639 4675
rect 24581 4635 24639 4641
rect 23661 4471 23719 4477
rect 23661 4437 23673 4471
rect 23707 4468 23719 4471
rect 24670 4468 24676 4480
rect 23707 4440 24676 4468
rect 23707 4437 23719 4440
rect 23661 4431 23719 4437
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 24820 4440 24865 4468
rect 24820 4428 24826 4440
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 23842 4264 23848 4276
rect 23803 4236 23848 4264
rect 23842 4224 23848 4236
rect 23900 4224 23906 4276
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24581 4063 24639 4069
rect 24581 4060 24593 4063
rect 23992 4032 24593 4060
rect 23992 4020 23998 4032
rect 24581 4029 24593 4032
rect 24627 4060 24639 4063
rect 25133 4063 25191 4069
rect 25133 4060 25145 4063
rect 24627 4032 25145 4060
rect 24627 4029 24639 4032
rect 24581 4023 24639 4029
rect 25133 4029 25145 4032
rect 25179 4029 25191 4063
rect 25133 4023 25191 4029
rect 24210 3952 24216 4004
rect 24268 3992 24274 4004
rect 24268 3964 24808 3992
rect 24268 3952 24274 3964
rect 24394 3924 24400 3936
rect 24355 3896 24400 3924
rect 24394 3884 24400 3896
rect 24452 3884 24458 3936
rect 24780 3933 24808 3964
rect 24765 3927 24823 3933
rect 24765 3893 24777 3927
rect 24811 3893 24823 3927
rect 24765 3887 24823 3893
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 23753 3655 23811 3661
rect 23753 3621 23765 3655
rect 23799 3652 23811 3655
rect 24394 3652 24400 3664
rect 23799 3624 24400 3652
rect 23799 3621 23811 3624
rect 23753 3615 23811 3621
rect 24394 3612 24400 3624
rect 24452 3612 24458 3664
rect 23474 3584 23480 3596
rect 23435 3556 23480 3584
rect 23474 3544 23480 3556
rect 23532 3544 23538 3596
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3584 24823 3587
rect 24854 3584 24860 3596
rect 24811 3556 24860 3584
rect 24811 3553 24823 3556
rect 24765 3547 24823 3553
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 24762 3340 24768 3392
rect 24820 3380 24826 3392
rect 24949 3383 25007 3389
rect 24949 3380 24961 3383
rect 24820 3352 24961 3380
rect 24820 3340 24826 3352
rect 24949 3349 24961 3352
rect 24995 3349 25007 3383
rect 24949 3343 25007 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 23109 3179 23167 3185
rect 23109 3145 23121 3179
rect 23155 3176 23167 3179
rect 23750 3176 23756 3188
rect 23155 3148 23756 3176
rect 23155 3145 23167 3148
rect 23109 3139 23167 3145
rect 22281 2975 22339 2981
rect 22281 2941 22293 2975
rect 22327 2972 22339 2975
rect 23124 2972 23152 3139
rect 23750 3136 23756 3148
rect 23808 3136 23814 3188
rect 24854 3176 24860 3188
rect 24815 3148 24860 3176
rect 24854 3136 24860 3148
rect 24912 3136 24918 3188
rect 23474 3108 23480 3120
rect 23435 3080 23480 3108
rect 23474 3068 23480 3080
rect 23532 3068 23538 3120
rect 23934 3040 23940 3052
rect 23895 3012 23940 3040
rect 23934 3000 23940 3012
rect 23992 3000 23998 3052
rect 24872 3040 24900 3136
rect 25133 3043 25191 3049
rect 25133 3040 25145 3043
rect 24872 3012 25145 3040
rect 25133 3009 25145 3012
rect 25179 3009 25191 3043
rect 25133 3003 25191 3009
rect 23658 2972 23664 2984
rect 22327 2944 23152 2972
rect 23619 2944 23664 2972
rect 22327 2941 22339 2944
rect 22281 2935 22339 2941
rect 23658 2932 23664 2944
rect 23716 2972 23722 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 23716 2944 24409 2972
rect 23716 2932 23722 2944
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 24946 2972 24952 2984
rect 24907 2944 24952 2972
rect 24397 2935 24455 2941
rect 24946 2932 24952 2944
rect 25004 2972 25010 2984
rect 25685 2975 25743 2981
rect 25685 2972 25697 2975
rect 25004 2944 25697 2972
rect 25004 2932 25010 2944
rect 25685 2941 25697 2944
rect 25731 2941 25743 2975
rect 25685 2935 25743 2941
rect 22554 2904 22560 2916
rect 22515 2876 22560 2904
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 22833 2499 22891 2505
rect 22833 2465 22845 2499
rect 22879 2496 22891 2499
rect 24026 2496 24032 2508
rect 22879 2468 23520 2496
rect 23987 2468 24032 2496
rect 22879 2465 22891 2468
rect 22833 2459 22891 2465
rect 23492 2437 23520 2468
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24084 2468 24777 2496
rect 24084 2456 24090 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 25314 2496 25320 2508
rect 25275 2468 25320 2496
rect 24765 2459 24823 2465
rect 25314 2456 25320 2468
rect 25372 2496 25378 2508
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25372 2468 25881 2496
rect 25372 2456 25378 2468
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2428 23535 2431
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 23523 2400 24225 2428
rect 23523 2397 23535 2400
rect 23477 2391 23535 2397
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 23014 2292 23020 2304
rect 22975 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2252 23078 2304
rect 25498 2292 25504 2304
rect 25459 2264 25504 2292
rect 25498 2252 25504 2264
rect 25556 2252 25562 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 20352 26936 20404 26988
rect 24768 26936 24820 26988
rect 19984 26392 20036 26444
rect 24768 26392 24820 26444
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 21548 25440 21600 25492
rect 23572 25440 23624 25492
rect 18696 25372 18748 25424
rect 23204 25304 23256 25356
rect 24768 25304 24820 25356
rect 19432 25279 19484 25288
rect 19432 25245 19441 25279
rect 19441 25245 19475 25279
rect 19475 25245 19484 25279
rect 19432 25236 19484 25245
rect 19616 25236 19668 25288
rect 14832 25100 14884 25152
rect 19340 25100 19392 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 19432 24896 19484 24948
rect 23664 24896 23716 24948
rect 24768 24896 24820 24948
rect 9680 24760 9732 24812
rect 10140 24760 10192 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 19616 24828 19668 24880
rect 20076 24828 20128 24880
rect 14372 24692 14424 24744
rect 18696 24692 18748 24744
rect 14004 24667 14056 24676
rect 14004 24633 14013 24667
rect 14013 24633 14047 24667
rect 14047 24633 14056 24667
rect 14004 24624 14056 24633
rect 14464 24624 14516 24676
rect 18512 24556 18564 24608
rect 19708 24624 19760 24676
rect 20168 24624 20220 24676
rect 19156 24599 19208 24608
rect 19156 24565 19165 24599
rect 19165 24565 19199 24599
rect 19199 24565 19208 24599
rect 19156 24556 19208 24565
rect 24676 24828 24728 24880
rect 22376 24599 22428 24608
rect 22376 24565 22385 24599
rect 22385 24565 22419 24599
rect 22419 24565 22428 24599
rect 22376 24556 22428 24565
rect 22928 24556 22980 24608
rect 23204 24556 23256 24608
rect 24032 24556 24084 24608
rect 24216 24624 24268 24676
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 14280 24352 14332 24404
rect 14832 24352 14884 24404
rect 15568 24352 15620 24404
rect 20260 24352 20312 24404
rect 25412 24395 25464 24404
rect 25412 24361 25421 24395
rect 25421 24361 25455 24395
rect 25455 24361 25464 24395
rect 25412 24352 25464 24361
rect 18604 24284 18656 24336
rect 10324 24216 10376 24268
rect 11244 24216 11296 24268
rect 11060 24148 11112 24200
rect 10784 24012 10836 24064
rect 11428 24012 11480 24064
rect 12532 24055 12584 24064
rect 12532 24021 12541 24055
rect 12541 24021 12575 24055
rect 12575 24021 12584 24055
rect 12532 24012 12584 24021
rect 13176 24012 13228 24064
rect 15844 24216 15896 24268
rect 21364 24216 21416 24268
rect 23020 24259 23072 24268
rect 23020 24225 23054 24259
rect 23054 24225 23072 24259
rect 25228 24259 25280 24268
rect 23020 24216 23072 24225
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 22744 24191 22796 24200
rect 18696 24123 18748 24132
rect 18696 24089 18705 24123
rect 18705 24089 18739 24123
rect 18739 24089 18748 24123
rect 18696 24080 18748 24089
rect 14372 24012 14424 24064
rect 19616 24012 19668 24064
rect 22744 24157 22753 24191
rect 22753 24157 22787 24191
rect 22787 24157 22796 24191
rect 22744 24148 22796 24157
rect 20168 24012 20220 24064
rect 24124 24055 24176 24064
rect 24124 24021 24133 24055
rect 24133 24021 24167 24055
rect 24167 24021 24176 24055
rect 24124 24012 24176 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 11244 23808 11296 23860
rect 16856 23851 16908 23860
rect 9864 23740 9916 23792
rect 11428 23715 11480 23724
rect 11428 23681 11437 23715
rect 11437 23681 11471 23715
rect 11471 23681 11480 23715
rect 11428 23672 11480 23681
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 16856 23817 16865 23851
rect 16865 23817 16899 23851
rect 16899 23817 16908 23851
rect 16856 23808 16908 23817
rect 20904 23808 20956 23860
rect 22744 23851 22796 23860
rect 22744 23817 22753 23851
rect 22753 23817 22787 23851
rect 22787 23817 22796 23851
rect 22744 23808 22796 23817
rect 23020 23808 23072 23860
rect 23388 23808 23440 23860
rect 24676 23808 24728 23860
rect 17776 23740 17828 23792
rect 18236 23672 18288 23724
rect 12164 23647 12216 23656
rect 10784 23468 10836 23520
rect 12164 23613 12173 23647
rect 12173 23613 12207 23647
rect 12207 23613 12216 23647
rect 12164 23604 12216 23613
rect 11428 23468 11480 23520
rect 12440 23468 12492 23520
rect 13820 23468 13872 23520
rect 14280 23604 14332 23656
rect 14832 23604 14884 23656
rect 18604 23647 18656 23656
rect 18604 23613 18613 23647
rect 18613 23613 18647 23647
rect 18647 23613 18656 23647
rect 18604 23604 18656 23613
rect 19156 23604 19208 23656
rect 20536 23740 20588 23792
rect 24676 23672 24728 23724
rect 25228 23672 25280 23724
rect 19616 23647 19668 23656
rect 18696 23536 18748 23588
rect 19616 23613 19650 23647
rect 19650 23613 19668 23647
rect 19616 23604 19668 23613
rect 23296 23536 23348 23588
rect 14188 23468 14240 23520
rect 14740 23468 14792 23520
rect 15292 23468 15344 23520
rect 15844 23468 15896 23520
rect 17224 23511 17276 23520
rect 17224 23477 17233 23511
rect 17233 23477 17267 23511
rect 17267 23477 17276 23511
rect 17224 23468 17276 23477
rect 19064 23468 19116 23520
rect 20720 23511 20772 23520
rect 20720 23477 20729 23511
rect 20729 23477 20763 23511
rect 20763 23477 20772 23511
rect 20720 23468 20772 23477
rect 21364 23511 21416 23520
rect 21364 23477 21373 23511
rect 21373 23477 21407 23511
rect 21407 23477 21416 23511
rect 21364 23468 21416 23477
rect 25228 23511 25280 23520
rect 25228 23477 25237 23511
rect 25237 23477 25271 23511
rect 25271 23477 25280 23511
rect 25228 23468 25280 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 10968 23264 11020 23316
rect 11244 23264 11296 23316
rect 14280 23264 14332 23316
rect 18696 23307 18748 23316
rect 18696 23273 18705 23307
rect 18705 23273 18739 23307
rect 18739 23273 18748 23307
rect 18696 23264 18748 23273
rect 10140 23060 10192 23112
rect 11428 23196 11480 23248
rect 12532 23196 12584 23248
rect 13084 23196 13136 23248
rect 10968 23128 11020 23180
rect 12440 23060 12492 23112
rect 13728 23128 13780 23180
rect 17776 23196 17828 23248
rect 18972 23196 19024 23248
rect 20352 23264 20404 23316
rect 22008 23264 22060 23316
rect 23480 23264 23532 23316
rect 19892 23239 19944 23248
rect 19892 23205 19901 23239
rect 19901 23205 19935 23239
rect 19935 23205 19944 23239
rect 19892 23196 19944 23205
rect 20076 23196 20128 23248
rect 20628 23196 20680 23248
rect 22928 23196 22980 23248
rect 23572 23196 23624 23248
rect 16948 23171 17000 23180
rect 16948 23137 16982 23171
rect 16982 23137 17000 23171
rect 16948 23128 17000 23137
rect 19524 23128 19576 23180
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 22836 23171 22888 23180
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 23848 23128 23900 23180
rect 14740 23060 14792 23112
rect 22284 23060 22336 23112
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 12992 22924 13044 22976
rect 13728 22924 13780 22976
rect 17316 22924 17368 22976
rect 19340 22967 19392 22976
rect 19340 22933 19349 22967
rect 19349 22933 19383 22967
rect 19383 22933 19392 22967
rect 19340 22924 19392 22933
rect 22560 22967 22612 22976
rect 22560 22933 22569 22967
rect 22569 22933 22603 22967
rect 22603 22933 22612 22967
rect 22560 22924 22612 22933
rect 23940 22924 23992 22976
rect 24124 22967 24176 22976
rect 24124 22933 24133 22967
rect 24133 22933 24167 22967
rect 24167 22933 24176 22967
rect 24124 22924 24176 22933
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10968 22763 11020 22772
rect 10968 22729 10977 22763
rect 10977 22729 11011 22763
rect 11011 22729 11020 22763
rect 10968 22720 11020 22729
rect 12440 22720 12492 22772
rect 13084 22763 13136 22772
rect 13084 22729 13093 22763
rect 13093 22729 13127 22763
rect 13127 22729 13136 22763
rect 13084 22720 13136 22729
rect 16948 22720 17000 22772
rect 17960 22720 18012 22772
rect 19892 22720 19944 22772
rect 22284 22720 22336 22772
rect 22928 22720 22980 22772
rect 23480 22763 23532 22772
rect 23480 22729 23489 22763
rect 23489 22729 23523 22763
rect 23523 22729 23532 22763
rect 23480 22720 23532 22729
rect 14556 22652 14608 22704
rect 16580 22652 16632 22704
rect 17500 22695 17552 22704
rect 17500 22661 17509 22695
rect 17509 22661 17543 22695
rect 17543 22661 17552 22695
rect 17500 22652 17552 22661
rect 17776 22652 17828 22704
rect 22100 22695 22152 22704
rect 22100 22661 22109 22695
rect 22109 22661 22143 22695
rect 22143 22661 22152 22695
rect 22100 22652 22152 22661
rect 23388 22652 23440 22704
rect 23756 22695 23808 22704
rect 23756 22661 23765 22695
rect 23765 22661 23799 22695
rect 23799 22661 23808 22695
rect 23756 22652 23808 22661
rect 14740 22627 14792 22636
rect 14740 22593 14749 22627
rect 14749 22593 14783 22627
rect 14783 22593 14792 22627
rect 14740 22584 14792 22593
rect 14648 22516 14700 22568
rect 15108 22584 15160 22636
rect 21824 22627 21876 22636
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 16856 22516 16908 22568
rect 14464 22448 14516 22500
rect 16120 22448 16172 22500
rect 10140 22380 10192 22432
rect 10692 22380 10744 22432
rect 17316 22448 17368 22500
rect 20536 22516 20588 22568
rect 18972 22423 19024 22432
rect 18972 22389 18981 22423
rect 18981 22389 19015 22423
rect 19015 22389 19024 22423
rect 18972 22380 19024 22389
rect 19892 22448 19944 22500
rect 22468 22448 22520 22500
rect 23572 22584 23624 22636
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 25596 22720 25648 22772
rect 24492 22584 24544 22636
rect 23848 22516 23900 22568
rect 23112 22448 23164 22500
rect 23940 22448 23992 22500
rect 25872 22491 25924 22500
rect 25872 22457 25881 22491
rect 25881 22457 25915 22491
rect 25915 22457 25924 22491
rect 25872 22448 25924 22457
rect 20628 22380 20680 22432
rect 23480 22380 23532 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 9956 22176 10008 22228
rect 14464 22176 14516 22228
rect 17408 22176 17460 22228
rect 19524 22176 19576 22228
rect 20904 22176 20956 22228
rect 23020 22176 23072 22228
rect 23664 22176 23716 22228
rect 24492 22176 24544 22228
rect 13636 22040 13688 22092
rect 16856 22108 16908 22160
rect 17040 22083 17092 22092
rect 17040 22049 17049 22083
rect 17049 22049 17083 22083
rect 17083 22049 17092 22083
rect 17040 22040 17092 22049
rect 17776 22040 17828 22092
rect 19984 22108 20036 22160
rect 22100 22108 22152 22160
rect 23296 22108 23348 22160
rect 22468 22040 22520 22092
rect 22560 22040 22612 22092
rect 23020 22083 23072 22092
rect 23020 22049 23029 22083
rect 23029 22049 23063 22083
rect 23063 22049 23072 22083
rect 24216 22083 24268 22092
rect 23020 22040 23072 22049
rect 24216 22049 24239 22083
rect 24239 22049 24268 22083
rect 24216 22040 24268 22049
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 14096 22015 14148 22024
rect 14096 21981 14105 22015
rect 14105 21981 14139 22015
rect 14139 21981 14148 22015
rect 14096 21972 14148 21981
rect 14280 22015 14332 22024
rect 14280 21981 14289 22015
rect 14289 21981 14323 22015
rect 14323 21981 14332 22015
rect 14280 21972 14332 21981
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 18880 22015 18932 22024
rect 18880 21981 18889 22015
rect 18889 21981 18923 22015
rect 18923 21981 18932 22015
rect 18880 21972 18932 21981
rect 22836 21972 22888 22024
rect 22928 21972 22980 22024
rect 23480 21904 23532 21956
rect 23664 21904 23716 21956
rect 10876 21836 10928 21888
rect 13728 21879 13780 21888
rect 13728 21845 13737 21879
rect 13737 21845 13771 21879
rect 13771 21845 13780 21879
rect 13728 21836 13780 21845
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 21732 21879 21784 21888
rect 21732 21845 21741 21879
rect 21741 21845 21775 21879
rect 21775 21845 21784 21879
rect 21732 21836 21784 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10784 21632 10836 21684
rect 13636 21675 13688 21684
rect 13636 21641 13645 21675
rect 13645 21641 13679 21675
rect 13679 21641 13688 21675
rect 13636 21632 13688 21641
rect 15568 21632 15620 21684
rect 16580 21632 16632 21684
rect 17776 21675 17828 21684
rect 17776 21641 17785 21675
rect 17785 21641 17819 21675
rect 17819 21641 17828 21675
rect 17776 21632 17828 21641
rect 18880 21632 18932 21684
rect 22008 21632 22060 21684
rect 23572 21632 23624 21684
rect 10048 21564 10100 21616
rect 14280 21564 14332 21616
rect 16764 21607 16816 21616
rect 16764 21573 16773 21607
rect 16773 21573 16807 21607
rect 16807 21573 16816 21607
rect 16764 21564 16816 21573
rect 17040 21607 17092 21616
rect 17040 21573 17049 21607
rect 17049 21573 17083 21607
rect 17083 21573 17092 21607
rect 17040 21564 17092 21573
rect 19248 21607 19300 21616
rect 19248 21573 19257 21607
rect 19257 21573 19291 21607
rect 19291 21573 19300 21607
rect 19248 21564 19300 21573
rect 23112 21607 23164 21616
rect 23112 21573 23121 21607
rect 23121 21573 23155 21607
rect 23155 21573 23164 21607
rect 23112 21564 23164 21573
rect 9956 21496 10008 21548
rect 10968 21539 11020 21548
rect 10968 21505 10977 21539
rect 10977 21505 11011 21539
rect 11011 21505 11020 21539
rect 10968 21496 11020 21505
rect 13820 21496 13872 21548
rect 14096 21496 14148 21548
rect 17960 21496 18012 21548
rect 20628 21496 20680 21548
rect 22468 21496 22520 21548
rect 23020 21496 23072 21548
rect 10692 21471 10744 21480
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 10876 21403 10928 21412
rect 10876 21369 10885 21403
rect 10885 21369 10919 21403
rect 10919 21369 10928 21403
rect 10876 21360 10928 21369
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 14004 21292 14056 21344
rect 14648 21471 14700 21480
rect 14648 21437 14682 21471
rect 14682 21437 14700 21471
rect 14648 21428 14700 21437
rect 19340 21428 19392 21480
rect 22928 21428 22980 21480
rect 23204 21428 23256 21480
rect 23388 21428 23440 21480
rect 23664 21471 23716 21480
rect 23664 21437 23673 21471
rect 23673 21437 23707 21471
rect 23707 21437 23716 21471
rect 23664 21428 23716 21437
rect 19432 21360 19484 21412
rect 23112 21360 23164 21412
rect 17316 21292 17368 21344
rect 17776 21292 17828 21344
rect 17960 21292 18012 21344
rect 21732 21292 21784 21344
rect 22744 21292 22796 21344
rect 24216 21292 24268 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 10968 21088 11020 21140
rect 13636 21088 13688 21140
rect 13912 21088 13964 21140
rect 14648 21088 14700 21140
rect 16488 21131 16540 21140
rect 16488 21097 16497 21131
rect 16497 21097 16531 21131
rect 16531 21097 16540 21131
rect 16488 21088 16540 21097
rect 18880 21131 18932 21140
rect 18880 21097 18889 21131
rect 18889 21097 18923 21131
rect 18923 21097 18932 21131
rect 18880 21088 18932 21097
rect 19432 21131 19484 21140
rect 19432 21097 19441 21131
rect 19441 21097 19475 21131
rect 19475 21097 19484 21131
rect 19432 21088 19484 21097
rect 20904 21088 20956 21140
rect 22560 21088 22612 21140
rect 23112 21088 23164 21140
rect 10876 21020 10928 21072
rect 11060 21020 11112 21072
rect 11704 21020 11756 21072
rect 13820 21063 13872 21072
rect 13820 21029 13829 21063
rect 13829 21029 13863 21063
rect 13863 21029 13872 21063
rect 13820 21020 13872 21029
rect 22468 21063 22520 21072
rect 22468 21029 22477 21063
rect 22477 21029 22511 21063
rect 22511 21029 22520 21063
rect 22468 21020 22520 21029
rect 23020 21020 23072 21072
rect 23204 21063 23256 21072
rect 23204 21029 23213 21063
rect 23213 21029 23247 21063
rect 23247 21029 23256 21063
rect 23204 21020 23256 21029
rect 24216 21088 24268 21140
rect 24768 21131 24820 21140
rect 24768 21097 24777 21131
rect 24777 21097 24811 21131
rect 24811 21097 24820 21131
rect 24768 21088 24820 21097
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 17776 20995 17828 21004
rect 17776 20961 17810 20995
rect 17810 20961 17828 20995
rect 17776 20952 17828 20961
rect 20904 20995 20956 21004
rect 20904 20961 20913 20995
rect 20913 20961 20947 20995
rect 20947 20961 20956 20995
rect 20904 20952 20956 20961
rect 25044 20952 25096 21004
rect 10140 20884 10192 20936
rect 10416 20927 10468 20936
rect 10416 20893 10425 20927
rect 10425 20893 10459 20927
rect 10459 20893 10468 20927
rect 10416 20884 10468 20893
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 16488 20927 16540 20936
rect 16488 20893 16497 20927
rect 16497 20893 16531 20927
rect 16531 20893 16540 20927
rect 16488 20884 16540 20893
rect 16580 20927 16632 20936
rect 16580 20893 16589 20927
rect 16589 20893 16623 20927
rect 16623 20893 16632 20927
rect 16580 20884 16632 20893
rect 22652 20884 22704 20936
rect 13728 20816 13780 20868
rect 22744 20859 22796 20868
rect 22744 20825 22753 20859
rect 22753 20825 22787 20859
rect 22787 20825 22796 20859
rect 22744 20816 22796 20825
rect 13544 20791 13596 20800
rect 13544 20757 13553 20791
rect 13553 20757 13587 20791
rect 13587 20757 13596 20791
rect 13544 20748 13596 20757
rect 16028 20791 16080 20800
rect 16028 20757 16037 20791
rect 16037 20757 16071 20791
rect 16071 20757 16080 20791
rect 16028 20748 16080 20757
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 20720 20748 20772 20800
rect 23664 20748 23716 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 13636 20544 13688 20596
rect 14096 20544 14148 20596
rect 16580 20544 16632 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 16488 20519 16540 20528
rect 16488 20485 16497 20519
rect 16497 20485 16531 20519
rect 16531 20485 16540 20519
rect 16488 20476 16540 20485
rect 20904 20544 20956 20596
rect 23112 20544 23164 20596
rect 25044 20587 25096 20596
rect 25044 20553 25053 20587
rect 25053 20553 25087 20587
rect 25087 20553 25096 20587
rect 25044 20544 25096 20553
rect 17960 20408 18012 20460
rect 10416 20272 10468 20324
rect 10784 20272 10836 20324
rect 10876 20247 10928 20256
rect 10876 20213 10885 20247
rect 10885 20213 10919 20247
rect 10919 20213 10928 20247
rect 10876 20204 10928 20213
rect 12808 20204 12860 20256
rect 13728 20383 13780 20392
rect 13728 20349 13762 20383
rect 13762 20349 13780 20383
rect 13728 20340 13780 20349
rect 16948 20315 17000 20324
rect 16948 20281 16957 20315
rect 16957 20281 16991 20315
rect 16991 20281 17000 20315
rect 16948 20272 17000 20281
rect 18880 20340 18932 20392
rect 20444 20315 20496 20324
rect 20444 20281 20453 20315
rect 20453 20281 20487 20315
rect 20487 20281 20496 20315
rect 20444 20272 20496 20281
rect 21180 20315 21232 20324
rect 21180 20281 21189 20315
rect 21189 20281 21223 20315
rect 21223 20281 21232 20315
rect 21180 20272 21232 20281
rect 25136 20272 25188 20324
rect 19432 20247 19484 20256
rect 19432 20213 19441 20247
rect 19441 20213 19475 20247
rect 19475 20213 19484 20247
rect 19432 20204 19484 20213
rect 20720 20204 20772 20256
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 24768 20204 24820 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 10876 20000 10928 20052
rect 13360 20000 13412 20052
rect 12900 19932 12952 19984
rect 13820 20000 13872 20052
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 20444 20000 20496 20052
rect 21180 20000 21232 20052
rect 23112 20043 23164 20052
rect 23112 20009 23121 20043
rect 23121 20009 23155 20043
rect 23155 20009 23164 20043
rect 23112 20000 23164 20009
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 14096 19932 14148 19984
rect 15568 19975 15620 19984
rect 15568 19941 15602 19975
rect 15602 19941 15620 19975
rect 15568 19932 15620 19941
rect 18328 19975 18380 19984
rect 18328 19941 18337 19975
rect 18337 19941 18371 19975
rect 18371 19941 18380 19975
rect 18328 19932 18380 19941
rect 22008 19975 22060 19984
rect 22008 19941 22020 19975
rect 22020 19941 22060 19975
rect 22008 19932 22060 19941
rect 23940 19932 23992 19984
rect 10692 19907 10744 19916
rect 10692 19873 10726 19907
rect 10726 19873 10744 19907
rect 10692 19864 10744 19873
rect 12808 19864 12860 19916
rect 14004 19864 14056 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 17776 19864 17828 19916
rect 20536 19864 20588 19916
rect 21824 19864 21876 19916
rect 24032 19864 24084 19916
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 18420 19839 18472 19848
rect 16948 19728 17000 19780
rect 18420 19805 18429 19839
rect 18429 19805 18463 19839
rect 18463 19805 18472 19839
rect 18420 19796 18472 19805
rect 18788 19728 18840 19780
rect 25136 19796 25188 19848
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 16672 19703 16724 19712
rect 16672 19669 16681 19703
rect 16681 19669 16715 19703
rect 16715 19669 16724 19703
rect 16672 19660 16724 19669
rect 24952 19660 25004 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 12900 19499 12952 19508
rect 12900 19465 12909 19499
rect 12909 19465 12943 19499
rect 12943 19465 12952 19499
rect 12900 19456 12952 19465
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 15568 19456 15620 19508
rect 16488 19456 16540 19508
rect 18420 19456 18472 19508
rect 22008 19456 22060 19508
rect 22100 19456 22152 19508
rect 23940 19499 23992 19508
rect 23940 19465 23949 19499
rect 23949 19465 23983 19499
rect 23983 19465 23992 19499
rect 23940 19456 23992 19465
rect 10416 19388 10468 19440
rect 10784 19388 10836 19440
rect 16580 19388 16632 19440
rect 17500 19388 17552 19440
rect 18328 19388 18380 19440
rect 10140 19184 10192 19236
rect 11244 19252 11296 19304
rect 12808 19252 12860 19304
rect 18788 19320 18840 19372
rect 18328 19252 18380 19304
rect 19064 19295 19116 19304
rect 19064 19261 19073 19295
rect 19073 19261 19107 19295
rect 19107 19261 19116 19295
rect 19064 19252 19116 19261
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 11152 19227 11204 19236
rect 11152 19193 11161 19227
rect 11161 19193 11195 19227
rect 11195 19193 11204 19227
rect 11152 19184 11204 19193
rect 13360 19184 13412 19236
rect 17776 19227 17828 19236
rect 17776 19193 17785 19227
rect 17785 19193 17819 19227
rect 17819 19193 17828 19227
rect 17776 19184 17828 19193
rect 18144 19227 18196 19236
rect 18144 19193 18169 19227
rect 18169 19193 18196 19227
rect 18144 19184 18196 19193
rect 18696 19227 18748 19236
rect 18696 19193 18705 19227
rect 18705 19193 18739 19227
rect 18739 19193 18748 19227
rect 18696 19184 18748 19193
rect 21640 19184 21692 19236
rect 21824 19184 21876 19236
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 13820 19116 13872 19168
rect 22100 19159 22152 19168
rect 22100 19125 22109 19159
rect 22109 19125 22143 19159
rect 22143 19125 22152 19159
rect 22100 19116 22152 19125
rect 23664 19116 23716 19168
rect 25320 19252 25372 19304
rect 26240 19252 26292 19304
rect 25136 19184 25188 19236
rect 25504 19159 25556 19168
rect 25504 19125 25513 19159
rect 25513 19125 25547 19159
rect 25547 19125 25556 19159
rect 25504 19116 25556 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 12992 18912 13044 18964
rect 14004 18912 14056 18964
rect 21824 18912 21876 18964
rect 25136 18955 25188 18964
rect 25136 18921 25145 18955
rect 25145 18921 25179 18955
rect 25179 18921 25188 18955
rect 25136 18912 25188 18921
rect 11152 18844 11204 18896
rect 13544 18887 13596 18896
rect 10784 18776 10836 18828
rect 11888 18776 11940 18828
rect 13544 18853 13553 18887
rect 13553 18853 13587 18887
rect 13587 18853 13596 18887
rect 13544 18844 13596 18853
rect 13820 18887 13872 18896
rect 13820 18853 13829 18887
rect 13829 18853 13863 18887
rect 13863 18853 13872 18887
rect 13820 18844 13872 18853
rect 16672 18844 16724 18896
rect 21364 18844 21416 18896
rect 13452 18776 13504 18828
rect 23480 18776 23532 18828
rect 10600 18708 10652 18760
rect 15292 18708 15344 18760
rect 16580 18708 16632 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 21640 18708 21692 18760
rect 23664 18708 23716 18760
rect 20720 18640 20772 18692
rect 10416 18615 10468 18624
rect 10416 18581 10425 18615
rect 10425 18581 10459 18615
rect 10459 18581 10468 18615
rect 10416 18572 10468 18581
rect 10692 18572 10744 18624
rect 13728 18572 13780 18624
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 18696 18572 18748 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10416 18368 10468 18420
rect 10968 18300 11020 18352
rect 13544 18368 13596 18420
rect 14004 18411 14056 18420
rect 14004 18377 14013 18411
rect 14013 18377 14047 18411
rect 14047 18377 14056 18411
rect 14004 18368 14056 18377
rect 15292 18368 15344 18420
rect 13820 18300 13872 18352
rect 15384 18343 15436 18352
rect 15384 18309 15393 18343
rect 15393 18309 15427 18343
rect 15427 18309 15436 18343
rect 15384 18300 15436 18309
rect 16672 18368 16724 18420
rect 21456 18368 21508 18420
rect 23480 18411 23532 18420
rect 23480 18377 23489 18411
rect 23489 18377 23523 18411
rect 23523 18377 23532 18411
rect 23480 18368 23532 18377
rect 16580 18300 16632 18352
rect 23664 18300 23716 18352
rect 24860 18275 24912 18284
rect 24860 18241 24869 18275
rect 24869 18241 24903 18275
rect 24903 18241 24912 18275
rect 24860 18232 24912 18241
rect 25504 18232 25556 18284
rect 10784 18096 10836 18148
rect 11244 18139 11296 18148
rect 11244 18105 11253 18139
rect 11253 18105 11287 18139
rect 11287 18105 11296 18139
rect 11244 18096 11296 18105
rect 16672 18164 16724 18216
rect 24952 18139 25004 18148
rect 24952 18105 24961 18139
rect 24961 18105 24995 18139
rect 24995 18105 25004 18139
rect 24952 18096 25004 18105
rect 10692 18028 10744 18080
rect 11888 18028 11940 18080
rect 13544 18071 13596 18080
rect 13544 18037 13553 18071
rect 13553 18037 13587 18071
rect 13587 18037 13596 18071
rect 13544 18028 13596 18037
rect 15476 18028 15528 18080
rect 16304 18028 16356 18080
rect 16580 18028 16632 18080
rect 17960 18028 18012 18080
rect 18696 18071 18748 18080
rect 18696 18037 18705 18071
rect 18705 18037 18739 18071
rect 18739 18037 18748 18071
rect 18696 18028 18748 18037
rect 21364 18071 21416 18080
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 21640 18071 21692 18080
rect 21640 18037 21649 18071
rect 21649 18037 21683 18071
rect 21683 18037 21692 18071
rect 21640 18028 21692 18037
rect 23388 18028 23440 18080
rect 23572 18028 23624 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 10784 17867 10836 17876
rect 10784 17833 10793 17867
rect 10793 17833 10827 17867
rect 10827 17833 10836 17867
rect 10784 17824 10836 17833
rect 11244 17867 11296 17876
rect 11244 17833 11253 17867
rect 11253 17833 11287 17867
rect 11287 17833 11296 17867
rect 11244 17824 11296 17833
rect 13544 17824 13596 17876
rect 15476 17867 15528 17876
rect 15476 17833 15485 17867
rect 15485 17833 15519 17867
rect 15519 17833 15528 17867
rect 15476 17824 15528 17833
rect 18144 17867 18196 17876
rect 18144 17833 18153 17867
rect 18153 17833 18187 17867
rect 18187 17833 18196 17867
rect 18144 17824 18196 17833
rect 24768 17824 24820 17876
rect 14464 17756 14516 17808
rect 21456 17799 21508 17808
rect 21456 17765 21465 17799
rect 21465 17765 21499 17799
rect 21499 17765 21508 17799
rect 21456 17756 21508 17765
rect 23204 17756 23256 17808
rect 17500 17688 17552 17740
rect 18052 17688 18104 17740
rect 22836 17688 22888 17740
rect 13820 17620 13872 17672
rect 17960 17620 18012 17672
rect 21548 17663 21600 17672
rect 21548 17629 21557 17663
rect 21557 17629 21591 17663
rect 21591 17629 21600 17663
rect 21548 17620 21600 17629
rect 23848 17663 23900 17672
rect 23848 17629 23857 17663
rect 23857 17629 23891 17663
rect 23891 17629 23900 17663
rect 23848 17620 23900 17629
rect 24216 17620 24268 17672
rect 21824 17552 21876 17604
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 16856 17484 16908 17536
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 21916 17484 21968 17536
rect 23480 17484 23532 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 15752 17280 15804 17332
rect 16304 17280 16356 17332
rect 17500 17323 17552 17332
rect 17500 17289 17509 17323
rect 17509 17289 17543 17323
rect 17543 17289 17552 17323
rect 17500 17280 17552 17289
rect 17960 17280 18012 17332
rect 18328 17280 18380 17332
rect 16120 17255 16172 17264
rect 16120 17221 16129 17255
rect 16129 17221 16163 17255
rect 16163 17221 16172 17255
rect 16120 17212 16172 17221
rect 16580 17212 16632 17264
rect 18144 17255 18196 17264
rect 18144 17221 18153 17255
rect 18153 17221 18187 17255
rect 18187 17221 18196 17255
rect 18144 17212 18196 17221
rect 12808 17076 12860 17128
rect 13820 17076 13872 17128
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 18696 17144 18748 17196
rect 20536 17280 20588 17332
rect 21088 17280 21140 17332
rect 21548 17280 21600 17332
rect 22836 17323 22888 17332
rect 22836 17289 22845 17323
rect 22845 17289 22879 17323
rect 22879 17289 22888 17323
rect 22836 17280 22888 17289
rect 24032 17212 24084 17264
rect 21456 17144 21508 17196
rect 24216 17187 24268 17196
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 23204 17119 23256 17128
rect 13360 17008 13412 17060
rect 23204 17085 23213 17119
rect 23213 17085 23247 17119
rect 23247 17085 23256 17119
rect 23204 17076 23256 17085
rect 16948 17051 17000 17060
rect 16948 17017 16957 17051
rect 16957 17017 16991 17051
rect 16991 17017 17000 17051
rect 16948 17008 17000 17017
rect 18236 17008 18288 17060
rect 18696 17051 18748 17060
rect 18696 17017 18705 17051
rect 18705 17017 18739 17051
rect 18739 17017 18748 17051
rect 18696 17008 18748 17017
rect 19708 17008 19760 17060
rect 23848 17008 23900 17060
rect 24400 17051 24452 17060
rect 24400 17017 24409 17051
rect 24409 17017 24443 17051
rect 24443 17017 24452 17051
rect 24400 17008 24452 17017
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 14464 16940 14516 16992
rect 15016 16983 15068 16992
rect 15016 16949 15025 16983
rect 15025 16949 15059 16983
rect 15059 16949 15068 16983
rect 15016 16940 15068 16949
rect 15936 16940 15988 16992
rect 21824 16940 21876 16992
rect 22008 16940 22060 16992
rect 24124 16940 24176 16992
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 11888 16736 11940 16788
rect 13360 16736 13412 16788
rect 13820 16736 13872 16788
rect 18696 16736 18748 16788
rect 24124 16736 24176 16788
rect 24860 16736 24912 16788
rect 13544 16668 13596 16720
rect 14372 16668 14424 16720
rect 15936 16668 15988 16720
rect 18788 16711 18840 16720
rect 18788 16677 18797 16711
rect 18797 16677 18831 16711
rect 18831 16677 18840 16711
rect 18788 16668 18840 16677
rect 21088 16668 21140 16720
rect 23112 16668 23164 16720
rect 24400 16668 24452 16720
rect 10692 16600 10744 16652
rect 11152 16643 11204 16652
rect 11152 16609 11186 16643
rect 11186 16609 11204 16643
rect 18604 16643 18656 16652
rect 11152 16600 11204 16609
rect 18604 16609 18613 16643
rect 18613 16609 18647 16643
rect 18647 16609 18656 16643
rect 18604 16600 18656 16609
rect 23388 16600 23440 16652
rect 24676 16600 24728 16652
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 16948 16532 17000 16584
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 13452 16439 13504 16448
rect 13452 16405 13461 16439
rect 13461 16405 13495 16439
rect 13495 16405 13504 16439
rect 13452 16396 13504 16405
rect 16764 16396 16816 16448
rect 18420 16396 18472 16448
rect 19156 16396 19208 16448
rect 20536 16396 20588 16448
rect 20996 16396 21048 16448
rect 22376 16439 22428 16448
rect 22376 16405 22385 16439
rect 22385 16405 22419 16439
rect 22419 16405 22428 16439
rect 22376 16396 22428 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 11152 16192 11204 16244
rect 13728 16192 13780 16244
rect 16948 16192 17000 16244
rect 18788 16192 18840 16244
rect 18880 16192 18932 16244
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 23572 16192 23624 16244
rect 10692 16124 10744 16176
rect 21824 16124 21876 16176
rect 23848 16124 23900 16176
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 24768 16192 24820 16244
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 25872 16235 25924 16244
rect 25872 16201 25881 16235
rect 25881 16201 25915 16235
rect 25915 16201 25924 16235
rect 25872 16192 25924 16201
rect 24676 16167 24728 16176
rect 24676 16133 24685 16167
rect 24685 16133 24719 16167
rect 24719 16133 24728 16167
rect 24676 16124 24728 16133
rect 14372 15920 14424 15972
rect 24032 16031 24084 16040
rect 21916 15920 21968 15972
rect 24032 15997 24041 16031
rect 24041 15997 24075 16031
rect 24075 15997 24084 16031
rect 24032 15988 24084 15997
rect 25872 15988 25924 16040
rect 22376 15920 22428 15972
rect 22836 15920 22888 15972
rect 23480 15920 23532 15972
rect 24216 15963 24268 15972
rect 24216 15929 24225 15963
rect 24225 15929 24259 15963
rect 24259 15929 24268 15963
rect 24216 15920 24268 15929
rect 15752 15852 15804 15904
rect 16304 15852 16356 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 13544 15648 13596 15700
rect 14372 15648 14424 15700
rect 16580 15648 16632 15700
rect 21088 15691 21140 15700
rect 21088 15657 21097 15691
rect 21097 15657 21131 15691
rect 21131 15657 21140 15691
rect 21088 15648 21140 15657
rect 21916 15691 21968 15700
rect 21916 15657 21925 15691
rect 21925 15657 21959 15691
rect 21959 15657 21968 15691
rect 21916 15648 21968 15657
rect 23112 15648 23164 15700
rect 24216 15648 24268 15700
rect 25228 15691 25280 15700
rect 25228 15657 25237 15691
rect 25237 15657 25271 15691
rect 25271 15657 25280 15691
rect 25228 15648 25280 15657
rect 16488 15580 16540 15632
rect 17132 15580 17184 15632
rect 17224 15580 17276 15632
rect 22008 15580 22060 15632
rect 17776 15555 17828 15564
rect 17776 15521 17785 15555
rect 17785 15521 17819 15555
rect 17819 15521 17828 15555
rect 17776 15512 17828 15521
rect 22836 15555 22888 15564
rect 22836 15521 22870 15555
rect 22870 15521 22888 15555
rect 22836 15512 22888 15521
rect 25044 15555 25096 15564
rect 25044 15521 25053 15555
rect 25053 15521 25087 15555
rect 25087 15521 25096 15555
rect 25044 15512 25096 15521
rect 16396 15444 16448 15496
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 20996 15444 21048 15496
rect 22560 15487 22612 15496
rect 22560 15453 22569 15487
rect 22569 15453 22603 15487
rect 22603 15453 22612 15487
rect 22560 15444 22612 15453
rect 16120 15308 16172 15360
rect 20168 15351 20220 15360
rect 20168 15317 20177 15351
rect 20177 15317 20211 15351
rect 20211 15317 20220 15351
rect 20168 15308 20220 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 16488 15104 16540 15156
rect 16580 15104 16632 15156
rect 17776 15104 17828 15156
rect 19156 15104 19208 15156
rect 13176 15011 13228 15020
rect 13176 14977 13185 15011
rect 13185 14977 13219 15011
rect 13219 14977 13228 15011
rect 13176 14968 13228 14977
rect 15844 15011 15896 15020
rect 15844 14977 15853 15011
rect 15853 14977 15887 15011
rect 15887 14977 15896 15011
rect 15844 14968 15896 14977
rect 19064 15011 19116 15020
rect 19064 14977 19073 15011
rect 19073 14977 19107 15011
rect 19107 14977 19116 15011
rect 19064 14968 19116 14977
rect 21640 15104 21692 15156
rect 22560 15147 22612 15156
rect 22560 15113 22569 15147
rect 22569 15113 22603 15147
rect 22603 15113 22612 15147
rect 22560 15104 22612 15113
rect 22836 15104 22888 15156
rect 25044 15147 25096 15156
rect 25044 15113 25053 15147
rect 25053 15113 25087 15147
rect 25087 15113 25096 15147
rect 25044 15104 25096 15113
rect 13728 14900 13780 14952
rect 20168 14832 20220 14884
rect 20904 14832 20956 14884
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 19064 14807 19116 14816
rect 19064 14773 19073 14807
rect 19073 14773 19107 14807
rect 19107 14773 19116 14807
rect 19064 14764 19116 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 16396 14560 16448 14612
rect 21364 14560 21416 14612
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 13636 14492 13688 14544
rect 14832 14424 14884 14476
rect 16580 14424 16632 14476
rect 16856 14492 16908 14544
rect 16948 14535 17000 14544
rect 16948 14501 16957 14535
rect 16957 14501 16991 14535
rect 16991 14501 17000 14535
rect 16948 14492 17000 14501
rect 19156 14492 19208 14544
rect 21272 14535 21324 14544
rect 21272 14501 21281 14535
rect 21281 14501 21315 14535
rect 21315 14501 21324 14535
rect 21272 14492 21324 14501
rect 18328 14467 18380 14476
rect 18328 14433 18337 14467
rect 18337 14433 18371 14467
rect 18371 14433 18380 14467
rect 18328 14424 18380 14433
rect 18604 14467 18656 14476
rect 18604 14433 18638 14467
rect 18638 14433 18656 14467
rect 18604 14424 18656 14433
rect 24584 14467 24636 14476
rect 24584 14433 24593 14467
rect 24593 14433 24627 14467
rect 24627 14433 24636 14467
rect 24584 14424 24636 14433
rect 14280 14399 14332 14408
rect 14280 14365 14289 14399
rect 14289 14365 14323 14399
rect 14323 14365 14332 14399
rect 14280 14356 14332 14365
rect 17316 14356 17368 14408
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 13728 14331 13780 14340
rect 13728 14297 13737 14331
rect 13737 14297 13771 14331
rect 13771 14297 13780 14331
rect 13728 14288 13780 14297
rect 15476 14288 15528 14340
rect 20996 14331 21048 14340
rect 20996 14297 21005 14331
rect 21005 14297 21039 14331
rect 21039 14297 21048 14331
rect 20996 14288 21048 14297
rect 19800 14220 19852 14272
rect 21548 14220 21600 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 13820 14016 13872 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 15292 13948 15344 14000
rect 16304 14016 16356 14068
rect 16856 14016 16908 14068
rect 16948 14016 17000 14068
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 20904 14059 20956 14068
rect 17316 13991 17368 14000
rect 17316 13957 17325 13991
rect 17325 13957 17359 13991
rect 17359 13957 17368 13991
rect 17316 13948 17368 13957
rect 18236 13948 18288 14000
rect 18604 13948 18656 14000
rect 20904 14025 20913 14059
rect 20913 14025 20947 14059
rect 20947 14025 20956 14059
rect 20904 14016 20956 14025
rect 21272 14016 21324 14068
rect 21548 14016 21600 14068
rect 24676 14059 24728 14068
rect 24676 14025 24685 14059
rect 24685 14025 24719 14059
rect 24719 14025 24728 14059
rect 24676 14016 24728 14025
rect 16948 13812 17000 13864
rect 19616 13812 19668 13864
rect 19800 13855 19852 13864
rect 19800 13821 19834 13855
rect 19834 13821 19852 13855
rect 19800 13812 19852 13821
rect 13176 13787 13228 13796
rect 13176 13753 13210 13787
rect 13210 13753 13228 13787
rect 13176 13744 13228 13753
rect 15292 13744 15344 13796
rect 16488 13744 16540 13796
rect 16764 13719 16816 13728
rect 16764 13685 16773 13719
rect 16773 13685 16807 13719
rect 16807 13685 16816 13719
rect 16764 13676 16816 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 13728 13472 13780 13524
rect 15292 13472 15344 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 21180 13515 21232 13524
rect 21180 13481 21189 13515
rect 21189 13481 21223 13515
rect 21223 13481 21232 13515
rect 21180 13472 21232 13481
rect 21364 13472 21416 13524
rect 14004 13404 14056 13456
rect 16764 13404 16816 13456
rect 13176 13336 13228 13388
rect 24584 13379 24636 13388
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 24584 13345 24593 13379
rect 24593 13345 24627 13379
rect 24627 13345 24636 13379
rect 24584 13336 24636 13345
rect 14464 13268 14516 13320
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 13636 13200 13688 13252
rect 24768 13243 24820 13252
rect 24768 13209 24777 13243
rect 24777 13209 24811 13243
rect 24811 13209 24820 13243
rect 24768 13200 24820 13209
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 16488 12971 16540 12980
rect 16488 12937 16497 12971
rect 16497 12937 16531 12971
rect 16531 12937 16540 12971
rect 16488 12928 16540 12937
rect 16856 12928 16908 12980
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 12808 12792 12860 12844
rect 16672 12792 16724 12844
rect 16764 12792 16816 12844
rect 13360 12699 13412 12708
rect 13360 12665 13394 12699
rect 13394 12665 13412 12699
rect 13360 12656 13412 12665
rect 16672 12656 16724 12708
rect 16856 12656 16908 12708
rect 16948 12699 17000 12708
rect 16948 12665 16957 12699
rect 16957 12665 16991 12699
rect 16991 12665 17000 12699
rect 16948 12656 17000 12665
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 16580 12588 16632 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 12808 12384 12860 12436
rect 14188 12384 14240 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 16764 12384 16816 12436
rect 25320 12384 25372 12436
rect 14004 12359 14056 12368
rect 14004 12325 14013 12359
rect 14013 12325 14047 12359
rect 14047 12325 14056 12359
rect 14004 12316 14056 12325
rect 16488 12316 16540 12368
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 13268 11883 13320 11892
rect 13268 11849 13277 11883
rect 13277 11849 13311 11883
rect 13311 11849 13320 11883
rect 13268 11840 13320 11849
rect 24676 11883 24728 11892
rect 24676 11849 24685 11883
rect 24685 11849 24719 11883
rect 24719 11849 24728 11883
rect 24676 11840 24728 11849
rect 13268 11636 13320 11688
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 12256 11067 12308 11076
rect 12256 11033 12265 11067
rect 12265 11033 12299 11067
rect 12299 11033 12308 11067
rect 12256 11024 12308 11033
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 11612 10752 11664 10804
rect 12072 10752 12124 10804
rect 11612 10548 11664 10600
rect 11428 10455 11480 10464
rect 11428 10421 11437 10455
rect 11437 10421 11471 10455
rect 11471 10421 11480 10455
rect 11428 10412 11480 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 9864 10072 9916 10124
rect 10968 10072 11020 10124
rect 10876 9979 10928 9988
rect 10876 9945 10885 9979
rect 10885 9945 10919 9979
rect 10919 9945 10928 9979
rect 10876 9936 10928 9945
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 10968 9707 11020 9716
rect 10968 9673 10977 9707
rect 10977 9673 11011 9707
rect 11011 9673 11020 9707
rect 10968 9664 11020 9673
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 9772 9460 9824 9512
rect 24584 9503 24636 9512
rect 24584 9469 24593 9503
rect 24593 9469 24627 9503
rect 24627 9469 24636 9503
rect 24584 9460 24636 9469
rect 24768 9367 24820 9376
rect 24768 9333 24777 9367
rect 24777 9333 24811 9367
rect 24811 9333 24820 9367
rect 24768 9324 24820 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 24584 9095 24636 9104
rect 24584 9061 24593 9095
rect 24593 9061 24627 9095
rect 24627 9061 24636 9095
rect 24584 9052 24636 9061
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 23664 8984 23716 9036
rect 24952 8984 25004 9036
rect 9864 8891 9916 8900
rect 9864 8857 9873 8891
rect 9873 8857 9907 8891
rect 9907 8857 9916 8891
rect 9864 8848 9916 8857
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 25320 8551 25372 8560
rect 25320 8517 25329 8551
rect 25329 8517 25363 8551
rect 25363 8517 25372 8551
rect 25320 8508 25372 8517
rect 23848 8415 23900 8424
rect 23848 8381 23857 8415
rect 23857 8381 23891 8415
rect 23891 8381 23900 8415
rect 23848 8372 23900 8381
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 19340 7939 19392 7948
rect 19340 7905 19349 7939
rect 19349 7905 19383 7939
rect 19383 7905 19392 7939
rect 19340 7896 19392 7905
rect 21824 7896 21876 7948
rect 22928 7939 22980 7948
rect 22928 7905 22937 7939
rect 22937 7905 22971 7939
rect 22971 7905 22980 7939
rect 22928 7896 22980 7905
rect 24216 7896 24268 7948
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 24768 7692 24820 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 19340 7531 19392 7540
rect 19340 7497 19349 7531
rect 19349 7497 19383 7531
rect 19383 7497 19392 7531
rect 19340 7488 19392 7497
rect 22928 7531 22980 7540
rect 22928 7497 22937 7531
rect 22937 7497 22971 7531
rect 22971 7497 22980 7531
rect 22928 7488 22980 7497
rect 24216 7488 24268 7540
rect 24584 7327 24636 7336
rect 24584 7293 24593 7327
rect 24593 7293 24627 7327
rect 24627 7293 24636 7327
rect 24584 7284 24636 7293
rect 24676 7148 24728 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 23480 6808 23532 6860
rect 24768 6808 24820 6860
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 24768 6443 24820 6452
rect 24768 6409 24777 6443
rect 24777 6409 24811 6443
rect 24811 6409 24820 6443
rect 24768 6400 24820 6409
rect 14556 6196 14608 6248
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 15200 6171 15252 6180
rect 15200 6137 15209 6171
rect 15209 6137 15243 6171
rect 15243 6137 15252 6171
rect 15200 6128 15252 6137
rect 26148 6060 26200 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 23664 5763 23716 5772
rect 23664 5729 23673 5763
rect 23673 5729 23707 5763
rect 23707 5729 23716 5763
rect 23664 5720 23716 5729
rect 24952 5763 25004 5772
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 23848 5652 23900 5661
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 23664 5312 23716 5364
rect 24952 5312 25004 5364
rect 23664 5151 23716 5160
rect 23664 5117 23673 5151
rect 23673 5117 23707 5151
rect 23707 5117 23716 5151
rect 23664 5108 23716 5117
rect 25136 5015 25188 5024
rect 25136 4981 25145 5015
rect 25145 4981 25179 5015
rect 25179 4981 25188 5015
rect 25136 4972 25188 4981
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 23848 4632 23900 4684
rect 24216 4632 24268 4684
rect 24676 4428 24728 4480
rect 24768 4471 24820 4480
rect 24768 4437 24777 4471
rect 24777 4437 24811 4471
rect 24811 4437 24820 4471
rect 24768 4428 24820 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 23848 4267 23900 4276
rect 23848 4233 23857 4267
rect 23857 4233 23891 4267
rect 23891 4233 23900 4267
rect 23848 4224 23900 4233
rect 23940 4020 23992 4072
rect 24216 3952 24268 4004
rect 24400 3927 24452 3936
rect 24400 3893 24409 3927
rect 24409 3893 24443 3927
rect 24443 3893 24452 3927
rect 24400 3884 24452 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 24400 3612 24452 3664
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 24860 3544 24912 3596
rect 24768 3340 24820 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 23756 3136 23808 3188
rect 24860 3179 24912 3188
rect 24860 3145 24869 3179
rect 24869 3145 24903 3179
rect 24903 3145 24912 3179
rect 24860 3136 24912 3145
rect 23480 3111 23532 3120
rect 23480 3077 23489 3111
rect 23489 3077 23523 3111
rect 23523 3077 23532 3111
rect 23480 3068 23532 3077
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 23664 2975 23716 2984
rect 23664 2941 23673 2975
rect 23673 2941 23707 2975
rect 23707 2941 23716 2975
rect 23664 2932 23716 2941
rect 24952 2975 25004 2984
rect 24952 2941 24961 2975
rect 24961 2941 24995 2975
rect 24995 2941 25004 2975
rect 24952 2932 25004 2941
rect 22560 2907 22612 2916
rect 22560 2873 22569 2907
rect 22569 2873 22603 2907
rect 22603 2873 22612 2907
rect 22560 2864 22612 2873
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 25320 2499 25372 2508
rect 25320 2465 25329 2499
rect 25329 2465 25363 2499
rect 25363 2465 25372 2499
rect 25320 2456 25372 2465
rect 23020 2295 23072 2304
rect 23020 2261 23029 2295
rect 23029 2261 23063 2295
rect 23063 2261 23072 2295
rect 23020 2252 23072 2261
rect 25504 2295 25556 2304
rect 25504 2261 25513 2295
rect 25513 2261 25547 2295
rect 25547 2261 25556 2295
rect 25504 2252 25556 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 938 27520 994 28000
rect 1582 27520 1638 28000
rect 2226 27520 2282 28000
rect 2870 27520 2926 28000
rect 3606 27520 3662 28000
rect 4250 27520 4306 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6274 27520 6330 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8206 27520 8262 28000
rect 8942 27520 8998 28000
rect 9586 27520 9642 28000
rect 10230 27520 10286 28000
rect 10874 27520 10930 28000
rect 11610 27520 11666 28000
rect 12254 27520 12310 28000
rect 12898 27520 12954 28000
rect 13542 27520 13598 28000
rect 14278 27520 14334 28000
rect 14922 27520 14978 28000
rect 15566 27520 15622 28000
rect 16210 27520 16266 28000
rect 16854 27520 16910 28000
rect 17590 27520 17646 28000
rect 18234 27520 18290 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20258 27520 20314 28000
rect 20902 27520 20958 28000
rect 21546 27520 21602 28000
rect 22190 27520 22246 28000
rect 22926 27520 22982 28000
rect 23570 27520 23626 28000
rect 24214 27520 24270 28000
rect 24766 27704 24822 27713
rect 24766 27639 24822 27648
rect 308 27418 336 27520
rect 308 27390 428 27418
rect 400 12753 428 27390
rect 952 23633 980 27520
rect 938 23624 994 23633
rect 938 23559 994 23568
rect 1596 22545 1624 27520
rect 1582 22536 1638 22545
rect 1582 22471 1638 22480
rect 2240 19825 2268 27520
rect 2226 19816 2282 19825
rect 2226 19751 2282 19760
rect 2884 17241 2912 27520
rect 3620 18873 3648 27520
rect 4264 23769 4292 27520
rect 4908 24177 4936 27520
rect 5552 24721 5580 27520
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5538 24712 5594 24721
rect 5538 24647 5594 24656
rect 4894 24168 4950 24177
rect 4894 24103 4950 24112
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 4250 23760 4306 23769
rect 4250 23695 4306 23704
rect 6288 23089 6316 27520
rect 6274 23080 6330 23089
rect 6274 23015 6330 23024
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6932 19281 6960 27520
rect 6918 19272 6974 19281
rect 6918 19207 6974 19216
rect 3606 18864 3662 18873
rect 3606 18799 3662 18808
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 7576 17785 7604 27520
rect 7562 17776 7618 17785
rect 7562 17711 7618 17720
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 2870 17232 2926 17241
rect 2870 17167 2926 17176
rect 8220 17105 8248 27520
rect 8956 19417 8984 27520
rect 8942 19408 8998 19417
rect 8942 19343 8998 19352
rect 8206 17096 8262 17105
rect 8206 17031 8262 17040
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 3330 16008 3386 16017
rect 3330 15943 3386 15952
rect 3344 14113 3372 15943
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 3330 14104 3386 14113
rect 5622 14096 5918 14116
rect 3330 14039 3386 14048
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 386 12744 442 12753
rect 386 12679 442 12688
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 9600 9602 9628 27520
rect 10244 25786 10272 27520
rect 10152 25758 10272 25786
rect 10152 24818 10180 25758
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 10140 24812 10192 24818
rect 10140 24754 10192 24760
rect 9692 9738 9720 24754
rect 10888 24698 10916 27520
rect 9784 24670 10916 24698
rect 9784 20074 9812 24670
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 10336 23866 10364 24210
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 9864 23792 9916 23798
rect 9864 23734 9916 23740
rect 9954 23760 10010 23769
rect 9876 20210 9904 23734
rect 9954 23695 10010 23704
rect 9968 22234 9996 23695
rect 10796 23526 10824 24006
rect 10784 23520 10836 23526
rect 11072 23474 11100 24142
rect 11256 23866 11284 24210
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 10784 23462 10836 23468
rect 10980 23446 11100 23474
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10980 23322 11008 23446
rect 11256 23322 11284 23802
rect 11440 23730 11468 24006
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 11428 23520 11480 23526
rect 11428 23462 11480 23468
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11440 23254 11468 23462
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 10152 22438 10180 23054
rect 10980 22778 11008 23122
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10692 22432 10744 22438
rect 10692 22374 10744 22380
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9968 21554 9996 22170
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9876 20182 9996 20210
rect 9784 20046 9904 20074
rect 9876 10130 9904 20046
rect 9864 10124 9916 10130
rect 9864 10066 9916 10072
rect 9692 9710 9812 9738
rect 9600 9574 9720 9602
rect 9692 9042 9720 9574
rect 9784 9518 9812 9710
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 9692 8634 9720 8978
rect 9862 8936 9918 8945
rect 9862 8871 9864 8880
rect 9916 8871 9918 8880
rect 9864 8842 9916 8848
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 9968 6361 9996 20182
rect 9954 6352 10010 6361
rect 9954 6287 10010 6296
rect 10060 5817 10088 21558
rect 10152 20942 10180 22374
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 21486 10732 22374
rect 10876 22024 10928 22030
rect 10874 21992 10876 22001
rect 10928 21992 10930 22001
rect 10796 21950 10874 21978
rect 10796 21690 10824 21950
rect 10874 21927 10930 21936
rect 10876 21888 10928 21894
rect 10876 21830 10928 21836
rect 10784 21684 10836 21690
rect 10784 21626 10836 21632
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10888 21418 10916 21830
rect 10980 21554 11008 22714
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10980 21146 11008 21490
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 11072 21078 11100 21966
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 11060 21072 11112 21078
rect 11060 21014 11112 21020
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10416 20936 10468 20942
rect 10416 20878 10468 20884
rect 10428 20330 10456 20878
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10784 20324 10836 20330
rect 10784 20266 10836 20272
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19446 10456 19790
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10140 19236 10192 19242
rect 10140 19178 10192 19184
rect 10152 18873 10180 19178
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10138 18864 10194 18873
rect 10138 18799 10194 18808
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 18426 10456 18566
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10612 18068 10640 18702
rect 10704 18630 10732 19858
rect 10796 19446 10824 20266
rect 10888 20262 10916 21014
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10888 20058 10916 20198
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10796 18834 10824 19382
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18902 11192 19178
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10968 18352 11020 18358
rect 10968 18294 11020 18300
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10692 18080 10744 18086
rect 10612 18040 10692 18068
rect 10692 18022 10744 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16697 10732 18022
rect 10796 17882 10824 18090
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10690 16688 10746 16697
rect 10690 16623 10692 16632
rect 10744 16623 10746 16632
rect 10692 16594 10744 16600
rect 10704 16182 10732 16594
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10704 16017 10732 16118
rect 10690 16008 10746 16017
rect 10690 15943 10746 15952
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10980 10282 11008 18294
rect 11256 18154 11284 19246
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11256 17882 11284 18090
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11164 16561 11192 16594
rect 11150 16552 11206 16561
rect 11150 16487 11206 16496
rect 11164 16250 11192 16487
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11624 10810 11652 27520
rect 12268 27418 12296 27520
rect 12084 27390 12296 27418
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11716 21078 11744 21286
rect 11704 21072 11756 21078
rect 11704 21014 11756 21020
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18834 11928 19110
rect 11888 18828 11940 18834
rect 11888 18770 11940 18776
rect 11900 18086 11928 18770
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 16794 11928 18022
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 12084 11218 12112 27390
rect 12162 24168 12218 24177
rect 12912 24154 12940 27520
rect 12912 24126 13308 24154
rect 12162 24103 12218 24112
rect 12176 23662 12204 24103
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 13176 24064 13228 24070
rect 13176 24006 13228 24012
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 23118 12480 23462
rect 12544 23254 12572 24006
rect 12990 23760 13046 23769
rect 12990 23695 12992 23704
rect 13044 23695 13046 23704
rect 12992 23666 13044 23672
rect 12532 23248 12584 23254
rect 12532 23190 12584 23196
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12452 22778 12480 23054
rect 13004 22982 13032 23666
rect 13084 23248 13136 23254
rect 13084 23190 13136 23196
rect 12992 22976 13044 22982
rect 12992 22918 13044 22924
rect 13096 22778 13124 23190
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12820 19922 12848 20198
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12820 19310 12848 19858
rect 12912 19825 12940 19926
rect 12898 19816 12954 19825
rect 12898 19751 12954 19760
rect 12912 19514 12940 19751
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12808 19304 12860 19310
rect 12808 19246 12860 19252
rect 12820 17134 12848 19246
rect 13004 18970 13032 19654
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12820 16998 12848 17070
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16697 12848 16934
rect 12806 16688 12862 16697
rect 12806 16623 12862 16632
rect 12820 14074 12848 16623
rect 13188 15026 13216 24006
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12820 12850 12848 14010
rect 13176 13796 13228 13802
rect 13176 13738 13228 13744
rect 13188 13394 13216 13738
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12442 12848 12786
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 13280 11898 13308 24126
rect 13556 22681 13584 27520
rect 14002 24712 14058 24721
rect 14002 24647 14004 24656
rect 14056 24647 14058 24656
rect 14004 24618 14056 24624
rect 14292 24410 14320 27520
rect 14936 25242 14964 27520
rect 14752 25214 14964 25242
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14280 24404 14332 24410
rect 14280 24346 14332 24352
rect 14384 24070 14412 24686
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 13820 23520 13872 23526
rect 13740 23468 13820 23474
rect 14188 23520 14240 23526
rect 13740 23462 13872 23468
rect 14094 23488 14150 23497
rect 13740 23446 13860 23462
rect 13740 23186 13768 23446
rect 14188 23462 14240 23468
rect 14094 23423 14150 23432
rect 13728 23180 13780 23186
rect 13728 23122 13780 23128
rect 13634 23080 13690 23089
rect 13634 23015 13690 23024
rect 13542 22672 13598 22681
rect 13542 22607 13598 22616
rect 13648 22098 13676 23015
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13636 22092 13688 22098
rect 13636 22034 13688 22040
rect 13648 21690 13676 22034
rect 13740 21978 13768 22918
rect 14108 22030 14136 23423
rect 14096 22024 14148 22030
rect 13740 21950 13952 21978
rect 14096 21966 14148 21972
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13636 21140 13688 21146
rect 13636 21082 13688 21088
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13372 19242 13400 19994
rect 13450 19952 13506 19961
rect 13450 19887 13506 19896
rect 13464 19854 13492 19887
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13360 19236 13412 19242
rect 13360 19178 13412 19184
rect 13464 18834 13492 19790
rect 13556 18902 13584 20742
rect 13648 20602 13676 21082
rect 13740 21049 13768 21830
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 13832 21078 13860 21490
rect 13924 21146 13952 21950
rect 14108 21554 14136 21966
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13820 21072 13872 21078
rect 13726 21040 13782 21049
rect 13820 21014 13872 21020
rect 13726 20975 13782 20984
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13740 20398 13768 20810
rect 13728 20392 13780 20398
rect 13726 20360 13728 20369
rect 13780 20360 13782 20369
rect 13726 20295 13782 20304
rect 13832 20058 13860 21014
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 14016 19922 14044 21286
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20602 14136 20878
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14108 19990 14136 20538
rect 14096 19984 14148 19990
rect 14096 19926 14148 19932
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13832 18902 13860 19110
rect 14200 18986 14228 23462
rect 14292 23322 14320 23598
rect 14384 23361 14412 24006
rect 14370 23352 14426 23361
rect 14280 23316 14332 23322
rect 14370 23287 14426 23296
rect 14280 23258 14332 23264
rect 14476 22506 14504 24618
rect 14752 23526 14780 25214
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24818 14872 25094
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14844 24410 14872 24754
rect 15580 24410 15608 27520
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 14844 23662 14872 24346
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 15856 23526 15884 24210
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 15292 23520 15344 23526
rect 15292 23462 15344 23468
rect 15844 23520 15896 23526
rect 15844 23462 15896 23468
rect 14740 23112 14792 23118
rect 14740 23054 14792 23060
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14476 22234 14504 22442
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14292 21622 14320 21966
rect 14280 21616 14332 21622
rect 14280 21558 14332 21564
rect 14004 18964 14056 18970
rect 14200 18958 14320 18986
rect 14004 18906 14056 18912
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13556 18426 13584 18838
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13556 17882 13584 18022
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13360 17060 13412 17066
rect 13360 17002 13412 17008
rect 13372 16794 13400 17002
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13556 16726 13584 17478
rect 13740 16810 13768 18566
rect 13832 18358 13860 18838
rect 14016 18426 14044 18906
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13832 17678 13860 18294
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17134 13860 17614
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13740 16794 13860 16810
rect 13740 16788 13872 16794
rect 13740 16782 13820 16788
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13280 11694 13308 11834
rect 13268 11688 13320 11694
rect 12898 11656 12954 11665
rect 13268 11630 13320 11636
rect 12898 11591 12954 11600
rect 12912 11558 12940 11591
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 10810 12112 11154
rect 12254 11112 12310 11121
rect 12254 11047 12256 11056
rect 12308 11047 12310 11056
rect 12256 11018 12308 11024
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11624 10606 11652 10746
rect 11612 10600 11664 10606
rect 11426 10568 11482 10577
rect 11612 10542 11664 10548
rect 11426 10503 11482 10512
rect 11440 10470 11468 10503
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 10796 10254 11008 10282
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10244 9489 10272 9590
rect 10230 9480 10286 9489
rect 10230 9415 10286 9424
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10046 5808 10102 5817
rect 10046 5743 10102 5752
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 10796 5137 10824 10254
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10874 10024 10930 10033
rect 10874 9959 10876 9968
rect 10928 9959 10930 9968
rect 10876 9930 10928 9936
rect 10980 9722 11008 10066
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 13372 8265 13400 12650
rect 13358 8256 13414 8265
rect 13358 8191 13414 8200
rect 10782 5128 10838 5137
rect 10782 5063 10838 5072
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 13464 2961 13492 16390
rect 13556 15706 13584 16662
rect 13740 16250 13768 16782
rect 13820 16730 13872 16736
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 14292 14906 14320 18958
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 14476 16998 14504 17750
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14384 16726 14412 16934
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14384 15978 14412 16662
rect 14372 15972 14424 15978
rect 14372 15914 14424 15920
rect 14384 15706 14412 15914
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13648 13258 13676 14486
rect 13740 14346 13768 14894
rect 14292 14878 14412 14906
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 14292 14074 14320 14350
rect 13820 14068 13872 14074
rect 13740 14028 13820 14056
rect 13740 13530 13768 14028
rect 13820 14010 13872 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 14004 13456 14056 13462
rect 14004 13398 14056 13404
rect 14186 13424 14242 13433
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 14016 12753 14044 13398
rect 14186 13359 14242 13368
rect 14200 13326 14228 13359
rect 14188 13320 14240 13326
rect 14384 13297 14412 14878
rect 14464 13320 14516 13326
rect 14188 13262 14240 13268
rect 14370 13288 14426 13297
rect 14002 12744 14058 12753
rect 14002 12679 14058 12688
rect 14016 12374 14044 12679
rect 14200 12442 14228 13262
rect 14464 13262 14516 13268
rect 14370 13223 14426 13232
rect 14476 12646 14504 13262
rect 14464 12640 14516 12646
rect 14464 12582 14516 12588
rect 14476 12442 14504 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 13450 2952 13506 2961
rect 13450 2887 13506 2896
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 14016 480 14044 8191
rect 14568 6254 14596 22646
rect 14752 22642 14780 23054
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22658 15332 23462
rect 15120 22642 15332 22658
rect 14740 22636 14792 22642
rect 14740 22578 14792 22584
rect 15108 22636 15332 22642
rect 15160 22630 15332 22636
rect 15108 22578 15160 22584
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14660 21486 14688 22510
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14660 21146 14688 21422
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 15474 21040 15530 21049
rect 15474 20975 15530 20984
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15304 19514 15332 19858
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15304 18426 15332 18702
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15028 16833 15056 16934
rect 15014 16824 15070 16833
rect 15014 16759 15070 16768
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14844 14074 14872 14418
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15304 13802 15332 13942
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 15304 13530 15332 13738
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15396 6497 15424 18294
rect 15488 18086 15516 20975
rect 15580 19990 15608 21626
rect 15568 19984 15620 19990
rect 15568 19926 15620 19932
rect 15580 19514 15608 19926
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15488 17882 15516 18022
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15764 16590 15792 17274
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15764 15910 15792 16526
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15856 15026 15884 23462
rect 16118 22536 16174 22545
rect 16118 22471 16120 22480
rect 16172 22471 16174 22480
rect 16120 22442 16172 22448
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16726 15976 16934
rect 15936 16720 15988 16726
rect 15936 16662 15988 16668
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15488 14346 15516 14758
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15382 6488 15438 6497
rect 15382 6423 15438 6432
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 15198 6216 15254 6225
rect 15198 6151 15200 6160
rect 15252 6151 15254 6160
rect 15200 6122 15252 6128
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 16040 2417 16068 20742
rect 16120 17264 16172 17270
rect 16118 17232 16120 17241
rect 16172 17232 16174 17241
rect 16118 17167 16174 17176
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 3097 16160 15302
rect 16224 15065 16252 27520
rect 16868 23866 16896 27520
rect 17604 27418 17632 27520
rect 17604 27390 17908 27418
rect 16856 23860 16908 23866
rect 16856 23802 16908 23808
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17038 23352 17094 23361
rect 17038 23287 17094 23296
rect 16948 23180 17000 23186
rect 16948 23122 17000 23128
rect 16960 22778 16988 23122
rect 16948 22772 17000 22778
rect 16948 22714 17000 22720
rect 16580 22704 16632 22710
rect 16580 22646 16632 22652
rect 16592 21690 16620 22646
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16868 22166 16896 22510
rect 16856 22160 16908 22166
rect 16856 22102 16908 22108
rect 16762 21992 16818 22001
rect 16762 21927 16818 21936
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16776 21622 16804 21927
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 16486 21176 16542 21185
rect 16486 21111 16488 21120
rect 16540 21111 16542 21120
rect 16488 21082 16540 21088
rect 16488 20936 16540 20942
rect 16488 20878 16540 20884
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16500 20534 16528 20878
rect 16592 20602 16620 20878
rect 16580 20596 16632 20602
rect 16580 20538 16632 20544
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16500 19514 16528 20470
rect 16592 20369 16620 20538
rect 16578 20360 16634 20369
rect 16578 20295 16634 20304
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 16592 18766 16620 19382
rect 16684 18902 16712 19654
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16592 18358 16620 18702
rect 16684 18426 16712 18838
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16592 18086 16620 18294
rect 16684 18222 16712 18362
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16304 18080 16356 18086
rect 16304 18022 16356 18028
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16316 17338 16344 18022
rect 16868 17542 16896 22102
rect 17052 22098 17080 23287
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 17052 21622 17080 22034
rect 17040 21616 17092 21622
rect 17040 21558 17092 21564
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 20330 16988 20742
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16960 19786 16988 20266
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16210 15056 16266 15065
rect 16210 14991 16266 15000
rect 16316 14074 16344 15846
rect 16592 15706 16620 17206
rect 16868 17202 16896 17478
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16960 16590 16988 17002
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 17130 16552 17186 16561
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 14618 16436 15438
rect 16500 15162 16528 15574
rect 16592 15162 16620 15642
rect 16776 15502 16804 16390
rect 16960 16250 16988 16526
rect 17130 16487 17132 16496
rect 17184 16487 17186 16496
rect 17132 16458 17184 16464
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 17144 15638 17172 16458
rect 17236 15638 17264 23462
rect 17788 23254 17816 23734
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17316 22976 17368 22982
rect 17316 22918 17368 22924
rect 17328 22506 17356 22918
rect 17788 22710 17816 23190
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17776 22704 17828 22710
rect 17776 22646 17828 22652
rect 17406 22536 17462 22545
rect 17316 22500 17368 22506
rect 17406 22471 17462 22480
rect 17316 22442 17368 22448
rect 17328 22030 17356 22442
rect 17420 22234 17448 22471
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17316 22024 17368 22030
rect 17420 22001 17448 22170
rect 17316 21966 17368 21972
rect 17406 21992 17462 22001
rect 17328 21350 17356 21966
rect 17406 21927 17462 21936
rect 17316 21344 17368 21350
rect 17316 21286 17368 21292
rect 17512 21010 17540 22646
rect 17776 22092 17828 22098
rect 17776 22034 17828 22040
rect 17788 21690 17816 22034
rect 17776 21684 17828 21690
rect 17776 21626 17828 21632
rect 17776 21344 17828 21350
rect 17776 21286 17828 21292
rect 17788 21010 17816 21286
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17512 20602 17540 20946
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17512 19446 17540 20538
rect 17788 19922 17816 20946
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17500 19440 17552 19446
rect 17500 19382 17552 19388
rect 17774 19272 17830 19281
rect 17774 19207 17776 19216
rect 17828 19207 17830 19216
rect 17776 19178 17828 19184
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17512 17338 17540 17682
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17880 16017 17908 27390
rect 18248 23730 18276 27520
rect 18696 25424 18748 25430
rect 18696 25366 18748 25372
rect 18708 24750 18736 25366
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18524 23497 18552 24550
rect 18604 24336 18656 24342
rect 18604 24278 18656 24284
rect 18616 23662 18644 24278
rect 18708 24138 18736 24686
rect 18696 24132 18748 24138
rect 18696 24074 18748 24080
rect 18604 23656 18656 23662
rect 18602 23624 18604 23633
rect 18656 23624 18658 23633
rect 18602 23559 18658 23568
rect 18696 23588 18748 23594
rect 18696 23530 18748 23536
rect 18510 23488 18566 23497
rect 18510 23423 18566 23432
rect 18708 23322 18736 23530
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18892 23225 18920 27520
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19156 24608 19208 24614
rect 19156 24550 19208 24556
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19076 23526 19104 24142
rect 19168 23769 19196 24550
rect 19154 23760 19210 23769
rect 19154 23695 19210 23704
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18972 23248 19024 23254
rect 18878 23216 18934 23225
rect 18972 23190 19024 23196
rect 18878 23151 18934 23160
rect 17960 22772 18012 22778
rect 17960 22714 18012 22720
rect 17972 21554 18000 22714
rect 18984 22438 19012 23190
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17972 20466 18000 21286
rect 18340 21185 18368 21830
rect 18892 21690 18920 21966
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18326 21176 18382 21185
rect 18892 21146 18920 21626
rect 18326 21111 18382 21120
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18892 20398 18920 21082
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18892 20058 18920 20334
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18328 19984 18380 19990
rect 18328 19926 18380 19932
rect 18340 19446 18368 19926
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18432 19514 18460 19790
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 18340 19310 18368 19382
rect 18800 19378 18828 19722
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17972 17678 18000 18022
rect 18064 17746 18092 18566
rect 18156 17882 18184 19178
rect 18708 18630 18736 19178
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18800 18193 18828 19314
rect 18786 18184 18842 18193
rect 18786 18119 18842 18128
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17972 17338 18000 17614
rect 18156 17354 18184 17818
rect 17960 17332 18012 17338
rect 18156 17326 18276 17354
rect 17960 17274 18012 17280
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 17866 16008 17922 16017
rect 17866 15943 17922 15952
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17776 15564 17828 15570
rect 17776 15506 17828 15512
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 17788 15162 17816 15506
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16868 14550 16896 14758
rect 16856 14544 16908 14550
rect 16856 14486 16908 14492
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16580 14476 16632 14482
rect 16408 14436 16580 14464
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 16408 13530 16436 14436
rect 16580 14418 16632 14424
rect 16960 14074 16988 14486
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16500 12986 16528 13738
rect 16764 13728 16816 13734
rect 16764 13670 16816 13676
rect 16776 13462 16804 13670
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16776 12850 16804 13398
rect 16868 13326 16896 14010
rect 16960 13870 16988 14010
rect 17328 14006 17356 14350
rect 17316 14000 17368 14006
rect 17316 13942 17368 13948
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12986 16896 13262
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16946 12880 17002 12889
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16764 12844 16816 12850
rect 16946 12815 17002 12824
rect 16764 12786 16816 12792
rect 16684 12714 16712 12786
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12640 16632 12646
rect 16500 12588 16580 12594
rect 16500 12582 16632 12588
rect 16500 12566 16620 12582
rect 16500 12374 16528 12566
rect 16776 12442 16804 12786
rect 16854 12744 16910 12753
rect 16960 12714 16988 12815
rect 16854 12679 16856 12688
rect 16908 12679 16910 12688
rect 16948 12708 17000 12714
rect 16856 12650 16908 12656
rect 16948 12650 17000 12656
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 18156 8401 18184 17206
rect 18248 17066 18276 17326
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18340 16402 18368 17274
rect 18708 17202 18736 18022
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18696 17060 18748 17066
rect 18696 17002 18748 17008
rect 18708 16794 18736 17002
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18800 16726 18828 18119
rect 18984 16833 19012 22374
rect 19076 20505 19104 23462
rect 19062 20496 19118 20505
rect 19062 20431 19118 20440
rect 19076 19961 19104 20431
rect 19062 19952 19118 19961
rect 19062 19887 19118 19896
rect 19064 19304 19116 19310
rect 19062 19272 19064 19281
rect 19116 19272 19118 19281
rect 19062 19207 19118 19216
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18420 16448 18472 16454
rect 18340 16396 18420 16402
rect 18340 16390 18472 16396
rect 18340 16374 18460 16390
rect 18616 16114 18644 16594
rect 18800 16250 18828 16662
rect 18880 16584 18932 16590
rect 19168 16561 19196 23598
rect 19352 23066 19380 25094
rect 19444 24954 19472 25230
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19536 24721 19564 27520
rect 19984 26444 20036 26450
rect 19984 26386 20036 26392
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19616 25288 19668 25294
rect 19616 25230 19668 25236
rect 19628 24886 19656 25230
rect 19616 24880 19668 24886
rect 19616 24822 19668 24828
rect 19522 24712 19578 24721
rect 19996 24698 20024 26386
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19720 24682 20024 24698
rect 19522 24647 19578 24656
rect 19708 24676 20024 24682
rect 19760 24670 20024 24676
rect 19708 24618 19760 24624
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19628 23662 19656 24006
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 20088 23254 20116 24822
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20180 24070 20208 24618
rect 20272 24410 20300 27520
rect 20352 26988 20404 26994
rect 20352 26930 20404 26936
rect 20260 24404 20312 24410
rect 20260 24346 20312 24352
rect 20168 24064 20220 24070
rect 20166 24032 20168 24041
rect 20220 24032 20222 24041
rect 20166 23967 20222 23976
rect 20364 23322 20392 26930
rect 20916 23866 20944 27520
rect 21560 25498 21588 27520
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 21364 24268 21416 24274
rect 21364 24210 21416 24216
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 20536 23792 20588 23798
rect 20536 23734 20588 23740
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 19892 23248 19944 23254
rect 19892 23190 19944 23196
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 19524 23180 19576 23186
rect 19524 23122 19576 23128
rect 19352 23038 19472 23066
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 18880 16526 18932 16532
rect 19154 16552 19210 16561
rect 18892 16250 18920 16526
rect 19154 16487 19210 16496
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19076 15026 19104 15438
rect 19168 15162 19196 16390
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14521 19104 14758
rect 19168 14550 19196 15098
rect 19156 14544 19208 14550
rect 19062 14512 19118 14521
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18604 14476 18656 14482
rect 19156 14486 19208 14492
rect 19062 14447 19118 14456
rect 18604 14418 18656 14424
rect 18340 14074 18368 14418
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18616 14006 18644 14418
rect 18236 14000 18288 14006
rect 18236 13942 18288 13948
rect 18604 14000 18656 14006
rect 18604 13942 18656 13948
rect 18248 13530 18276 13942
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18142 8392 18198 8401
rect 18142 8327 18198 8336
rect 19260 3505 19288 21558
rect 19352 21486 19380 22918
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19444 21418 19472 23038
rect 19536 22234 19564 23122
rect 19904 22778 19932 23190
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 19904 22506 19932 22714
rect 20548 22574 20576 23734
rect 21376 23526 21404 24210
rect 20720 23520 20772 23526
rect 20640 23468 20720 23474
rect 20640 23462 20772 23468
rect 21364 23520 21416 23526
rect 22204 23474 22232 27520
rect 22940 24614 22968 27520
rect 23110 27160 23166 27169
rect 23110 27095 23166 27104
rect 22376 24608 22428 24614
rect 22376 24550 22428 24556
rect 22928 24608 22980 24614
rect 22928 24550 22980 24556
rect 21364 23462 21416 23468
rect 20640 23446 20760 23462
rect 20640 23254 20668 23446
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 19892 22500 19944 22506
rect 19944 22460 20024 22488
rect 19892 22442 19944 22448
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19524 22228 19576 22234
rect 19524 22170 19576 22176
rect 19996 22166 20024 22460
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19432 21412 19484 21418
rect 19432 21354 19484 21360
rect 19444 21146 19472 21354
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19432 21140 19484 21146
rect 19432 21082 19484 21088
rect 19430 20360 19486 20369
rect 19430 20295 19486 20304
rect 20444 20324 20496 20330
rect 19444 20262 19472 20295
rect 20444 20266 20496 20272
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 20456 20058 20484 20266
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20548 19922 20576 22510
rect 20628 22432 20680 22438
rect 20628 22374 20680 22380
rect 20640 21554 20668 22374
rect 20916 22234 20944 23122
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20916 21146 20944 22170
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20262 20760 20742
rect 20916 20602 20944 20946
rect 21376 20641 21404 23462
rect 22020 23446 22232 23474
rect 22020 23322 22048 23446
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22296 22778 22324 23054
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22100 22704 22152 22710
rect 21822 22672 21878 22681
rect 21822 22607 21824 22616
rect 21876 22607 21878 22616
rect 22020 22652 22100 22658
rect 22020 22646 22152 22652
rect 22020 22630 22140 22646
rect 21824 22578 21876 22584
rect 22020 22114 22048 22630
rect 22100 22160 22152 22166
rect 22020 22108 22100 22114
rect 22020 22102 22152 22108
rect 22020 22086 22140 22102
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21744 21350 21772 21830
rect 22020 21690 22048 22086
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21362 20632 21418 20641
rect 20904 20596 20956 20602
rect 21362 20567 21418 20576
rect 20904 20538 20956 20544
rect 22388 20369 22416 24550
rect 23020 24268 23072 24274
rect 23020 24210 23072 24216
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22756 23866 22784 24142
rect 23032 23866 23060 24210
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 22466 23760 22522 23769
rect 22466 23695 22522 23704
rect 22480 22506 22508 23695
rect 22928 23248 22980 23254
rect 23124 23202 23152 27095
rect 23584 25498 23612 27520
rect 23938 26072 23994 26081
rect 23938 26007 23994 26016
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23204 25356 23256 25362
rect 23204 25298 23256 25304
rect 23216 24614 23244 25298
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23570 24848 23626 24857
rect 23570 24783 23626 24792
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 22928 23190 22980 23196
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22848 23089 22876 23122
rect 22834 23080 22890 23089
rect 22834 23015 22890 23024
rect 22560 22976 22612 22982
rect 22560 22918 22612 22924
rect 22468 22500 22520 22506
rect 22468 22442 22520 22448
rect 22480 22098 22508 22442
rect 22572 22098 22600 22918
rect 22940 22778 22968 23190
rect 23032 23174 23152 23202
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22940 22545 22968 22714
rect 22926 22536 22982 22545
rect 22926 22471 22982 22480
rect 23032 22234 23060 23174
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23124 22506 23152 23054
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 23020 22228 23072 22234
rect 23020 22170 23072 22176
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 23020 22092 23072 22098
rect 23020 22034 23072 22040
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22480 21078 22508 21490
rect 22572 21146 22600 22034
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22928 22024 22980 22030
rect 22928 21966 22980 21972
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22652 20936 22704 20942
rect 22652 20878 22704 20884
rect 22664 20754 22692 20878
rect 22756 20874 22784 21286
rect 22744 20868 22796 20874
rect 22744 20810 22796 20816
rect 22664 20726 22784 20754
rect 22374 20360 22430 20369
rect 21180 20324 21232 20330
rect 22374 20295 22430 20304
rect 21180 20266 21232 20272
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 19310 20576 19858
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19720 17066 19748 17478
rect 20548 17338 20576 19246
rect 20732 18698 20760 20198
rect 21192 20058 21220 20266
rect 22756 20262 22784 20726
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 22008 19984 22060 19990
rect 22008 19926 22060 19932
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21454 19408 21510 19417
rect 21454 19343 21510 19352
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 21376 18086 21404 18838
rect 21468 18766 21496 19343
rect 21836 19242 21864 19858
rect 22020 19514 22048 19926
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21652 18766 21680 19178
rect 21836 18970 21864 19178
rect 22112 19174 22140 19450
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21824 18964 21876 18970
rect 21824 18906 21876 18912
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21468 18426 21496 18702
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21652 18086 21680 18702
rect 22756 18193 22784 20198
rect 22742 18184 22798 18193
rect 22742 18119 22798 18128
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 20536 17332 20588 17338
rect 20536 17274 20588 17280
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 19708 17060 19760 17066
rect 19708 17002 19760 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 20548 16454 20576 17274
rect 21100 16726 21128 17274
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20536 16448 20588 16454
rect 20536 16390 20588 16396
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16250 21036 16390
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 21008 15502 21036 16186
rect 21100 15706 21128 16662
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 20168 15360 20220 15366
rect 20168 15302 20220 15308
rect 20180 14890 20208 15302
rect 21270 15056 21326 15065
rect 21270 14991 21326 15000
rect 20168 14884 20220 14890
rect 20168 14826 20220 14832
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19812 13870 19840 14214
rect 20916 14074 20944 14826
rect 21284 14550 21312 14991
rect 21376 14618 21404 18022
rect 21456 17808 21508 17814
rect 21454 17776 21456 17785
rect 21508 17776 21510 17785
rect 21454 17711 21510 17720
rect 21468 17202 21496 17711
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21560 17338 21588 17614
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 21456 17196 21508 17202
rect 21456 17138 21508 17144
rect 21652 15162 21680 18022
rect 22848 17746 22876 21966
rect 22940 21486 22968 21966
rect 23032 21554 23060 22034
rect 23124 21622 23152 22442
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23020 21548 23072 21554
rect 23020 21490 23072 21496
rect 22928 21480 22980 21486
rect 22928 21422 22980 21428
rect 23124 21418 23152 21558
rect 23216 21486 23244 24550
rect 23388 23860 23440 23866
rect 23388 23802 23440 23808
rect 23296 23588 23348 23594
rect 23296 23530 23348 23536
rect 23308 22250 23336 23530
rect 23400 22710 23428 23802
rect 23480 23316 23532 23322
rect 23480 23258 23532 23264
rect 23492 23225 23520 23258
rect 23584 23254 23612 24783
rect 23572 23248 23624 23254
rect 23478 23216 23534 23225
rect 23572 23190 23624 23196
rect 23478 23151 23534 23160
rect 23478 23080 23534 23089
rect 23478 23015 23534 23024
rect 23492 22778 23520 23015
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 23480 22432 23532 22438
rect 23480 22374 23532 22380
rect 23308 22222 23428 22250
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23124 21146 23152 21354
rect 23308 21332 23336 22102
rect 23400 21842 23428 22222
rect 23492 21962 23520 22374
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23400 21814 23520 21842
rect 23492 21570 23520 21814
rect 23584 21690 23612 22578
rect 23676 22409 23704 24890
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23662 22400 23718 22409
rect 23662 22335 23718 22344
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 23676 21962 23704 22170
rect 23664 21956 23716 21962
rect 23664 21898 23716 21904
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23492 21542 23612 21570
rect 23388 21480 23440 21486
rect 23388 21422 23440 21428
rect 23216 21304 23336 21332
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23020 21072 23072 21078
rect 23020 21014 23072 21020
rect 23032 20262 23060 21014
rect 23124 20602 23152 21082
rect 23216 21078 23244 21304
rect 23204 21072 23256 21078
rect 23204 21014 23256 21020
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23032 19281 23060 20198
rect 23124 20058 23152 20538
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23018 19272 23074 19281
rect 23018 19207 23074 19216
rect 23400 19145 23428 21422
rect 23386 19136 23442 19145
rect 23386 19071 23442 19080
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23492 18426 23520 18770
rect 23584 18737 23612 21542
rect 23664 21480 23716 21486
rect 23664 21422 23716 21428
rect 23676 20806 23704 21422
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 19174 23704 20742
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23676 18766 23704 19110
rect 23664 18760 23716 18766
rect 23570 18728 23626 18737
rect 23664 18702 23716 18708
rect 23570 18663 23626 18672
rect 23676 18578 23704 18702
rect 23584 18550 23704 18578
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 22836 17740 22888 17746
rect 22836 17682 22888 17688
rect 21824 17604 21876 17610
rect 21824 17546 21876 17552
rect 21836 16998 21864 17546
rect 21916 17536 21968 17542
rect 21916 17478 21968 17484
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21836 16697 21864 16934
rect 21822 16688 21878 16697
rect 21822 16623 21878 16632
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21272 14544 21324 14550
rect 20994 14512 21050 14521
rect 21272 14486 21324 14492
rect 20994 14447 21050 14456
rect 21008 14346 21036 14447
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21284 14074 21312 14486
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 19616 13864 19668 13870
rect 19536 13812 19616 13818
rect 19536 13806 19668 13812
rect 19800 13864 19852 13870
rect 19800 13806 19852 13812
rect 19536 13790 19656 13806
rect 19536 13530 19564 13790
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 21376 13530 21404 14554
rect 21548 14408 21600 14414
rect 21548 14350 21600 14356
rect 21560 14278 21588 14350
rect 21548 14272 21600 14278
rect 21548 14214 21600 14220
rect 21560 14074 21588 14214
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21364 13524 21416 13530
rect 21364 13466 21416 13472
rect 21192 12889 21220 13466
rect 21362 13424 21418 13433
rect 21362 13359 21418 13368
rect 21376 12889 21404 13359
rect 21178 12880 21234 12889
rect 21178 12815 21234 12824
rect 21362 12880 21418 12889
rect 21362 12815 21418 12824
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19338 8392 19394 8401
rect 19338 8327 19394 8336
rect 19352 7954 19380 8327
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 21836 7954 21864 16118
rect 21928 15978 21956 17478
rect 22848 17338 22876 17682
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 23216 17134 23244 17750
rect 23204 17128 23256 17134
rect 23202 17096 23204 17105
rect 23256 17096 23258 17105
rect 23202 17031 23258 17040
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22020 16114 22048 16934
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21928 15706 21956 15914
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 22020 15638 22048 16050
rect 22388 15978 22416 16390
rect 23124 16250 23152 16662
rect 23400 16658 23428 18022
rect 23492 17626 23520 18362
rect 23584 18086 23612 18550
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23492 17598 23612 17626
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23388 16652 23440 16658
rect 23388 16594 23440 16600
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 22848 15570 22876 15914
rect 23124 15706 23152 16186
rect 23492 15978 23520 17478
rect 23584 16250 23612 17598
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23480 15972 23532 15978
rect 23480 15914 23532 15920
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22560 15496 22612 15502
rect 22560 15438 22612 15444
rect 22572 15162 22600 15438
rect 22848 15162 22876 15506
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 23676 9042 23704 18294
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22928 7948 22980 7954
rect 22928 7890 22980 7896
rect 19352 7546 19380 7890
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 19340 7540 19392 7546
rect 19340 7482 19392 7488
rect 19628 7449 19656 7822
rect 22940 7546 22968 7890
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 19614 7440 19670 7449
rect 19614 7375 19670 7384
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23492 6497 23520 6802
rect 23478 6488 23534 6497
rect 23478 6423 23480 6432
rect 23532 6423 23534 6432
rect 23480 6394 23532 6400
rect 23662 6352 23718 6361
rect 23662 6287 23718 6296
rect 23676 6254 23704 6287
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 23662 5808 23718 5817
rect 23662 5743 23664 5752
rect 23716 5743 23718 5752
rect 23664 5714 23716 5720
rect 23676 5370 23704 5714
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23664 5160 23716 5166
rect 23662 5128 23664 5137
rect 23716 5128 23718 5137
rect 23662 5063 23718 5072
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 19246 3496 19302 3505
rect 19246 3431 19302 3440
rect 23492 3126 23520 3538
rect 23768 3194 23796 22646
rect 23860 22574 23888 23122
rect 23952 23089 23980 26007
rect 24228 24682 24256 27520
rect 24780 26994 24808 27639
rect 24858 27520 24914 28000
rect 25594 27520 25650 28000
rect 26238 27520 26294 28000
rect 26882 27520 26938 28000
rect 27526 27520 27582 28000
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24766 26616 24822 26625
rect 24766 26551 24822 26560
rect 24780 26450 24808 26551
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24674 25392 24730 25401
rect 24674 25327 24730 25336
rect 24768 25356 24820 25362
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24886 24716 25327
rect 24768 25298 24820 25304
rect 24780 24954 24808 25298
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24676 24880 24728 24886
rect 24872 24834 24900 27520
rect 24676 24822 24728 24828
rect 24780 24806 24900 24834
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 23938 23080 23994 23089
rect 23938 23015 23994 23024
rect 23940 22976 23992 22982
rect 23940 22918 23992 22924
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23860 19394 23888 22510
rect 23952 22506 23980 22918
rect 24044 22522 24072 24550
rect 24214 24304 24270 24313
rect 24214 24239 24270 24248
rect 24124 24064 24176 24070
rect 24122 24032 24124 24041
rect 24176 24032 24178 24041
rect 24122 23967 24178 23976
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24136 22642 24164 22918
rect 24228 22658 24256 24239
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24674 23896 24730 23905
rect 24674 23831 24676 23840
rect 24728 23831 24730 23840
rect 24676 23802 24728 23808
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24124 22636 24176 22642
rect 24228 22630 24440 22658
rect 24124 22578 24176 22584
rect 23940 22500 23992 22506
rect 24044 22494 24164 22522
rect 23940 22442 23992 22448
rect 23938 22400 23994 22409
rect 23938 22335 23994 22344
rect 23952 20913 23980 22335
rect 24030 21992 24086 22001
rect 24030 21927 24086 21936
rect 23938 20904 23994 20913
rect 23938 20839 23994 20848
rect 24044 20505 24072 21927
rect 24136 21457 24164 22494
rect 24216 22092 24268 22098
rect 24216 22034 24268 22040
rect 24122 21448 24178 21457
rect 24122 21383 24178 21392
rect 24228 21350 24256 22034
rect 24412 22001 24440 22630
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24504 22234 24532 22578
rect 24492 22228 24544 22234
rect 24492 22170 24544 22176
rect 24398 21992 24454 22001
rect 24398 21927 24454 21936
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24228 21146 24256 21286
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24122 20632 24178 20641
rect 24289 20624 24585 20644
rect 24122 20567 24178 20576
rect 24030 20496 24086 20505
rect 24030 20431 24086 20440
rect 24044 20058 24072 20431
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 23952 19553 23980 19926
rect 24044 19922 24072 19994
rect 24032 19916 24084 19922
rect 24032 19858 24084 19864
rect 23938 19544 23994 19553
rect 23938 19479 23940 19488
rect 23992 19479 23994 19488
rect 23940 19450 23992 19456
rect 23860 19366 23980 19394
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23860 17066 23888 17614
rect 23848 17060 23900 17066
rect 23848 17002 23900 17008
rect 23952 16833 23980 19366
rect 24030 18184 24086 18193
rect 24030 18119 24086 18128
rect 24044 17898 24072 18119
rect 24136 18057 24164 20567
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24122 18048 24178 18057
rect 24122 17983 24178 17992
rect 24044 17870 24164 17898
rect 24032 17264 24084 17270
rect 24032 17206 24084 17212
rect 23938 16824 23994 16833
rect 23938 16759 23994 16768
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23860 8430 23888 16118
rect 24044 16046 24072 17206
rect 24136 16998 24164 17870
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 24228 17202 24256 17614
rect 24688 17513 24716 23666
rect 24780 21146 24808 24806
rect 25410 24712 25466 24721
rect 25410 24647 25466 24656
rect 25424 24410 25452 24647
rect 25412 24404 25464 24410
rect 25412 24346 25464 24352
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25240 23730 25268 24210
rect 25228 23724 25280 23730
rect 25228 23666 25280 23672
rect 25228 23520 25280 23526
rect 25226 23488 25228 23497
rect 25280 23488 25282 23497
rect 25226 23423 25282 23432
rect 25608 22778 25636 27520
rect 26252 23905 26280 27520
rect 26238 23896 26294 23905
rect 26238 23831 26294 23840
rect 26896 23202 26924 27520
rect 26252 23174 26924 23202
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25870 22536 25926 22545
rect 25870 22471 25872 22480
rect 25924 22471 25926 22480
rect 25872 22442 25924 22448
rect 25042 21992 25098 22001
rect 25042 21927 25098 21936
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 25056 21010 25084 21927
rect 25044 21004 25096 21010
rect 25044 20946 25096 20952
rect 25056 20602 25084 20946
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24780 18578 24808 20198
rect 25148 19854 25176 20266
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24780 18550 24900 18578
rect 24872 18290 24900 18550
rect 24860 18284 24912 18290
rect 24860 18226 24912 18232
rect 24872 18034 24900 18226
rect 24964 18154 24992 19654
rect 25148 19242 25176 19790
rect 26252 19310 26280 23174
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 25136 19236 25188 19242
rect 25136 19178 25188 19184
rect 25148 18970 25176 19178
rect 25136 18964 25188 18970
rect 25136 18906 25188 18912
rect 24952 18148 25004 18154
rect 24952 18090 25004 18096
rect 24780 18006 24900 18034
rect 24780 17882 24808 18006
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24674 17504 24730 17513
rect 24289 17436 24585 17456
rect 24674 17439 24730 17448
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 16794 24164 16934
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24032 16040 24084 16046
rect 24032 15982 24084 15988
rect 23848 8424 23900 8430
rect 23848 8366 23900 8372
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23860 4690 23888 5646
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23860 4282 23888 4626
rect 23848 4276 23900 4282
rect 23848 4218 23900 4224
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23480 3120 23532 3126
rect 16118 3088 16174 3097
rect 16118 3023 16174 3032
rect 23478 3088 23480 3097
rect 23532 3088 23534 3097
rect 23952 3058 23980 4014
rect 23478 3023 23534 3032
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 23664 2984 23716 2990
rect 23662 2952 23664 2961
rect 23716 2952 23718 2961
rect 22560 2916 22612 2922
rect 23662 2887 23718 2896
rect 22560 2858 22612 2864
rect 22572 2825 22600 2858
rect 22558 2816 22614 2825
rect 19622 2748 19918 2768
rect 22558 2751 22614 2760
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 2417 24072 2450
rect 16026 2408 16082 2417
rect 16026 2343 16082 2352
rect 24030 2408 24086 2417
rect 24030 2343 24086 2352
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 23032 2009 23060 2246
rect 23018 2000 23074 2009
rect 23018 1935 23074 1944
rect 14002 0 14058 480
rect 24136 377 24164 16730
rect 24412 16726 24440 17002
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24400 16720 24452 16726
rect 24872 16674 24900 16730
rect 24400 16662 24452 16668
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 24780 16646 24900 16674
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24688 16182 24716 16594
rect 24780 16250 24808 16646
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 25226 16008 25282 16017
rect 24216 15972 24268 15978
rect 25226 15943 25282 15952
rect 24216 15914 24268 15920
rect 24228 15706 24256 15914
rect 25042 15736 25098 15745
rect 24216 15700 24268 15706
rect 25240 15706 25268 15943
rect 25042 15671 25098 15680
rect 25228 15700 25280 15706
rect 24216 15642 24268 15648
rect 25056 15570 25084 15671
rect 25228 15642 25280 15648
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 25056 15162 25084 15506
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 24766 14920 24822 14929
rect 24766 14855 24822 14864
rect 24582 14648 24638 14657
rect 24780 14618 24808 14855
rect 24582 14583 24638 14592
rect 24768 14612 24820 14618
rect 24596 14482 24624 14583
rect 24768 14554 24820 14560
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24596 14362 24624 14418
rect 24596 14334 24716 14362
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24688 14074 24716 14334
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 24214 13968 24270 13977
rect 24214 13903 24270 13912
rect 24228 12753 24256 13903
rect 24582 13424 24638 13433
rect 24582 13359 24584 13368
rect 24636 13359 24638 13368
rect 24584 13330 24636 13336
rect 24596 13274 24624 13330
rect 24766 13288 24822 13297
rect 24596 13246 24716 13274
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24688 12986 24716 13246
rect 24766 13223 24768 13232
rect 24820 13223 24822 13232
rect 24768 13194 24820 13200
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24214 12744 24270 12753
rect 24214 12679 24270 12688
rect 25332 12442 25360 19246
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25516 18873 25544 19110
rect 27540 18873 27568 27520
rect 25502 18864 25558 18873
rect 25502 18799 25558 18808
rect 27526 18864 27582 18873
rect 27526 18799 27582 18808
rect 25516 18290 25544 18799
rect 25504 18284 25556 18290
rect 25504 18226 25556 18232
rect 25410 16552 25466 16561
rect 25410 16487 25466 16496
rect 25424 16250 25452 16487
rect 25870 16280 25926 16289
rect 25412 16244 25464 16250
rect 25870 16215 25872 16224
rect 25412 16186 25464 16192
rect 25924 16215 25926 16224
rect 25872 16186 25924 16192
rect 25884 16046 25912 16186
rect 25872 16040 25924 16046
rect 25872 15982 25924 15988
rect 25320 12436 25372 12442
rect 25320 12378 25372 12384
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24596 12209 24624 12242
rect 24582 12200 24638 12209
rect 24638 12158 24716 12186
rect 24582 12135 24638 12144
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24688 11898 24716 12158
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24584 9512 24636 9518
rect 24584 9454 24636 9460
rect 24596 9110 24624 9454
rect 24768 9376 24820 9382
rect 24768 9318 24820 9324
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24780 8265 24808 9318
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24964 8634 24992 8978
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 24766 8256 24822 8265
rect 24766 8191 24822 8200
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24228 7546 24256 7890
rect 24768 7744 24820 7750
rect 25332 7721 25360 8502
rect 24768 7686 24820 7692
rect 25318 7712 25374 7721
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24582 7440 24638 7449
rect 24582 7375 24638 7384
rect 24596 7342 24624 7375
rect 24584 7336 24636 7342
rect 24584 7278 24636 7284
rect 24676 7200 24728 7206
rect 24780 7177 24808 7686
rect 25318 7647 25374 7656
rect 24676 7142 24728 7148
rect 24766 7168 24822 7177
rect 24688 6633 24716 7142
rect 24766 7103 24822 7112
rect 24768 6860 24820 6866
rect 24768 6802 24820 6808
rect 24674 6624 24730 6633
rect 24289 6556 24585 6576
rect 24674 6559 24730 6568
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24780 6458 24808 6802
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24950 6216 25006 6225
rect 24950 6151 25006 6160
rect 24964 5778 24992 6151
rect 25148 6089 25176 6598
rect 26148 6112 26200 6118
rect 25134 6080 25190 6089
rect 26148 6054 26200 6060
rect 25134 6015 25190 6024
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24964 5370 24992 5714
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25148 5409 25176 5510
rect 25134 5400 25190 5409
rect 24952 5364 25004 5370
rect 25134 5335 25190 5344
rect 24952 5306 25004 5312
rect 25136 5024 25188 5030
rect 25136 4966 25188 4972
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 24228 4162 24256 4626
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4321 24716 4422
rect 24674 4312 24730 4321
rect 24674 4247 24730 4256
rect 24228 4134 24440 4162
rect 24216 4004 24268 4010
rect 24216 3946 24268 3952
rect 24228 2553 24256 3946
rect 24412 3942 24440 4134
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 24412 3670 24440 3878
rect 24400 3664 24452 3670
rect 24400 3606 24452 3612
rect 24780 3482 24808 4422
rect 25148 3777 25176 4966
rect 26160 4865 26188 6054
rect 26146 4856 26202 4865
rect 26146 4791 26202 4800
rect 25134 3768 25190 3777
rect 25134 3703 25190 3712
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 24688 3454 24808 3482
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24688 3233 24716 3454
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24674 3224 24730 3233
rect 24674 3159 24730 3168
rect 24214 2544 24270 2553
rect 24214 2479 24270 2488
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24780 1465 24808 3334
rect 24872 3194 24900 3538
rect 24950 3496 25006 3505
rect 24950 3431 25006 3440
rect 24860 3188 24912 3194
rect 24860 3130 24912 3136
rect 24964 2990 24992 3431
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 25318 2816 25374 2825
rect 25318 2751 25374 2760
rect 25332 2514 25360 2751
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25504 2304 25556 2310
rect 25504 2246 25556 2252
rect 24766 1456 24822 1465
rect 24766 1391 24822 1400
rect 25516 921 25544 2246
rect 25502 912 25558 921
rect 25502 847 25558 856
rect 24122 368 24178 377
rect 24122 303 24178 312
<< via2 >>
rect 24766 27648 24822 27704
rect 938 23568 994 23624
rect 1582 22480 1638 22536
rect 2226 19760 2282 19816
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5538 24656 5594 24712
rect 4894 24112 4950 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 4250 23704 4306 23760
rect 6274 23024 6330 23080
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6918 19216 6974 19272
rect 3606 18808 3662 18864
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 7562 17720 7618 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 2870 17176 2926 17232
rect 8942 19352 8998 19408
rect 8206 17040 8262 17096
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 3330 15952 3386 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 3330 14048 3386 14104
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 386 12688 442 12744
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9954 23704 10010 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 9862 8900 9918 8936
rect 9862 8880 9864 8900
rect 9864 8880 9916 8900
rect 9916 8880 9918 8900
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 9954 6296 10010 6352
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10874 21972 10876 21992
rect 10876 21972 10928 21992
rect 10928 21972 10930 21992
rect 10874 21936 10930 21972
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10138 18808 10194 18864
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10690 16652 10746 16688
rect 10690 16632 10692 16652
rect 10692 16632 10744 16652
rect 10744 16632 10746 16652
rect 10690 15952 10746 16008
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 11150 16496 11206 16552
rect 12162 24112 12218 24168
rect 12990 23724 13046 23760
rect 12990 23704 12992 23724
rect 12992 23704 13044 23724
rect 13044 23704 13046 23724
rect 12898 19760 12954 19816
rect 12806 16632 12862 16688
rect 14002 24676 14058 24712
rect 14002 24656 14004 24676
rect 14004 24656 14056 24676
rect 14056 24656 14058 24676
rect 14094 23432 14150 23488
rect 13634 23024 13690 23080
rect 13542 22616 13598 22672
rect 13450 19896 13506 19952
rect 13726 20984 13782 21040
rect 13726 20340 13728 20360
rect 13728 20340 13780 20360
rect 13780 20340 13782 20360
rect 13726 20304 13782 20340
rect 14370 23296 14426 23352
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 12898 11600 12954 11656
rect 12254 11076 12310 11112
rect 12254 11056 12256 11076
rect 12256 11056 12308 11076
rect 12308 11056 12310 11076
rect 11426 10512 11482 10568
rect 10230 9424 10286 9480
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10046 5752 10102 5808
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 10874 9988 10930 10024
rect 10874 9968 10876 9988
rect 10876 9968 10928 9988
rect 10928 9968 10930 9988
rect 13358 8200 13414 8256
rect 10782 5072 10838 5128
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 14186 13368 14242 13424
rect 14002 12688 14058 12744
rect 14370 13232 14426 13288
rect 14002 8200 14058 8256
rect 13450 2896 13506 2952
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15474 20984 15530 21040
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15014 16768 15070 16824
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 16118 22500 16174 22536
rect 16118 22480 16120 22500
rect 16120 22480 16172 22500
rect 16172 22480 16174 22500
rect 15382 6432 15438 6488
rect 15198 6180 15254 6216
rect 15198 6160 15200 6180
rect 15200 6160 15252 6180
rect 15252 6160 15254 6180
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 16118 17212 16120 17232
rect 16120 17212 16172 17232
rect 16172 17212 16174 17232
rect 16118 17176 16174 17212
rect 17038 23296 17094 23352
rect 16762 21936 16818 21992
rect 16486 21140 16542 21176
rect 16486 21120 16488 21140
rect 16488 21120 16540 21140
rect 16540 21120 16542 21140
rect 16578 20304 16634 20360
rect 16210 15000 16266 15056
rect 17130 16516 17186 16552
rect 17130 16496 17132 16516
rect 17132 16496 17184 16516
rect 17184 16496 17186 16516
rect 17406 22480 17462 22536
rect 17406 21936 17462 21992
rect 17774 19236 17830 19272
rect 17774 19216 17776 19236
rect 17776 19216 17828 19236
rect 17828 19216 17830 19236
rect 18602 23604 18604 23624
rect 18604 23604 18656 23624
rect 18656 23604 18658 23624
rect 18602 23568 18658 23604
rect 18510 23432 18566 23488
rect 19154 23704 19210 23760
rect 18878 23160 18934 23216
rect 18326 21120 18382 21176
rect 18786 18128 18842 18184
rect 17866 15952 17922 16008
rect 16946 12824 17002 12880
rect 16854 12708 16910 12744
rect 16854 12688 16856 12708
rect 16856 12688 16908 12708
rect 16908 12688 16910 12708
rect 19062 20440 19118 20496
rect 19062 19896 19118 19952
rect 19062 19252 19064 19272
rect 19064 19252 19116 19272
rect 19116 19252 19118 19272
rect 19062 19216 19118 19252
rect 18970 16768 19026 16824
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19522 24656 19578 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 20166 24012 20168 24032
rect 20168 24012 20220 24032
rect 20220 24012 20222 24032
rect 20166 23976 20222 24012
rect 19154 16496 19210 16552
rect 19062 14456 19118 14512
rect 18142 8336 18198 8392
rect 23110 27104 23166 27160
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19430 20304 19486 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 21822 22636 21878 22672
rect 21822 22616 21824 22636
rect 21824 22616 21876 22636
rect 21876 22616 21878 22636
rect 21362 20576 21418 20632
rect 22466 23704 22522 23760
rect 23938 26016 23994 26072
rect 23570 24792 23626 24848
rect 22834 23024 22890 23080
rect 22926 22480 22982 22536
rect 22374 20304 22430 20360
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 21454 19352 21510 19408
rect 22742 18128 22798 18184
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 21270 15000 21326 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 21454 17756 21456 17776
rect 21456 17756 21508 17776
rect 21508 17756 21510 17776
rect 21454 17720 21510 17756
rect 23478 23160 23534 23216
rect 23478 23024 23534 23080
rect 23662 22344 23718 22400
rect 23018 19216 23074 19272
rect 23386 19080 23442 19136
rect 23570 18672 23626 18728
rect 21822 16632 21878 16688
rect 20994 14456 21050 14512
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 21362 13368 21418 13424
rect 21178 12824 21234 12880
rect 21362 12824 21418 12880
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19338 8336 19394 8392
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 23202 17076 23204 17096
rect 23204 17076 23256 17096
rect 23256 17076 23258 17096
rect 23202 17040 23258 17076
rect 19614 7384 19670 7440
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 23478 6452 23534 6488
rect 23478 6432 23480 6452
rect 23480 6432 23532 6452
rect 23532 6432 23534 6452
rect 23662 6296 23718 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 23662 5772 23718 5808
rect 23662 5752 23664 5772
rect 23664 5752 23716 5772
rect 23716 5752 23718 5772
rect 23662 5108 23664 5128
rect 23664 5108 23716 5128
rect 23716 5108 23718 5128
rect 23662 5072 23718 5108
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19246 3440 19302 3496
rect 24766 26560 24822 26616
rect 24674 25336 24730 25392
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 23938 23024 23994 23080
rect 24214 24248 24270 24304
rect 24122 24012 24124 24032
rect 24124 24012 24176 24032
rect 24176 24012 24178 24032
rect 24122 23976 24178 24012
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24674 23860 24730 23896
rect 24674 23840 24676 23860
rect 24676 23840 24728 23860
rect 24728 23840 24730 23860
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23938 22344 23994 22400
rect 24030 21936 24086 21992
rect 23938 20848 23994 20904
rect 24122 21392 24178 21448
rect 24398 21936 24454 21992
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24122 20576 24178 20632
rect 24030 20440 24086 20496
rect 23938 19508 23994 19544
rect 23938 19488 23940 19508
rect 23940 19488 23992 19508
rect 23992 19488 23994 19508
rect 24030 18128 24086 18184
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24122 17992 24178 18048
rect 23938 16768 23994 16824
rect 25410 24656 25466 24712
rect 25226 23468 25228 23488
rect 25228 23468 25280 23488
rect 25280 23468 25282 23488
rect 25226 23432 25282 23468
rect 26238 23840 26294 23896
rect 25870 22500 25926 22536
rect 25870 22480 25872 22500
rect 25872 22480 25924 22500
rect 25924 22480 25926 22500
rect 25042 21936 25098 21992
rect 24674 17448 24730 17504
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 16118 3032 16174 3088
rect 23478 3068 23480 3088
rect 23480 3068 23532 3088
rect 23532 3068 23534 3088
rect 23478 3032 23534 3068
rect 23662 2932 23664 2952
rect 23664 2932 23716 2952
rect 23716 2932 23718 2952
rect 23662 2896 23718 2932
rect 22558 2760 22614 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 16026 2352 16082 2408
rect 24030 2352 24086 2408
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 23018 1944 23074 2000
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 25226 15952 25282 16008
rect 25042 15680 25098 15736
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24766 14864 24822 14920
rect 24582 14592 24638 14648
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24214 13912 24270 13968
rect 24582 13388 24638 13424
rect 24582 13368 24584 13388
rect 24584 13368 24636 13388
rect 24636 13368 24638 13388
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24766 13252 24822 13288
rect 24766 13232 24768 13252
rect 24768 13232 24820 13252
rect 24820 13232 24822 13252
rect 24214 12688 24270 12744
rect 25502 18808 25558 18864
rect 27526 18808 27582 18864
rect 25410 16496 25466 16552
rect 25870 16244 25926 16280
rect 25870 16224 25872 16244
rect 25872 16224 25924 16244
rect 25924 16224 25926 16244
rect 24582 12144 24638 12200
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24766 8200 24822 8256
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24582 7384 24638 7440
rect 25318 7656 25374 7712
rect 24766 7112 24822 7168
rect 24674 6568 24730 6624
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24950 6160 25006 6216
rect 25134 6024 25190 6080
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 25134 5344 25190 5400
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24674 4256 24730 4312
rect 26146 4800 26202 4856
rect 25134 3712 25190 3768
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24674 3168 24730 3224
rect 24214 2488 24270 2544
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24950 3440 25006 3496
rect 25318 2760 25374 2816
rect 24766 1400 24822 1456
rect 25502 856 25558 912
rect 24122 312 24178 368
<< metal3 >>
rect 24761 27706 24827 27709
rect 27520 27706 28000 27736
rect 24761 27704 28000 27706
rect 24761 27648 24766 27704
rect 24822 27648 28000 27704
rect 24761 27646 28000 27648
rect 24761 27643 24827 27646
rect 27520 27616 28000 27646
rect 23105 27162 23171 27165
rect 27520 27162 28000 27192
rect 23105 27160 28000 27162
rect 23105 27104 23110 27160
rect 23166 27104 28000 27160
rect 23105 27102 28000 27104
rect 23105 27099 23171 27102
rect 27520 27072 28000 27102
rect 24761 26618 24827 26621
rect 27520 26618 28000 26648
rect 24761 26616 28000 26618
rect 24761 26560 24766 26616
rect 24822 26560 28000 26616
rect 24761 26558 28000 26560
rect 24761 26555 24827 26558
rect 27520 26528 28000 26558
rect 23933 26074 23999 26077
rect 27520 26074 28000 26104
rect 23933 26072 28000 26074
rect 23933 26016 23938 26072
rect 23994 26016 28000 26072
rect 23933 26014 28000 26016
rect 23933 26011 23999 26014
rect 27520 25984 28000 26014
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 24669 25394 24735 25397
rect 27520 25394 28000 25424
rect 24669 25392 28000 25394
rect 24669 25336 24674 25392
rect 24730 25336 28000 25392
rect 24669 25334 28000 25336
rect 24669 25331 24735 25334
rect 27520 25304 28000 25334
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 23565 24850 23631 24853
rect 27520 24850 28000 24880
rect 23565 24848 28000 24850
rect 23565 24792 23570 24848
rect 23626 24792 28000 24848
rect 23565 24790 28000 24792
rect 23565 24787 23631 24790
rect 27520 24760 28000 24790
rect 5533 24714 5599 24717
rect 13997 24714 14063 24717
rect 5533 24712 14063 24714
rect 5533 24656 5538 24712
rect 5594 24656 14002 24712
rect 14058 24656 14063 24712
rect 5533 24654 14063 24656
rect 5533 24651 5599 24654
rect 13997 24651 14063 24654
rect 19517 24714 19583 24717
rect 25405 24714 25471 24717
rect 19517 24712 25471 24714
rect 19517 24656 19522 24712
rect 19578 24656 25410 24712
rect 25466 24656 25471 24712
rect 19517 24654 25471 24656
rect 19517 24651 19583 24654
rect 25405 24651 25471 24654
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24209 24306 24275 24309
rect 27520 24306 28000 24336
rect 24209 24304 28000 24306
rect 24209 24248 24214 24304
rect 24270 24248 28000 24304
rect 24209 24246 28000 24248
rect 24209 24243 24275 24246
rect 27520 24216 28000 24246
rect 4889 24170 4955 24173
rect 12157 24170 12223 24173
rect 4889 24168 12223 24170
rect 4889 24112 4894 24168
rect 4950 24112 12162 24168
rect 12218 24112 12223 24168
rect 4889 24110 12223 24112
rect 4889 24107 4955 24110
rect 12157 24107 12223 24110
rect 20161 24034 20227 24037
rect 24117 24034 24183 24037
rect 20161 24032 24183 24034
rect 20161 23976 20166 24032
rect 20222 23976 24122 24032
rect 24178 23976 24183 24032
rect 20161 23974 24183 23976
rect 20161 23971 20227 23974
rect 24117 23971 24183 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 24669 23898 24735 23901
rect 26233 23898 26299 23901
rect 24669 23896 26299 23898
rect 24669 23840 24674 23896
rect 24730 23840 26238 23896
rect 26294 23840 26299 23896
rect 24669 23838 26299 23840
rect 24669 23835 24735 23838
rect 26233 23835 26299 23838
rect 4245 23762 4311 23765
rect 9949 23762 10015 23765
rect 4245 23760 10015 23762
rect 4245 23704 4250 23760
rect 4306 23704 9954 23760
rect 10010 23704 10015 23760
rect 4245 23702 10015 23704
rect 4245 23699 4311 23702
rect 9949 23699 10015 23702
rect 12985 23762 13051 23765
rect 19149 23762 19215 23765
rect 12985 23760 19215 23762
rect 12985 23704 12990 23760
rect 13046 23704 19154 23760
rect 19210 23704 19215 23760
rect 12985 23702 19215 23704
rect 12985 23699 13051 23702
rect 19149 23699 19215 23702
rect 22461 23762 22527 23765
rect 27520 23762 28000 23792
rect 22461 23760 28000 23762
rect 22461 23704 22466 23760
rect 22522 23704 28000 23760
rect 22461 23702 28000 23704
rect 22461 23699 22527 23702
rect 27520 23672 28000 23702
rect 933 23626 999 23629
rect 18597 23626 18663 23629
rect 933 23624 18663 23626
rect 933 23568 938 23624
rect 994 23568 18602 23624
rect 18658 23568 18663 23624
rect 933 23566 18663 23568
rect 933 23563 999 23566
rect 18597 23563 18663 23566
rect 14089 23490 14155 23493
rect 18505 23490 18571 23493
rect 14089 23488 18571 23490
rect 14089 23432 14094 23488
rect 14150 23432 18510 23488
rect 18566 23432 18571 23488
rect 14089 23430 18571 23432
rect 14089 23427 14155 23430
rect 18505 23427 18571 23430
rect 25221 23490 25287 23493
rect 25221 23488 25330 23490
rect 25221 23432 25226 23488
rect 25282 23432 25330 23488
rect 25221 23427 25330 23432
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 14365 23354 14431 23357
rect 17033 23354 17099 23357
rect 14365 23352 18706 23354
rect 14365 23296 14370 23352
rect 14426 23296 17038 23352
rect 17094 23296 18706 23352
rect 14365 23294 18706 23296
rect 14365 23291 14431 23294
rect 17033 23291 17099 23294
rect 6269 23082 6335 23085
rect 13629 23082 13695 23085
rect 6269 23080 13695 23082
rect 6269 23024 6274 23080
rect 6330 23024 13634 23080
rect 13690 23024 13695 23080
rect 6269 23022 13695 23024
rect 18646 23082 18706 23294
rect 18873 23218 18939 23221
rect 23473 23218 23539 23221
rect 18873 23216 23539 23218
rect 18873 23160 18878 23216
rect 18934 23160 23478 23216
rect 23534 23160 23539 23216
rect 18873 23158 23539 23160
rect 25270 23218 25330 23427
rect 27520 23218 28000 23248
rect 25270 23158 28000 23218
rect 18873 23155 18939 23158
rect 23473 23155 23539 23158
rect 27520 23128 28000 23158
rect 22829 23082 22895 23085
rect 23473 23082 23539 23085
rect 23933 23082 23999 23085
rect 18646 23080 23999 23082
rect 18646 23024 22834 23080
rect 22890 23024 23478 23080
rect 23534 23024 23938 23080
rect 23994 23024 23999 23080
rect 18646 23022 23999 23024
rect 6269 23019 6335 23022
rect 13629 23019 13695 23022
rect 22829 23019 22895 23022
rect 23473 23019 23539 23022
rect 23933 23019 23999 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 13537 22674 13603 22677
rect 21817 22674 21883 22677
rect 13537 22672 21883 22674
rect 13537 22616 13542 22672
rect 13598 22616 21822 22672
rect 21878 22616 21883 22672
rect 13537 22614 21883 22616
rect 13537 22611 13603 22614
rect 21817 22611 21883 22614
rect 1577 22538 1643 22541
rect 16113 22538 16179 22541
rect 1577 22536 16179 22538
rect 1577 22480 1582 22536
rect 1638 22480 16118 22536
rect 16174 22480 16179 22536
rect 1577 22478 16179 22480
rect 1577 22475 1643 22478
rect 16113 22475 16179 22478
rect 17401 22538 17467 22541
rect 22921 22538 22987 22541
rect 17401 22536 22987 22538
rect 17401 22480 17406 22536
rect 17462 22480 22926 22536
rect 22982 22480 22987 22536
rect 17401 22478 22987 22480
rect 17401 22475 17467 22478
rect 22921 22475 22987 22478
rect 25865 22538 25931 22541
rect 27520 22538 28000 22568
rect 25865 22536 28000 22538
rect 25865 22480 25870 22536
rect 25926 22480 28000 22536
rect 25865 22478 28000 22480
rect 25865 22475 25931 22478
rect 27520 22448 28000 22478
rect 23657 22402 23723 22405
rect 23933 22402 23999 22405
rect 23657 22400 23999 22402
rect 23657 22344 23662 22400
rect 23718 22344 23938 22400
rect 23994 22344 23999 22400
rect 23657 22342 23999 22344
rect 23657 22339 23723 22342
rect 23933 22339 23999 22342
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 10869 21994 10935 21997
rect 16757 21994 16823 21997
rect 17401 21994 17467 21997
rect 10869 21992 17467 21994
rect 10869 21936 10874 21992
rect 10930 21936 16762 21992
rect 16818 21936 17406 21992
rect 17462 21936 17467 21992
rect 10869 21934 17467 21936
rect 10869 21931 10935 21934
rect 16757 21931 16823 21934
rect 17401 21931 17467 21934
rect 24025 21994 24091 21997
rect 24393 21994 24459 21997
rect 24025 21992 24459 21994
rect 24025 21936 24030 21992
rect 24086 21936 24398 21992
rect 24454 21936 24459 21992
rect 24025 21934 24459 21936
rect 24025 21931 24091 21934
rect 24393 21931 24459 21934
rect 25037 21994 25103 21997
rect 27520 21994 28000 22024
rect 25037 21992 28000 21994
rect 25037 21936 25042 21992
rect 25098 21936 28000 21992
rect 25037 21934 28000 21936
rect 25037 21931 25103 21934
rect 27520 21904 28000 21934
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 24117 21450 24183 21453
rect 27520 21450 28000 21480
rect 24117 21448 28000 21450
rect 24117 21392 24122 21448
rect 24178 21392 28000 21448
rect 24117 21390 28000 21392
rect 24117 21387 24183 21390
rect 27520 21360 28000 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 16481 21178 16547 21181
rect 18321 21178 18387 21181
rect 16481 21176 18387 21178
rect 16481 21120 16486 21176
rect 16542 21120 18326 21176
rect 18382 21120 18387 21176
rect 16481 21118 18387 21120
rect 16481 21115 16547 21118
rect 18321 21115 18387 21118
rect 13721 21042 13787 21045
rect 15469 21042 15535 21045
rect 13721 21040 15535 21042
rect 13721 20984 13726 21040
rect 13782 20984 15474 21040
rect 15530 20984 15535 21040
rect 13721 20982 15535 20984
rect 13721 20979 13787 20982
rect 15469 20979 15535 20982
rect 23933 20906 23999 20909
rect 27520 20906 28000 20936
rect 23933 20904 28000 20906
rect 23933 20848 23938 20904
rect 23994 20848 28000 20904
rect 23933 20846 28000 20848
rect 23933 20843 23999 20846
rect 27520 20816 28000 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 21357 20634 21423 20637
rect 24117 20634 24183 20637
rect 21357 20632 24183 20634
rect 21357 20576 21362 20632
rect 21418 20576 24122 20632
rect 24178 20576 24183 20632
rect 21357 20574 24183 20576
rect 21357 20571 21423 20574
rect 24117 20571 24183 20574
rect 19057 20498 19123 20501
rect 24025 20498 24091 20501
rect 19057 20496 24091 20498
rect 19057 20440 19062 20496
rect 19118 20440 24030 20496
rect 24086 20440 24091 20496
rect 19057 20438 24091 20440
rect 19057 20435 19123 20438
rect 24025 20435 24091 20438
rect 13721 20362 13787 20365
rect 16573 20362 16639 20365
rect 19425 20362 19491 20365
rect 13721 20360 19491 20362
rect 13721 20304 13726 20360
rect 13782 20304 16578 20360
rect 16634 20304 19430 20360
rect 19486 20304 19491 20360
rect 13721 20302 19491 20304
rect 13721 20299 13787 20302
rect 16573 20299 16639 20302
rect 19425 20299 19491 20302
rect 22369 20362 22435 20365
rect 27520 20362 28000 20392
rect 22369 20360 28000 20362
rect 22369 20304 22374 20360
rect 22430 20304 28000 20360
rect 22369 20302 28000 20304
rect 22369 20299 22435 20302
rect 27520 20272 28000 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 13445 19954 13511 19957
rect 19057 19954 19123 19957
rect 13445 19952 19123 19954
rect 13445 19896 13450 19952
rect 13506 19896 19062 19952
rect 19118 19896 19123 19952
rect 13445 19894 19123 19896
rect 13445 19891 13511 19894
rect 19057 19891 19123 19894
rect 2221 19818 2287 19821
rect 12893 19818 12959 19821
rect 2221 19816 12959 19818
rect 2221 19760 2226 19816
rect 2282 19760 12898 19816
rect 12954 19760 12959 19816
rect 2221 19758 12959 19760
rect 2221 19755 2287 19758
rect 12893 19755 12959 19758
rect 27520 19682 28000 19712
rect 24902 19622 28000 19682
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 23933 19546 23999 19549
rect 15334 19544 23999 19546
rect 15334 19488 23938 19544
rect 23994 19488 23999 19544
rect 15334 19486 23999 19488
rect 8937 19410 9003 19413
rect 15334 19410 15394 19486
rect 23933 19483 23999 19486
rect 8937 19408 15394 19410
rect 8937 19352 8942 19408
rect 8998 19352 15394 19408
rect 8937 19350 15394 19352
rect 21449 19410 21515 19413
rect 24902 19410 24962 19622
rect 27520 19592 28000 19622
rect 21449 19408 24962 19410
rect 21449 19352 21454 19408
rect 21510 19352 24962 19408
rect 21449 19350 24962 19352
rect 8937 19347 9003 19350
rect 21449 19347 21515 19350
rect 6913 19274 6979 19277
rect 17769 19274 17835 19277
rect 6913 19272 17835 19274
rect 6913 19216 6918 19272
rect 6974 19216 17774 19272
rect 17830 19216 17835 19272
rect 6913 19214 17835 19216
rect 6913 19211 6979 19214
rect 17769 19211 17835 19214
rect 19057 19274 19123 19277
rect 23013 19274 23079 19277
rect 19057 19272 23079 19274
rect 19057 19216 19062 19272
rect 19118 19216 23018 19272
rect 23074 19216 23079 19272
rect 19057 19214 23079 19216
rect 19057 19211 19123 19214
rect 23013 19211 23079 19214
rect 23381 19138 23447 19141
rect 27520 19138 28000 19168
rect 23381 19136 28000 19138
rect 23381 19080 23386 19136
rect 23442 19080 28000 19136
rect 23381 19078 28000 19080
rect 23381 19075 23447 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 3601 18866 3667 18869
rect 10133 18866 10199 18869
rect 3601 18864 10199 18866
rect 3601 18808 3606 18864
rect 3662 18808 10138 18864
rect 10194 18808 10199 18864
rect 3601 18806 10199 18808
rect 3601 18803 3667 18806
rect 10133 18803 10199 18806
rect 25497 18866 25563 18869
rect 27521 18866 27587 18869
rect 25497 18864 27587 18866
rect 25497 18808 25502 18864
rect 25558 18808 27526 18864
rect 27582 18808 27587 18864
rect 25497 18806 27587 18808
rect 25497 18803 25563 18806
rect 27521 18803 27587 18806
rect 23565 18730 23631 18733
rect 23565 18728 24824 18730
rect 23565 18672 23570 18728
rect 23626 18672 24824 18728
rect 23565 18670 24824 18672
rect 23565 18667 23631 18670
rect 24764 18594 24824 18670
rect 27520 18594 28000 18624
rect 24764 18534 28000 18594
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 27520 18504 28000 18534
rect 24277 18463 24597 18464
rect 18781 18186 18847 18189
rect 22737 18186 22803 18189
rect 24025 18186 24091 18189
rect 18781 18184 24091 18186
rect 18781 18128 18786 18184
rect 18842 18128 22742 18184
rect 22798 18128 24030 18184
rect 24086 18128 24091 18184
rect 18781 18126 24091 18128
rect 18781 18123 18847 18126
rect 22737 18123 22803 18126
rect 24025 18123 24091 18126
rect 24117 18050 24183 18053
rect 27520 18050 28000 18080
rect 24117 18048 28000 18050
rect 24117 17992 24122 18048
rect 24178 17992 28000 18048
rect 24117 17990 28000 17992
rect 24117 17987 24183 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 27520 17960 28000 17990
rect 19610 17919 19930 17920
rect 7557 17778 7623 17781
rect 21449 17778 21515 17781
rect 7557 17776 21515 17778
rect 7557 17720 7562 17776
rect 7618 17720 21454 17776
rect 21510 17720 21515 17776
rect 7557 17718 21515 17720
rect 7557 17715 7623 17718
rect 21449 17715 21515 17718
rect 24669 17506 24735 17509
rect 27520 17506 28000 17536
rect 24669 17504 28000 17506
rect 24669 17448 24674 17504
rect 24730 17448 28000 17504
rect 24669 17446 28000 17448
rect 24669 17443 24735 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 27520 17416 28000 17446
rect 24277 17375 24597 17376
rect 2865 17234 2931 17237
rect 16113 17234 16179 17237
rect 2865 17232 16179 17234
rect 2865 17176 2870 17232
rect 2926 17176 16118 17232
rect 16174 17176 16179 17232
rect 2865 17174 16179 17176
rect 2865 17171 2931 17174
rect 16113 17171 16179 17174
rect 8201 17098 8267 17101
rect 23197 17098 23263 17101
rect 8201 17096 23263 17098
rect 8201 17040 8206 17096
rect 8262 17040 23202 17096
rect 23258 17040 23263 17096
rect 8201 17038 23263 17040
rect 8201 17035 8267 17038
rect 23197 17035 23263 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 15009 16826 15075 16829
rect 18965 16826 19031 16829
rect 23933 16826 23999 16829
rect 27520 16826 28000 16856
rect 15009 16824 19442 16826
rect 15009 16768 15014 16824
rect 15070 16768 18970 16824
rect 19026 16768 19442 16824
rect 15009 16766 19442 16768
rect 15009 16763 15075 16766
rect 18965 16763 19031 16766
rect 10685 16690 10751 16693
rect 12801 16690 12867 16693
rect 10685 16688 12867 16690
rect 10685 16632 10690 16688
rect 10746 16632 12806 16688
rect 12862 16632 12867 16688
rect 10685 16630 12867 16632
rect 19382 16690 19442 16766
rect 23933 16824 28000 16826
rect 23933 16768 23938 16824
rect 23994 16768 28000 16824
rect 23933 16766 28000 16768
rect 23933 16763 23999 16766
rect 27520 16736 28000 16766
rect 21817 16690 21883 16693
rect 19382 16688 21883 16690
rect 19382 16632 21822 16688
rect 21878 16632 21883 16688
rect 19382 16630 21883 16632
rect 10685 16627 10751 16630
rect 12801 16627 12867 16630
rect 21817 16627 21883 16630
rect 11145 16554 11211 16557
rect 17125 16554 17191 16557
rect 11145 16552 17191 16554
rect 11145 16496 11150 16552
rect 11206 16496 17130 16552
rect 17186 16496 17191 16552
rect 11145 16494 17191 16496
rect 11145 16491 11211 16494
rect 17125 16491 17191 16494
rect 19149 16554 19215 16557
rect 25405 16554 25471 16557
rect 19149 16552 25471 16554
rect 19149 16496 19154 16552
rect 19210 16496 25410 16552
rect 25466 16496 25471 16552
rect 19149 16494 25471 16496
rect 19149 16491 19215 16494
rect 25405 16491 25471 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 25865 16282 25931 16285
rect 27520 16282 28000 16312
rect 25865 16280 28000 16282
rect 25865 16224 25870 16280
rect 25926 16224 28000 16280
rect 25865 16222 28000 16224
rect 25865 16219 25931 16222
rect 27520 16192 28000 16222
rect 3325 16010 3391 16013
rect 10685 16010 10751 16013
rect 3325 16008 10751 16010
rect 3325 15952 3330 16008
rect 3386 15952 10690 16008
rect 10746 15952 10751 16008
rect 3325 15950 10751 15952
rect 3325 15947 3391 15950
rect 10685 15947 10751 15950
rect 17861 16010 17927 16013
rect 25221 16010 25287 16013
rect 17861 16008 25287 16010
rect 17861 15952 17866 16008
rect 17922 15952 25226 16008
rect 25282 15952 25287 16008
rect 17861 15950 25287 15952
rect 17861 15947 17927 15950
rect 25221 15947 25287 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 25037 15738 25103 15741
rect 27520 15738 28000 15768
rect 25037 15736 28000 15738
rect 25037 15680 25042 15736
rect 25098 15680 28000 15736
rect 25037 15678 28000 15680
rect 25037 15675 25103 15678
rect 27520 15648 28000 15678
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 27520 15194 28000 15224
rect 24902 15134 28000 15194
rect 16205 15058 16271 15061
rect 21265 15058 21331 15061
rect 24902 15058 24962 15134
rect 27520 15104 28000 15134
rect 16205 15056 20730 15058
rect 16205 15000 16210 15056
rect 16266 15000 20730 15056
rect 16205 14998 20730 15000
rect 16205 14995 16271 14998
rect 20670 14922 20730 14998
rect 21265 15056 24962 15058
rect 21265 15000 21270 15056
rect 21326 15000 24962 15056
rect 21265 14998 24962 15000
rect 21265 14995 21331 14998
rect 24761 14922 24827 14925
rect 20670 14920 24827 14922
rect 20670 14864 24766 14920
rect 24822 14864 24827 14920
rect 20670 14862 24827 14864
rect 24761 14859 24827 14862
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 24577 14650 24643 14653
rect 27520 14650 28000 14680
rect 24577 14648 28000 14650
rect 24577 14592 24582 14648
rect 24638 14592 28000 14648
rect 24577 14590 28000 14592
rect 24577 14587 24643 14590
rect 27520 14560 28000 14590
rect 19057 14514 19123 14517
rect 20989 14514 21055 14517
rect 19057 14512 21055 14514
rect 19057 14456 19062 14512
rect 19118 14456 20994 14512
rect 21050 14456 21055 14512
rect 19057 14454 21055 14456
rect 19057 14451 19123 14454
rect 20989 14451 21055 14454
rect 5610 14176 5930 14177
rect 0 14106 480 14136
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 3325 14106 3391 14109
rect 0 14104 3391 14106
rect 0 14048 3330 14104
rect 3386 14048 3391 14104
rect 0 14046 3391 14048
rect 0 14016 480 14046
rect 3325 14043 3391 14046
rect 24209 13970 24275 13973
rect 27520 13970 28000 14000
rect 24209 13968 28000 13970
rect 24209 13912 24214 13968
rect 24270 13912 28000 13968
rect 24209 13910 28000 13912
rect 24209 13907 24275 13910
rect 27520 13880 28000 13910
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 14181 13426 14247 13429
rect 21357 13426 21423 13429
rect 14181 13424 21423 13426
rect 14181 13368 14186 13424
rect 14242 13368 21362 13424
rect 21418 13368 21423 13424
rect 14181 13366 21423 13368
rect 14181 13363 14247 13366
rect 21357 13363 21423 13366
rect 24577 13426 24643 13429
rect 27520 13426 28000 13456
rect 24577 13424 28000 13426
rect 24577 13368 24582 13424
rect 24638 13368 28000 13424
rect 24577 13366 28000 13368
rect 24577 13363 24643 13366
rect 27520 13336 28000 13366
rect 14365 13290 14431 13293
rect 24761 13290 24827 13293
rect 14365 13288 24827 13290
rect 14365 13232 14370 13288
rect 14426 13232 24766 13288
rect 24822 13232 24827 13288
rect 14365 13230 24827 13232
rect 14365 13227 14431 13230
rect 24761 13227 24827 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 16941 12882 17007 12885
rect 21173 12882 21239 12885
rect 16941 12880 21239 12882
rect 16941 12824 16946 12880
rect 17002 12824 21178 12880
rect 21234 12824 21239 12880
rect 16941 12822 21239 12824
rect 16941 12819 17007 12822
rect 21173 12819 21239 12822
rect 21357 12882 21423 12885
rect 27520 12882 28000 12912
rect 21357 12880 28000 12882
rect 21357 12824 21362 12880
rect 21418 12824 28000 12880
rect 21357 12822 28000 12824
rect 21357 12819 21423 12822
rect 27520 12792 28000 12822
rect 381 12746 447 12749
rect 13997 12746 14063 12749
rect 381 12744 14063 12746
rect 381 12688 386 12744
rect 442 12688 14002 12744
rect 14058 12688 14063 12744
rect 381 12686 14063 12688
rect 381 12683 447 12686
rect 13997 12683 14063 12686
rect 16849 12746 16915 12749
rect 24209 12746 24275 12749
rect 16849 12744 24275 12746
rect 16849 12688 16854 12744
rect 16910 12688 24214 12744
rect 24270 12688 24275 12744
rect 16849 12686 24275 12688
rect 16849 12683 16915 12686
rect 24209 12683 24275 12686
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 27520 12338 28000 12368
rect 26374 12278 28000 12338
rect 24577 12202 24643 12205
rect 26374 12202 26434 12278
rect 27520 12248 28000 12278
rect 24577 12200 26434 12202
rect 24577 12144 24582 12200
rect 24638 12144 26434 12200
rect 24577 12142 26434 12144
rect 24577 12139 24643 12142
rect 5610 12000 5930 12001
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 27520 11794 28000 11824
rect 27478 11704 28000 11794
rect 12893 11658 12959 11661
rect 27478 11658 27538 11704
rect 12893 11656 27538 11658
rect 12893 11600 12898 11656
rect 12954 11600 27538 11656
rect 12893 11598 27538 11600
rect 12893 11595 12959 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 12249 11114 12315 11117
rect 27520 11114 28000 11144
rect 12249 11112 28000 11114
rect 12249 11056 12254 11112
rect 12310 11056 28000 11112
rect 12249 11054 28000 11056
rect 12249 11051 12315 11054
rect 27520 11024 28000 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 11421 10570 11487 10573
rect 27520 10570 28000 10600
rect 11421 10568 28000 10570
rect 11421 10512 11426 10568
rect 11482 10512 28000 10568
rect 11421 10510 28000 10512
rect 11421 10507 11487 10510
rect 27520 10480 28000 10510
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 10869 10026 10935 10029
rect 27520 10026 28000 10056
rect 10869 10024 28000 10026
rect 10869 9968 10874 10024
rect 10930 9968 28000 10024
rect 10869 9966 28000 9968
rect 10869 9963 10935 9966
rect 27520 9936 28000 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 10225 9482 10291 9485
rect 27520 9482 28000 9512
rect 10225 9480 28000 9482
rect 10225 9424 10230 9480
rect 10286 9424 28000 9480
rect 10225 9422 28000 9424
rect 10225 9419 10291 9422
rect 27520 9392 28000 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 9857 8938 9923 8941
rect 27520 8938 28000 8968
rect 9857 8936 28000 8938
rect 9857 8880 9862 8936
rect 9918 8880 28000 8936
rect 9857 8878 28000 8880
rect 9857 8875 9923 8878
rect 27520 8848 28000 8878
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 18137 8394 18203 8397
rect 19333 8394 19399 8397
rect 18137 8392 19399 8394
rect 18137 8336 18142 8392
rect 18198 8336 19338 8392
rect 19394 8336 19399 8392
rect 18137 8334 19399 8336
rect 18137 8331 18203 8334
rect 19333 8331 19399 8334
rect 13353 8258 13419 8261
rect 13997 8258 14063 8261
rect 13353 8256 14063 8258
rect 13353 8200 13358 8256
rect 13414 8200 14002 8256
rect 14058 8200 14063 8256
rect 13353 8198 14063 8200
rect 13353 8195 13419 8198
rect 13997 8195 14063 8198
rect 24761 8258 24827 8261
rect 27520 8258 28000 8288
rect 24761 8256 28000 8258
rect 24761 8200 24766 8256
rect 24822 8200 28000 8256
rect 24761 8198 28000 8200
rect 24761 8195 24827 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 25313 7714 25379 7717
rect 27520 7714 28000 7744
rect 25313 7712 28000 7714
rect 25313 7656 25318 7712
rect 25374 7656 28000 7712
rect 25313 7654 28000 7656
rect 25313 7651 25379 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 19609 7442 19675 7445
rect 24577 7442 24643 7445
rect 19609 7440 24643 7442
rect 19609 7384 19614 7440
rect 19670 7384 24582 7440
rect 24638 7384 24643 7440
rect 19609 7382 24643 7384
rect 19609 7379 19675 7382
rect 24577 7379 24643 7382
rect 24761 7170 24827 7173
rect 27520 7170 28000 7200
rect 24761 7168 28000 7170
rect 24761 7112 24766 7168
rect 24822 7112 28000 7168
rect 24761 7110 28000 7112
rect 24761 7107 24827 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 27520 7080 28000 7110
rect 19610 7039 19930 7040
rect 24669 6626 24735 6629
rect 27520 6626 28000 6656
rect 24669 6624 28000 6626
rect 24669 6568 24674 6624
rect 24730 6568 28000 6624
rect 24669 6566 28000 6568
rect 24669 6563 24735 6566
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 27520 6536 28000 6566
rect 24277 6495 24597 6496
rect 15377 6490 15443 6493
rect 23473 6490 23539 6493
rect 15377 6488 23539 6490
rect 15377 6432 15382 6488
rect 15438 6432 23478 6488
rect 23534 6432 23539 6488
rect 15377 6430 23539 6432
rect 15377 6427 15443 6430
rect 23473 6427 23539 6430
rect 9949 6354 10015 6357
rect 23657 6354 23723 6357
rect 9949 6352 23723 6354
rect 9949 6296 9954 6352
rect 10010 6296 23662 6352
rect 23718 6296 23723 6352
rect 9949 6294 23723 6296
rect 9949 6291 10015 6294
rect 23657 6291 23723 6294
rect 15193 6218 15259 6221
rect 24945 6218 25011 6221
rect 15193 6216 25011 6218
rect 15193 6160 15198 6216
rect 15254 6160 24950 6216
rect 25006 6160 25011 6216
rect 15193 6158 25011 6160
rect 15193 6155 15259 6158
rect 24945 6155 25011 6158
rect 25129 6082 25195 6085
rect 27520 6082 28000 6112
rect 25129 6080 28000 6082
rect 25129 6024 25134 6080
rect 25190 6024 28000 6080
rect 25129 6022 28000 6024
rect 25129 6019 25195 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 10041 5810 10107 5813
rect 23657 5810 23723 5813
rect 10041 5808 23723 5810
rect 10041 5752 10046 5808
rect 10102 5752 23662 5808
rect 23718 5752 23723 5808
rect 10041 5750 23723 5752
rect 10041 5747 10107 5750
rect 23657 5747 23723 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 25129 5402 25195 5405
rect 27520 5402 28000 5432
rect 25129 5400 28000 5402
rect 25129 5344 25134 5400
rect 25190 5344 28000 5400
rect 25129 5342 28000 5344
rect 25129 5339 25195 5342
rect 27520 5312 28000 5342
rect 10777 5130 10843 5133
rect 23657 5130 23723 5133
rect 10777 5128 23723 5130
rect 10777 5072 10782 5128
rect 10838 5072 23662 5128
rect 23718 5072 23723 5128
rect 10777 5070 23723 5072
rect 10777 5067 10843 5070
rect 23657 5067 23723 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 26141 4858 26207 4861
rect 27520 4858 28000 4888
rect 26141 4856 28000 4858
rect 26141 4800 26146 4856
rect 26202 4800 28000 4856
rect 26141 4798 28000 4800
rect 26141 4795 26207 4798
rect 27520 4768 28000 4798
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 24669 4314 24735 4317
rect 27520 4314 28000 4344
rect 24669 4312 28000 4314
rect 24669 4256 24674 4312
rect 24730 4256 28000 4312
rect 24669 4254 28000 4256
rect 24669 4251 24735 4254
rect 27520 4224 28000 4254
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 25129 3770 25195 3773
rect 27520 3770 28000 3800
rect 25129 3768 28000 3770
rect 25129 3712 25134 3768
rect 25190 3712 28000 3768
rect 25129 3710 28000 3712
rect 25129 3707 25195 3710
rect 27520 3680 28000 3710
rect 19241 3498 19307 3501
rect 24945 3498 25011 3501
rect 19241 3496 25011 3498
rect 19241 3440 19246 3496
rect 19302 3440 24950 3496
rect 25006 3440 25011 3496
rect 19241 3438 25011 3440
rect 19241 3435 19307 3438
rect 24945 3435 25011 3438
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 24669 3226 24735 3229
rect 27520 3226 28000 3256
rect 24669 3224 28000 3226
rect 24669 3168 24674 3224
rect 24730 3168 28000 3224
rect 24669 3166 28000 3168
rect 24669 3163 24735 3166
rect 27520 3136 28000 3166
rect 16113 3090 16179 3093
rect 23473 3090 23539 3093
rect 16113 3088 23539 3090
rect 16113 3032 16118 3088
rect 16174 3032 23478 3088
rect 23534 3032 23539 3088
rect 16113 3030 23539 3032
rect 16113 3027 16179 3030
rect 23473 3027 23539 3030
rect 13445 2954 13511 2957
rect 23657 2954 23723 2957
rect 13445 2952 23723 2954
rect 13445 2896 13450 2952
rect 13506 2896 23662 2952
rect 23718 2896 23723 2952
rect 13445 2894 23723 2896
rect 13445 2891 13511 2894
rect 23657 2891 23723 2894
rect 22553 2818 22619 2821
rect 25313 2818 25379 2821
rect 22553 2816 25379 2818
rect 22553 2760 22558 2816
rect 22614 2760 25318 2816
rect 25374 2760 25379 2816
rect 22553 2758 25379 2760
rect 22553 2755 22619 2758
rect 25313 2755 25379 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 24209 2546 24275 2549
rect 27520 2546 28000 2576
rect 24209 2544 28000 2546
rect 24209 2488 24214 2544
rect 24270 2488 28000 2544
rect 24209 2486 28000 2488
rect 24209 2483 24275 2486
rect 27520 2456 28000 2486
rect 16021 2410 16087 2413
rect 24025 2410 24091 2413
rect 16021 2408 24091 2410
rect 16021 2352 16026 2408
rect 16082 2352 24030 2408
rect 24086 2352 24091 2408
rect 16021 2350 24091 2352
rect 16021 2347 16087 2350
rect 24025 2347 24091 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 23013 2002 23079 2005
rect 27520 2002 28000 2032
rect 23013 2000 28000 2002
rect 23013 1944 23018 2000
rect 23074 1944 28000 2000
rect 23013 1942 28000 1944
rect 23013 1939 23079 1942
rect 27520 1912 28000 1942
rect 24761 1458 24827 1461
rect 27520 1458 28000 1488
rect 24761 1456 28000 1458
rect 24761 1400 24766 1456
rect 24822 1400 28000 1456
rect 24761 1398 28000 1400
rect 24761 1395 24827 1398
rect 27520 1368 28000 1398
rect 25497 914 25563 917
rect 27520 914 28000 944
rect 25497 912 28000 914
rect 25497 856 25502 912
rect 25558 856 28000 912
rect 25497 854 28000 856
rect 25497 851 25563 854
rect 27520 824 28000 854
rect 24117 370 24183 373
rect 27520 370 28000 400
rect 24117 368 28000 370
rect 24117 312 24122 368
rect 24178 312 28000 368
rect 24117 310 28000 312
rect 24117 307 24183 310
rect 27520 280 28000 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
use scs8hd_decap_3  PHY_0 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_15
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_3
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_15
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_27 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_27
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_56 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_59 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_74
timestamp 1586364061
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_87
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_106
timestamp 1586364061
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_118
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_137
timestamp 1586364061
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _53_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_4  mux_right_track_0.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.scs8hd_buf_4_0__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_8  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_228
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_6.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use scs8hd_buf_4  mux_right_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_265
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_4  mux_right_track_2.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 590 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_decap_6  FILLER_0_271
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_68
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_129
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_141
timestamp 1586364061
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_202
timestamp 1586364061
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _54_
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_right_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23460 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_4  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_261
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_15
timestamp 1586364061
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_27
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_39
timestamp 1586364061
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_3_59
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_74
timestamp 1586364061
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_98
timestamp 1586364061
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_110
timestamp 1586364061
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_123
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_135
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_147
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_159
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_171
timestamp 1586364061
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_208
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_220
timestamp 1586364061
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_232
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_259
timestamp 1586364061
transform 1 0 24932 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_263
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_275
timestamp 1586364061
transform 1 0 26404 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_56
timestamp 1586364061
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_68
timestamp 1586364061
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_80
timestamp 1586364061
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_105
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_117
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_129
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_190
timestamp 1586364061
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_202
timestamp 1586364061
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_227
timestamp 1586364061
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_239
timestamp 1586364061
transform 1 0 23092 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_8  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_271
timestamp 1586364061
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_51
timestamp 1586364061
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_59
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_74
timestamp 1586364061
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_86
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_98
timestamp 1586364061
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_110
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_135
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_147
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_159
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_184
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_196
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 774 592
use scs8hd_buf_4  mux_right_track_10.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__47__A
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_251
timestamp 1586364061
transform 1 0 24196 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_255
timestamp 1586364061
transform 1 0 24564 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 24932 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 25484 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_263
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_267
timestamp 1586364061
transform 1 0 25668 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_12  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_27
timestamp 1586364061
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_44
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_56
timestamp 1586364061
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_51
timestamp 1586364061
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_59
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_74
timestamp 1586364061
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_80
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_86
timestamp 1586364061
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_98
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_105
timestamp 1586364061
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_117
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_129
timestamp 1586364061
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_135
timestamp 1586364061
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_16.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_166
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_178
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_172
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_190
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_7_180
timestamp 1586364061
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_196
timestamp 1586364061
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_208
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_232
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_buf_4  mux_right_track_14.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 590 592
use scs8hd_buf_4  mux_right_track_12.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_255
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_251
timestamp 1586364061
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24380 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__46__A
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_267
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_263
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 406 592
use scs8hd_buf_2  _47_
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_275
timestamp 1586364061
transform 1 0 26404 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_15
timestamp 1586364061
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_68
timestamp 1586364061
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_80
timestamp 1586364061
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_105
timestamp 1586364061
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_117
timestamp 1586364061
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_166
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_18.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_6  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 590 592
use scs8hd_decap_8  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_2  _46_
timestamp 1586364061
transform 1 0 24932 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_15
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_39
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_59
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_74
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_86
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_110
timestamp 1586364061
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_135
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_147
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_200
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_212
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22908 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_224
timestamp 1586364061
transform 1 0 21712 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 130 592
use scs8hd_buf_2  _45_
timestamp 1586364061
transform 1 0 24564 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__44__A
timestamp 1586364061
transform 1 0 24288 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_239
timestamp 1586364061
transform 1 0 23092 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_243
timestamp 1586364061
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_251
timestamp 1586364061
transform 1 0 24196 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 130 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__45__A
timestamp 1586364061
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_259
timestamp 1586364061
transform 1 0 24932 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_263
timestamp 1586364061
transform 1 0 25300 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_275
timestamp 1586364061
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_15
timestamp 1586364061
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_44
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_56
timestamp 1586364061
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_68
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_80
timestamp 1586364061
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_178
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_20.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19320 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_212
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_22.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22908 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_235
timestamp 1586364061
transform 1 0 22724 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _44_
timestamp 1586364061
transform 1 0 24288 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_243
timestamp 1586364061
transform 1 0 23460 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_256
timestamp 1586364061
transform 1 0 24656 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_268
timestamp 1586364061
transform 1 0 25760 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_274
timestamp 1586364061
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_27
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_39
timestamp 1586364061
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_51
timestamp 1586364061
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__41__A
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_86
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_107
timestamp 1586364061
transform 1 0 10948 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_11_119
timestamp 1586364061
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23828 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_253
timestamp 1586364061
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _43_
timestamp 1586364061
transform 1 0 25116 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__43__A
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_265
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_15
timestamp 1586364061
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_68
timestamp 1586364061
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _41_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_80
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_97
timestamp 1586364061
transform 1 0 10028 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_109
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_121
timestamp 1586364061
transform 1 0 12236 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_4  mux_right_track_26.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24288 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_12_270
timestamp 1586364061
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_274
timestamp 1586364061
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _40_
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _39_
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__40__A
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__39__A
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_105
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_14_101
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_121
timestamp 1586364061
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_120
timestamp 1586364061
transform 1 0 12144 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_132
timestamp 1586364061
transform 1 0 13248 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_144
timestamp 1586364061
transform 1 0 14352 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_152
timestamp 1586364061
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _42_
timestamp 1586364061
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_253
timestamp 1586364061
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__42__A
timestamp 1586364061
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_259
timestamp 1586364061
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_263
timestamp 1586364061
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_13_275
timestamp 1586364061
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_buf_2  _38_
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__38__A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__37__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _37_
timestamp 1586364061
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_123
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_147
timestamp 1586364061
transform 1 0 14628 0 -1 11424
box -38 -48 590 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_buf_2  _36_
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__36__A
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_134
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_146
timestamp 1586364061
transform 1 0 14536 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_170
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_253
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_132
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_138
timestamp 1586364061
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_142
timestamp 1586364061
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16836 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_173
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_185
timestamp 1586364061
transform 1 0 18124 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_209
timestamp 1586364061
transform 1 0 20332 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 24564 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_259
timestamp 1586364061
transform 1 0 24932 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_271
timestamp 1586364061
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_68
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_19_127
timestamp 1586364061
transform 1 0 12788 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12880 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_20_130
timestamp 1586364061
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_mux2_2  mux_top_track_0.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13064 0 1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_157
timestamp 1586364061
transform 1 0 15548 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16836 0 -1 13600
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_162
timestamp 1586364061
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_20_198
timestamp 1586364061
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_219
timestamp 1586364061
transform 1 0 21252 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_231
timestamp 1586364061
transform 1 0 22356 0 -1 13600
box -38 -48 1142 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 24564 0 -1 13600
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 24564 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_253
timestamp 1586364061
transform 1 0 24380 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_243
timestamp 1586364061
transform 1 0 23460 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_259
timestamp 1586364061
transform 1 0 24932 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_271
timestamp 1586364061
transform 1 0 26036 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_21_3
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_27
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_39
timestamp 1586364061
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12696 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_top_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_174
timestamp 1586364061
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_178
timestamp 1586364061
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_182
timestamp 1586364061
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17664 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_3  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_189
timestamp 1586364061
transform 1 0 18492 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19504 0 1 13600
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_223
timestamp 1586364061
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_227
timestamp 1586364061
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 24564 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_239
timestamp 1586364061
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_243
timestamp 1586364061
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_21_253
timestamp 1586364061
transform 1 0 24380 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_15
timestamp 1586364061
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 774 592
use scs8hd_conb_1  _19_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_128
timestamp 1586364061
transform 1 0 12880 0 -1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_145
timestamp 1586364061
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_8  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use scs8hd_mux2_2  mux_top_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_162
timestamp 1586364061
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_175
timestamp 1586364061
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_top_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 1786 592
use scs8hd_mux2_2  mux_top_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_206
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_12  FILLER_22_224
timestamp 1586364061
transform 1 0 21712 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_236
timestamp 1586364061
transform 1 0 22816 0 -1 14688
box -38 -48 1142 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_6  FILLER_22_248
timestamp 1586364061
transform 1 0 23920 0 -1 14688
box -38 -48 590 592
use scs8hd_fill_1  FILLER_22_254
timestamp 1586364061
transform 1 0 24472 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_259
timestamp 1586364061
transform 1 0 24932 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_271
timestamp 1586364061
transform 1 0 26036 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_0.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 12880 0 1 14688
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_127
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_134
timestamp 1586364061
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 1142 592
use scs8hd_buf_4  mux_top_track_4.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15548 0 1 14688
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_4.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_150
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_154
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 130 592
use scs8hd_conb_1  _21_
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_163
timestamp 1586364061
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_167
timestamp 1586364061
transform 1 0 16468 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_174
timestamp 1586364061
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use scs8hd_mux2_2  mux_top_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_decap_6  FILLER_23_198
timestamp 1586364061
transform 1 0 19320 0 1 14688
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 20056 0 1 14688
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22540 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_225
timestamp 1586364061
transform 1 0 21804 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_235
timestamp 1586364061
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_239
timestamp 1586364061
transform 1 0 23092 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_243
timestamp 1586364061
transform 1 0 23460 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_23_262
timestamp 1586364061
transform 1 0 25208 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_23_274
timestamp 1586364061
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_6  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_144
timestamp 1586364061
transform 1 0 14352 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_24_152
timestamp 1586364061
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_8.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 866 592
use scs8hd_fill_2  FILLER_24_162
timestamp 1586364061
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_173
timestamp 1586364061
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use scs8hd_conb_1  _22_
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 314 592
use scs8hd_buf_4  mux_top_track_8.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 17756 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_8  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_208
timestamp 1586364061
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22540 0 -1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_219
timestamp 1586364061
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_223
timestamp 1586364061
transform 1 0 21620 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_252
timestamp 1586364061
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_256
timestamp 1586364061
transform 1 0 24656 0 -1 15776
box -38 -48 406 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 25024 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_264
timestamp 1586364061
transform 1 0 25392 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_272
timestamp 1586364061
transform 1 0 26128 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_108
timestamp 1586364061
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_112
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_120
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use scs8hd_fill_2  FILLER_25_131
timestamp 1586364061
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_139
timestamp 1586364061
transform 1 0 13892 0 1 15776
box -38 -48 130 592
use scs8hd_conb_1  _18_
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_8.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_161
timestamp 1586364061
transform 1 0 15916 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_165
timestamp 1586364061
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_169
timestamp 1586364061
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_174
timestamp 1586364061
transform 1 0 17112 0 1 15776
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18584 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 18952 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_188
timestamp 1586364061
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_192
timestamp 1586364061
transform 1 0 18768 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_218
timestamp 1586364061
transform 1 0 21160 0 1 15776
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_22.mux_l2_in_0_
timestamp 1586364061
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_230
timestamp 1586364061
transform 1 0 22264 0 1 15776
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_240
timestamp 1586364061
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_254
timestamp 1586364061
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_258
timestamp 1586364061
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_266
timestamp 1586364061
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_270
timestamp 1586364061
transform 1 0 25944 0 1 15776
box -38 -48 590 592
use scs8hd_fill_1  FILLER_25_276
timestamp 1586364061
transform 1 0 26496 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10856 0 -1 16864
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_6.mux_l3_in_0_
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 13156 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_125
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 590 592
use scs8hd_decap_4  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_142
timestamp 1586364061
transform 1 0 14168 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_4  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_158
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_148
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_152
timestamp 1586364061
transform 1 0 15088 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_158
timestamp 1586364061
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_right_track_8.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_161
timestamp 1586364061
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_174
timestamp 1586364061
transform 1 0 17112 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_8.mux_l1_in_1_
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_20.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_197
timestamp 1586364061
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_195
timestamp 1586364061
transform 1 0 19044 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_22.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20976 0 -1 16864
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_22.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_203
timestamp 1586364061
transform 1 0 19780 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_211
timestamp 1586364061
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21528 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_224
timestamp 1586364061
transform 1 0 21712 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21896 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 406 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 22080 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_27_235
timestamp 1586364061
transform 1 0 22724 0 1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_235
timestamp 1586364061
transform 1 0 22724 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_238
timestamp 1586364061
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_242
timestamp 1586364061
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_242
timestamp 1586364061
transform 1 0 23368 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23736 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_1_
timestamp 1586364061
transform 1 0 23736 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_255
timestamp 1586364061
transform 1 0 24564 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23920 0 -1 16864
box -38 -48 1786 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_267
timestamp 1586364061
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_27_259
timestamp 1586364061
transform 1 0 24932 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_27_271
timestamp 1586364061
transform 1 0 26036 0 1 16864
box -38 -48 590 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_112
timestamp 1586364061
transform 1 0 11408 0 -1 17952
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_6.mux_l2_in_1_
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_124
timestamp 1586364061
transform 1 0 12512 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_143
timestamp 1586364061
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_151
timestamp 1586364061
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_158
timestamp 1586364061
transform 1 0 15640 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_164
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_167
timestamp 1586364061
transform 1 0 16468 0 -1 17952
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 18308 0 -1 17952
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_179
timestamp 1586364061
transform 1 0 17572 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_183
timestamp 1586364061
transform 1 0 17940 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_22.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_206
timestamp 1586364061
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_224
timestamp 1586364061
transform 1 0 21712 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_28_236
timestamp 1586364061
transform 1 0 22816 0 -1 17952
box -38 -48 406 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 24748 0 -1 17952
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 23184 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 24564 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_249
timestamp 1586364061
transform 1 0 24012 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_253
timestamp 1586364061
transform 1 0 24380 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_260
timestamp 1586364061
transform 1 0 25024 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_28_272
timestamp 1586364061
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_96
timestamp 1586364061
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_10.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_10.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_100
timestamp 1586364061
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_113
timestamp 1586364061
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_117
timestamp 1586364061
transform 1 0 11868 0 1 17952
box -38 -48 406 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_121
timestamp 1586364061
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_29_129
timestamp 1586364061
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_133
timestamp 1586364061
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_138
timestamp 1586364061
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_18.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_142
timestamp 1586364061
transform 1 0 14168 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_150
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_20.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 590 592
use scs8hd_fill_2  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_175
timestamp 1586364061
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 18676 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_6  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use scs8hd_fill_1  FILLER_29_190
timestamp 1586364061
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_194
timestamp 1586364061
transform 1 0 18952 0 1 17952
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_206
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_29_214
timestamp 1586364061
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_217
timestamp 1586364061
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_221
timestamp 1586364061
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_225
timestamp 1586364061
transform 1 0 21804 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_29_237
timestamp 1586364061
transform 1 0 22908 0 1 17952
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_26.mux_l2_in_0_
timestamp 1586364061
transform 1 0 24380 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 24196 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_29_241
timestamp 1586364061
transform 1 0 23276 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_249
timestamp 1586364061
transform 1 0 24012 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_262
timestamp 1586364061
transform 1 0 25208 0 1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_29_266
timestamp 1586364061
transform 1 0 25576 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_29_274
timestamp 1586364061
transform 1 0 26312 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_10.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_103
timestamp 1586364061
transform 1 0 10580 0 -1 19040
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_6.mux_l2_in_0_
timestamp 1586364061
transform 1 0 13156 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_123
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_127
timestamp 1586364061
transform 1 0 12788 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_130
timestamp 1586364061
transform 1 0 13064 0 -1 19040
box -38 -48 130 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_140
timestamp 1586364061
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_152
timestamp 1586364061
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_158
timestamp 1586364061
transform 1 0 15640 0 -1 19040
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_20.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16652 0 -1 19040
box -38 -48 1786 592
use scs8hd_decap_3  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_192
timestamp 1586364061
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use scs8hd_mux2_2  mux_top_track_24.mux_l1_in_0_
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_204
timestamp 1586364061
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_224
timestamp 1586364061
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_228
timestamp 1586364061
transform 1 0 22080 0 -1 19040
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 23736 0 -1 19040
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_30_240
timestamp 1586364061
transform 1 0 23184 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_265
timestamp 1586364061
transform 1 0 25484 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_273
timestamp 1586364061
transform 1 0 26220 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_94
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_97
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_10.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_101
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_114
timestamp 1586364061
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_118
timestamp 1586364061
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 13156 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_31_127
timestamp 1586364061
transform 1 0 12788 0 1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_31_130
timestamp 1586364061
transform 1 0 13064 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_150
timestamp 1586364061
transform 1 0 14904 0 1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_160
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_164
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 774 592
use scs8hd_fill_1  FILLER_31_172
timestamp 1586364061
transform 1 0 16928 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_20.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_193
timestamp 1586364061
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_197
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_top_track_24.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 20700 0 1 19040
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_24.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 20148 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_201
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 590 592
use scs8hd_fill_2  FILLER_31_209
timestamp 1586364061
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 22632 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_236
timestamp 1586364061
transform 1 0 22816 0 1 19040
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_right_track_26.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 24104 0 1 19040
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 23920 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_32_120
timestamp 1586364061
transform 1 0 12144 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_2  FILLER_32_137
timestamp 1586364061
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 14260 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_173
timestamp 1586364061
transform 1 0 17020 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_177
timestamp 1586364061
transform 1 0 17388 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_2_
timestamp 1586364061
transform 1 0 17756 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_180
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_194
timestamp 1586364061
transform 1 0 18952 0 -1 20128
box -38 -48 774 592
use scs8hd_conb_1  _20_
timestamp 1586364061
transform 1 0 19780 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_210
timestamp 1586364061
transform 1 0 20424 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_213
timestamp 1586364061
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 21712 0 -1 20128
box -38 -48 1786 592
use scs8hd_fill_1  FILLER_32_223
timestamp 1586364061
transform 1 0 21620 0 -1 20128
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_26.mux_l1_in_0_
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 24012 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_26.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23644 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_243
timestamp 1586364061
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_247
timestamp 1586364061
transform 1 0 23828 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_260
timestamp 1586364061
transform 1 0 25024 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_32_272
timestamp 1586364061
transform 1 0 26128 0 -1 20128
box -38 -48 314 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_12.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_12.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_103
timestamp 1586364061
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_107
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use scs8hd_decap_8  FILLER_34_120
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_1  FILLER_33_127
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_130
timestamp 1586364061
transform 1 0 13064 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13248 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_6.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_6.mux_l1_in_1_
timestamp 1586364061
transform 1 0 13432 0 -1 21216
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_6.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13432 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_153
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_158
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_143
timestamp 1586364061
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_147
timestamp 1586364061
transform 1 0 14628 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_4  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_158
timestamp 1586364061
transform 1 0 15640 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_162
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_4.mux_l3_in_0_
timestamp 1586364061
transform 1 0 15916 0 -1 21216
box -38 -48 866 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_1_
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use scs8hd_decap_4  FILLER_34_174
timestamp 1586364061
transform 1 0 17112 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_34_170
timestamp 1586364061
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 16928 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_197
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_201
timestamp 1586364061
transform 1 0 19596 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_6  FILLER_33_203
timestamp 1586364061
transform 1 0 19780 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 19412 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_213
timestamp 1586364061
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_209
timestamp 1586364061
transform 1 0 20332 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_buf_4  mux_top_track_24.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use scs8hd_mux2_2  mux_top_track_24.mux_l2_in_0_
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 866 592
use scs8hd_fill_2  FILLER_34_225
timestamp 1586364061
transform 1 0 21804 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_221
timestamp 1586364061
transform 1 0 21436 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_224
timestamp 1586364061
transform 1 0 21712 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_24.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21528 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_233
timestamp 1586364061
transform 1 0 22540 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_229
timestamp 1586364061
transform 1 0 22172 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_236
timestamp 1586364061
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 22356 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_2_
timestamp 1586364061
transform 1 0 22632 0 -1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_34_243
timestamp 1586364061
transform 1 0 23460 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_240
timestamp 1586364061
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_34_250
timestamp 1586364061
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_247
timestamp 1586364061
transform 1 0 23828 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 24196 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 23920 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_254
timestamp 1586364061
transform 1 0 24472 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_253
timestamp 1586364061
transform 1 0 24380 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 24564 0 -1 21216
box -38 -48 406 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 24472 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 24932 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_261
timestamp 1586364061
transform 1 0 25116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_273
timestamp 1586364061
transform 1 0 26220 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_259
timestamp 1586364061
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_271
timestamp 1586364061
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_92
timestamp 1586364061
transform 1 0 9568 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_96
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_12.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10304 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12052 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_109
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_113
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_117
timestamp 1586364061
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 406 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_127
timestamp 1586364061
transform 1 0 12788 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_130
timestamp 1586364061
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_138
timestamp 1586364061
transform 1 0 13800 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_134
timestamp 1586364061
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_18.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 14352 0 1 21216
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_right_track_18.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 16652 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 17020 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_163
timestamp 1586364061
transform 1 0 16100 0 1 21216
box -38 -48 590 592
use scs8hd_fill_2  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_175
timestamp 1586364061
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use scs8hd_conb_1  _34_
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use scs8hd_mux2_2  mux_right_track_2.mux_l3_in_0_
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 18952 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18492 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_179
timestamp 1586364061
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_191
timestamp 1586364061
transform 1 0 18676 0 1 21216
box -38 -48 314 592
use scs8hd_conb_1  _23_
timestamp 1586364061
transform 1 0 20976 0 1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_205
timestamp 1586364061
transform 1 0 19964 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_209
timestamp 1586364061
transform 1 0 20332 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_215
timestamp 1586364061
transform 1 0 20884 0 1 21216
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_1_
timestamp 1586364061
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_219
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_223
timestamp 1586364061
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_236
timestamp 1586364061
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_0.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_240
timestamp 1586364061
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_264
timestamp 1586364061
transform 1 0 25392 0 1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_35_276
timestamp 1586364061
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_12.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_110
timestamp 1586364061
transform 1 0 11224 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_18.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13616 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_12  FILLER_36_122
timestamp 1586364061
transform 1 0 12328 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_36_134
timestamp 1586364061
transform 1 0 13432 0 -1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_145
timestamp 1586364061
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_149
timestamp 1586364061
transform 1 0 14812 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_1_
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_168
timestamp 1586364061
transform 1 0 16560 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 590 592
use scs8hd_mux2_2  mux_right_track_4.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18216 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 19228 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_195
timestamp 1586364061
transform 1 0 19044 0 -1 22304
box -38 -48 222 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 19780 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 19596 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 21068 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_199
timestamp 1586364061
transform 1 0 19412 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_206
timestamp 1586364061
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l2_in_0_
timestamp 1586364061
transform 1 0 22356 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 21620 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_219
timestamp 1586364061
transform 1 0 21252 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_36_225
timestamp 1586364061
transform 1 0 21804 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_229
timestamp 1586364061
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_0.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 23920 0 -1 22304
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_240
timestamp 1586364061
transform 1 0 23184 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_244
timestamp 1586364061
transform 1 0 23552 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_247
timestamp 1586364061
transform 1 0 23828 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_8  FILLER_36_267
timestamp 1586364061
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 130 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 10488 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10948 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_101
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_105
timestamp 1586364061
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_109
timestamp 1586364061
transform 1 0 11132 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_121
timestamp 1586364061
transform 1 0 12236 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_fill_2  FILLER_37_128
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_132
timestamp 1586364061
transform 1 0 13248 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_138
timestamp 1586364061
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_16.mux_l2_in_0_
timestamp 1586364061
transform 1 0 14168 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_37_151
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_4.mux_l1_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_4.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15824 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_162
timestamp 1586364061
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_175
timestamp 1586364061
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 19320 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 18584 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_179
timestamp 1586364061
transform 1 0 17572 0 1 22304
box -38 -48 406 592
use scs8hd_decap_6  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 590 592
use scs8hd_fill_2  FILLER_37_192
timestamp 1586364061
transform 1 0 18768 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 1786 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_0_
timestamp 1586364061
transform 1 0 21988 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 21804 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_219
timestamp 1586364061
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_223
timestamp 1586364061
transform 1 0 21620 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_236
timestamp 1586364061
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_0.mux_l3_in_0_
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_240
timestamp 1586364061
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_254
timestamp 1586364061
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_258
timestamp 1586364061
transform 1 0 24840 0 1 22304
box -38 -48 406 592
use scs8hd_fill_2  FILLER_37_266
timestamp 1586364061
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_37_270
timestamp 1586364061
transform 1 0 25944 0 1 22304
box -38 -48 590 592
use scs8hd_fill_1  FILLER_37_276
timestamp 1586364061
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 10212 0 -1 23392
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 590 592
use scs8hd_decap_4  FILLER_38_118
timestamp 1586364061
transform 1 0 11960 0 -1 23392
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_122
timestamp 1586364061
transform 1 0 12328 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_125
timestamp 1586364061
transform 1 0 12604 0 -1 23392
box -38 -48 130 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_145
timestamp 1586364061
transform 1 0 14444 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_8  FILLER_38_157
timestamp 1586364061
transform 1 0 15548 0 -1 23392
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_right_track_4.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 16652 0 -1 23392
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_165
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_168
timestamp 1586364061
transform 1 0 16560 0 -1 23392
box -38 -48 130 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_1_
timestamp 1586364061
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_188
timestamp 1586364061
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_192
timestamp 1586364061
transform 1 0 18768 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_196
timestamp 1586364061
transform 1 0 19136 0 -1 23392
box -38 -48 130 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_38_206
timestamp 1586364061
transform 1 0 20056 0 -1 23392
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_0.mux_l1_in_1_
timestamp 1586364061
transform 1 0 22448 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_38_219
timestamp 1586364061
transform 1 0 21252 0 -1 23392
box -38 -48 774 592
use scs8hd_decap_3  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 314 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 23644 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 24012 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_241
timestamp 1586364061
transform 1 0 23276 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_38_247
timestamp 1586364061
transform 1 0 23828 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_259
timestamp 1586364061
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_38_271
timestamp 1586364061
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 9752 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_97
timestamp 1586364061
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_107
timestamp 1586364061
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_103
timestamp 1586364061
transform 1 0 10580 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_101
timestamp 1586364061
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_14.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_14.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_right_track_14.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11132 0 -1 24480
box -38 -48 1786 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 13616 0 -1 24480
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_14.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13432 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_132
timestamp 1586364061
transform 1 0 13248 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_136
timestamp 1586364061
transform 1 0 13616 0 1 23392
box -38 -48 406 592
use scs8hd_decap_6  FILLER_40_128
timestamp 1586364061
transform 1 0 12880 0 -1 24480
box -38 -48 590 592
use scs8hd_decap_4  FILLER_40_148
timestamp 1586364061
transform 1 0 14720 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_40_144
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_140
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14536 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14168 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_16.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 13984 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_158
timestamp 1586364061
transform 1 0 15640 0 -1 24480
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_16.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14168 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 16652 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_161
timestamp 1586364061
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_165
timestamp 1586364061
transform 1 0 16284 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_177
timestamp 1586364061
transform 1 0 17388 0 1 23392
box -38 -48 590 592
use scs8hd_decap_12  FILLER_40_170
timestamp 1586364061
transform 1 0 16744 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_40_182
timestamp 1586364061
transform 1 0 17848 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 18216 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_0_
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 19320 0 1 23392
box -38 -48 1786 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 19964 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_217
timestamp 1586364061
transform 1 0 21068 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_199
timestamp 1586364061
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_40_203
timestamp 1586364061
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_6  FILLER_40_207
timestamp 1586364061
transform 1 0 20148 0 -1 24480
box -38 -48 590 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_221
timestamp 1586364061
transform 1 0 21436 0 1 23392
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 21252 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 21804 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_40_231
timestamp 1586364061
transform 1 0 22356 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_237
timestamp 1586364061
transform 1 0 22908 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_233
timestamp 1586364061
transform 1 0 22540 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_229
timestamp 1586364061
transform 1 0 22172 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 22724 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 22356 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_219
timestamp 1586364061
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_right_track_2.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 22724 0 -1 24480
box -38 -48 1786 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_right_track_2.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_241
timestamp 1586364061
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_253
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_254
timestamp 1586364061
transform 1 0 24472 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_8  FILLER_40_266
timestamp 1586364061
transform 1 0 25576 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_263
timestamp 1586364061
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_259
timestamp 1586364061
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 25484 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 25208 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_274
timestamp 1586364061
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_275
timestamp 1586364061
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_267
timestamp 1586364061
transform 1 0 25668 0 1 23392
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use scs8hd_mux2_2  mux_right_track_16.mux_l1_in_0_
timestamp 1586364061
transform 1 0 14168 0 1 24480
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use scs8hd_fill_1  FILLER_41_139
timestamp 1586364061
transform 1 0 13892 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_151
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_163
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_175
timestamp 1586364061
transform 1 0 17204 0 1 24480
box -38 -48 774 592
use scs8hd_mux2_2  mux_right_track_2.mux_l1_in_1_
timestamp 1586364061
transform 1 0 19228 0 1 24480
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 18676 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18308 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_41_189
timestamp 1586364061
transform 1 0 18492 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_193
timestamp 1586364061
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_206
timestamp 1586364061
transform 1 0 20056 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_210
timestamp 1586364061
transform 1 0 20424 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_214
timestamp 1586364061
transform 1 0 20792 0 1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 22264 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_226
timestamp 1586364061
transform 1 0 21896 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_236
timestamp 1586364061
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_240
timestamp 1586364061
transform 1 0 23184 0 1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_259
timestamp 1586364061
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_263
timestamp 1586364061
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_41_275
timestamp 1586364061
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14168 0 -1 25568
box -38 -48 222 592
use scs8hd_fill_1  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_144
timestamp 1586364061
transform 1 0 14352 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_3  FILLER_42_152
timestamp 1586364061
transform 1 0 15088 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_mux2_2  mux_right_track_2.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18860 0 -1 25568
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_6  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_202
timestamp 1586364061
transform 1 0 19688 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_42_214
timestamp 1586364061
transform 1 0 20792 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_6  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 590 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_8  FILLER_42_240
timestamp 1586364061
transform 1 0 23184 0 -1 25568
box -38 -48 774 592
use scs8hd_decap_6  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_259
timestamp 1586364061
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_271
timestamp 1586364061
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 14002 0 14058 480 6 ccff_head
port 0 nsew default input
rlabel metal2 s 27526 27520 27582 28000 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 27520 12248 28000 12368 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 27520 17960 28000 18080 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 27520 19592 28000 19712 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 27520 20816 28000 20936 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 27520 21360 28000 21480 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 27520 21904 28000 22024 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 27520 23128 28000 23248 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 27520 12792 28000 12912 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 27520 13336 28000 13456 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 27520 14560 28000 14680 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 27520 15104 28000 15224 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 27520 15648 28000 15768 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 27520 16192 28000 16312 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 27520 16736 28000 16856 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 27520 17416 28000 17536 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 27520 824 28000 944 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 27520 6536 28000 6656 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 27520 7080 28000 7200 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 27520 7624 28000 7744 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 27520 8848 28000 8968 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 27520 10480 28000 10600 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 27520 11024 28000 11144 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 27520 11704 28000 11824 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 27520 2456 28000 2576 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 27520 4224 28000 4344 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 27520 4768 28000 4888 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 27520 5312 28000 5432 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 938 27520 994 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 8942 27520 8998 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10230 27520 10286 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11610 27520 11666 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 12898 27520 12954 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 13542 27520 13598 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1582 27520 1638 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 2226 27520 2282 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2870 27520 2926 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 6274 27520 6330 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 22190 27520 22246 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 22926 27520 22982 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25594 27520 25650 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26238 27520 26294 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 26882 27520 26938 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 15566 27520 15622 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 16854 27520 16910 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 18234 27520 18290 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 prog_clk
port 82 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 27520 23672 28000 23792 6 right_top_grid_pin_42_
port 84 nsew default input
rlabel metal3 s 27520 24216 28000 24336 6 right_top_grid_pin_43_
port 85 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 86 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 87 nsew default input
rlabel metal3 s 27520 25984 28000 26104 6 right_top_grid_pin_46_
port 88 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 89 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 90 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 91 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 93 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
