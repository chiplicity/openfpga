magic
tech EFS8A
magscale 1 2
timestamp 1603803895
<< locali >>
rect 4169 8279 4203 8381
rect 29101 7191 29135 7497
rect 32505 7191 32539 7293
rect 3525 5559 3559 5661
rect 30573 5151 30607 5253
rect 17601 3995 17635 4165
rect 10057 2975 10091 3145
rect 23213 2975 23247 3145
<< viali >>
rect 1593 13481 1627 13515
rect 1409 13345 1443 13379
rect 1593 12937 1627 12971
rect 2421 12937 2455 12971
rect 1409 12733 1443 12767
rect 24292 12733 24326 12767
rect 2053 12597 2087 12631
rect 24363 12597 24397 12631
rect 24777 12597 24811 12631
rect 35633 12393 35667 12427
rect 1752 12257 1786 12291
rect 2764 12257 2798 12291
rect 11044 12257 11078 12291
rect 19165 12257 19199 12291
rect 24108 12257 24142 12291
rect 25120 12257 25154 12291
rect 34412 12257 34446 12291
rect 35449 12257 35483 12291
rect 29561 12189 29595 12223
rect 1823 12053 1857 12087
rect 2835 12053 2869 12087
rect 10149 12053 10183 12087
rect 11115 12053 11149 12087
rect 19349 12053 19383 12087
rect 24179 12053 24213 12087
rect 25191 12053 25225 12087
rect 34483 12053 34517 12087
rect 1593 11849 1627 11883
rect 20867 11849 20901 11883
rect 31769 11849 31803 11883
rect 35357 11849 35391 11883
rect 35633 11849 35667 11883
rect 36691 11849 36725 11883
rect 2053 11781 2087 11815
rect 18797 11781 18831 11815
rect 3341 11713 3375 11747
rect 1409 11645 1443 11679
rect 2580 11645 2614 11679
rect 10333 11645 10367 11679
rect 10609 11645 10643 11679
rect 18613 11645 18647 11679
rect 19073 11645 19107 11679
rect 20796 11645 20830 11679
rect 24444 11645 24478 11679
rect 24869 11645 24903 11679
rect 30088 11645 30122 11679
rect 31284 11645 31318 11679
rect 33860 11645 33894 11679
rect 34253 11645 34287 11679
rect 35449 11645 35483 11679
rect 36001 11645 36035 11679
rect 36588 11645 36622 11679
rect 37013 11645 37047 11679
rect 10793 11577 10827 11611
rect 30573 11577 30607 11611
rect 34621 11577 34655 11611
rect 2421 11509 2455 11543
rect 2651 11509 2685 11543
rect 3065 11509 3099 11543
rect 9965 11509 9999 11543
rect 11161 11509 11195 11543
rect 15669 11509 15703 11543
rect 19441 11509 19475 11543
rect 19717 11509 19751 11543
rect 21281 11509 21315 11543
rect 24133 11509 24167 11543
rect 24547 11509 24581 11543
rect 25237 11509 25271 11543
rect 25421 11509 25455 11543
rect 30159 11509 30193 11543
rect 31355 11509 31389 11543
rect 33931 11509 33965 11543
rect 2697 11305 2731 11339
rect 10149 11305 10183 11339
rect 15761 11305 15795 11339
rect 26663 11305 26697 11339
rect 31493 11305 31527 11339
rect 35633 11305 35667 11339
rect 11621 11237 11655 11271
rect 21097 11237 21131 11271
rect 24409 11237 24443 11271
rect 24501 11237 24535 11271
rect 29837 11237 29871 11271
rect 29929 11237 29963 11271
rect 30481 11237 30515 11271
rect 1409 11169 1443 11203
rect 2519 11169 2553 11203
rect 4144 11169 4178 11203
rect 8585 11169 8619 11203
rect 10057 11169 10091 11203
rect 10425 11169 10459 11203
rect 13001 11169 13035 11203
rect 15485 11169 15519 11203
rect 15945 11169 15979 11203
rect 18220 11169 18254 11203
rect 19349 11169 19383 11203
rect 19625 11169 19659 11203
rect 23372 11169 23406 11203
rect 26592 11169 26626 11203
rect 28089 11169 28123 11203
rect 28273 11169 28307 11203
rect 32137 11169 32171 11203
rect 32597 11169 32631 11203
rect 34345 11169 34379 11203
rect 35449 11169 35483 11203
rect 36553 11169 36587 11203
rect 11529 11101 11563 11135
rect 11805 11101 11839 11135
rect 19901 11101 19935 11135
rect 21005 11101 21039 11135
rect 21649 11101 21683 11135
rect 25053 11101 25087 11135
rect 28549 11101 28583 11135
rect 32689 11101 32723 11135
rect 34989 11101 35023 11135
rect 1593 11033 1627 11067
rect 4215 11033 4249 11067
rect 8769 11033 8803 11067
rect 13185 11033 13219 11067
rect 18291 11033 18325 11067
rect 36737 11033 36771 11067
rect 10885 10965 10919 10999
rect 12541 10965 12575 10999
rect 20177 10965 20211 10999
rect 23443 10965 23477 10999
rect 27629 10965 27663 10999
rect 34529 10965 34563 10999
rect 35265 10965 35299 10999
rect 4813 10761 4847 10795
rect 8953 10761 8987 10795
rect 11529 10761 11563 10795
rect 16727 10761 16761 10795
rect 19809 10761 19843 10795
rect 21741 10761 21775 10795
rect 23121 10761 23155 10795
rect 24041 10761 24075 10795
rect 27077 10761 27111 10795
rect 29745 10761 29779 10795
rect 34345 10761 34379 10795
rect 35909 10761 35943 10795
rect 36645 10761 36679 10795
rect 37013 10761 37047 10795
rect 8309 10693 8343 10727
rect 29101 10693 29135 10727
rect 36277 10693 36311 10727
rect 9275 10625 9309 10659
rect 11805 10625 11839 10659
rect 15393 10625 15427 10659
rect 20085 10625 20119 10659
rect 20729 10625 20763 10659
rect 24593 10625 24627 10659
rect 25513 10625 25547 10659
rect 30481 10625 30515 10659
rect 31585 10625 31619 10659
rect 1409 10557 1443 10591
rect 2580 10557 2614 10591
rect 3065 10557 3099 10591
rect 3960 10557 3994 10591
rect 8125 10557 8159 10591
rect 8585 10557 8619 10591
rect 9188 10557 9222 10591
rect 9689 10557 9723 10591
rect 12725 10557 12759 10591
rect 13001 10557 13035 10591
rect 16624 10557 16658 10591
rect 17049 10557 17083 10591
rect 17877 10557 17911 10591
rect 18429 10557 18463 10591
rect 18981 10557 19015 10591
rect 21557 10557 21591 10591
rect 22017 10557 22051 10591
rect 22636 10557 22670 10591
rect 25973 10557 26007 10591
rect 26065 10557 26099 10591
rect 26525 10557 26559 10591
rect 27537 10557 27571 10591
rect 27629 10557 27663 10591
rect 28089 10557 28123 10591
rect 33057 10557 33091 10591
rect 33517 10557 33551 10591
rect 36461 10557 36495 10591
rect 37600 10557 37634 10591
rect 38025 10557 38059 10591
rect 10241 10489 10275 10523
rect 10333 10489 10367 10523
rect 10885 10489 10919 10523
rect 15117 10489 15151 10523
rect 15209 10489 15243 10523
rect 16129 10489 16163 10523
rect 19165 10489 19199 10523
rect 20177 10489 20211 10523
rect 24685 10489 24719 10523
rect 25237 10489 25271 10523
rect 28365 10489 28399 10523
rect 30021 10489 30055 10523
rect 30113 10489 30147 10523
rect 31309 10489 31343 10523
rect 31677 10489 31711 10523
rect 32229 10489 32263 10523
rect 33793 10489 33827 10523
rect 34989 10489 35023 10523
rect 35081 10489 35115 10523
rect 35633 10489 35667 10523
rect 1593 10421 1627 10455
rect 2053 10421 2087 10455
rect 2651 10421 2685 10455
rect 3433 10421 3467 10455
rect 4031 10421 4065 10455
rect 4445 10421 4479 10455
rect 6837 10421 6871 10455
rect 10057 10421 10091 10455
rect 12173 10421 12207 10455
rect 12541 10421 12575 10455
rect 13461 10421 13495 10455
rect 14013 10421 14047 10455
rect 14933 10421 14967 10455
rect 18245 10421 18279 10455
rect 19533 10421 19567 10455
rect 21005 10421 21039 10455
rect 21465 10421 21499 10455
rect 22707 10421 22741 10455
rect 23489 10421 23523 10455
rect 24409 10421 24443 10455
rect 26341 10421 26375 10455
rect 28641 10421 28675 10455
rect 31033 10421 31067 10455
rect 32505 10421 32539 10455
rect 32873 10421 32907 10455
rect 37703 10421 37737 10455
rect 2053 10217 2087 10251
rect 4951 10217 4985 10251
rect 9965 10217 9999 10251
rect 10333 10217 10367 10251
rect 15117 10217 15151 10251
rect 15577 10217 15611 10251
rect 19073 10217 19107 10251
rect 19441 10217 19475 10251
rect 20177 10217 20211 10251
rect 26157 10217 26191 10251
rect 27905 10217 27939 10251
rect 29469 10217 29503 10251
rect 31585 10217 31619 10251
rect 32689 10217 32723 10251
rect 34069 10217 34103 10251
rect 36277 10217 36311 10251
rect 36645 10217 36679 10251
rect 10609 10149 10643 10183
rect 12081 10149 12115 10183
rect 12173 10149 12207 10183
rect 12725 10149 12759 10183
rect 15945 10149 15979 10183
rect 16037 10149 16071 10183
rect 18705 10149 18739 10183
rect 21097 10149 21131 10183
rect 23213 10149 23247 10183
rect 23305 10149 23339 10183
rect 24501 10149 24535 10183
rect 24777 10149 24811 10183
rect 24869 10149 24903 10183
rect 26617 10149 26651 10183
rect 26709 10149 26743 10183
rect 28870 10149 28904 10183
rect 29745 10149 29779 10183
rect 30481 10149 30515 10183
rect 30573 10149 30607 10183
rect 33149 10149 33183 10183
rect 33701 10149 33735 10183
rect 34713 10149 34747 10183
rect 2145 10081 2179 10115
rect 2421 10081 2455 10115
rect 4880 10081 4914 10115
rect 7608 10081 7642 10115
rect 8620 10081 8654 10115
rect 13921 10081 13955 10115
rect 14197 10081 14231 10115
rect 17601 10081 17635 10115
rect 18153 10081 18187 10115
rect 19349 10081 19383 10115
rect 19717 10081 19751 10115
rect 21649 10081 21683 10115
rect 36093 10081 36127 10115
rect 1685 10013 1719 10047
rect 6561 10013 6595 10047
rect 10517 10013 10551 10047
rect 11161 10013 11195 10047
rect 14381 10013 14415 10047
rect 16221 10013 16255 10047
rect 18337 10013 18371 10047
rect 21005 10013 21039 10047
rect 23489 10013 23523 10047
rect 25053 10013 25087 10047
rect 26893 10013 26927 10047
rect 28549 10013 28583 10047
rect 31125 10013 31159 10047
rect 33057 10013 33091 10047
rect 34621 10013 34655 10047
rect 34897 10013 34931 10047
rect 7711 9877 7745 9911
rect 8723 9877 8757 9911
rect 9045 9877 9079 9911
rect 24133 9877 24167 9911
rect 30113 9877 30147 9911
rect 32413 9877 32447 9911
rect 5181 9673 5215 9707
rect 9597 9673 9631 9707
rect 11437 9673 11471 9707
rect 11805 9673 11839 9707
rect 13737 9673 13771 9707
rect 16221 9673 16255 9707
rect 18797 9673 18831 9707
rect 20177 9673 20211 9707
rect 21925 9673 21959 9707
rect 22753 9673 22787 9707
rect 24961 9673 24995 9707
rect 25237 9673 25271 9707
rect 30849 9673 30883 9707
rect 33241 9673 33275 9707
rect 33517 9673 33551 9707
rect 2053 9605 2087 9639
rect 3985 9605 4019 9639
rect 5871 9605 5905 9639
rect 11069 9605 11103 9639
rect 12173 9605 12207 9639
rect 13093 9605 13127 9639
rect 15945 9605 15979 9639
rect 16589 9605 16623 9639
rect 17877 9605 17911 9639
rect 23121 9605 23155 9639
rect 24593 9605 24627 9639
rect 27169 9605 27203 9639
rect 28733 9605 28767 9639
rect 30205 9605 30239 9639
rect 30573 9605 30607 9639
rect 31447 9605 31481 9639
rect 33977 9605 34011 9639
rect 2329 9537 2363 9571
rect 3249 9537 3283 9571
rect 6653 9537 6687 9571
rect 8677 9537 8711 9571
rect 9321 9537 9355 9571
rect 10149 9537 10183 9571
rect 12541 9537 12575 9571
rect 15025 9537 15059 9571
rect 19257 9537 19291 9571
rect 21005 9537 21039 9571
rect 22201 9537 22235 9571
rect 25513 9537 25547 9571
rect 25789 9537 25823 9571
rect 28365 9537 28399 9571
rect 29285 9537 29319 9571
rect 32321 9537 32355 9571
rect 34989 9537 35023 9571
rect 35265 9537 35299 9571
rect 36829 9537 36863 9571
rect 3709 9469 3743 9503
rect 4445 9469 4479 9503
rect 4629 9469 4663 9503
rect 5641 9469 5675 9503
rect 5768 9469 5802 9503
rect 6837 9469 6871 9503
rect 7297 9469 7331 9503
rect 14048 9469 14082 9503
rect 14473 9469 14507 9503
rect 16992 9469 17026 9503
rect 17417 9469 17451 9503
rect 18312 9469 18346 9503
rect 23673 9469 23707 9503
rect 27905 9469 27939 9503
rect 28089 9469 28123 9503
rect 31344 9469 31378 9503
rect 31861 9469 31895 9503
rect 36093 9469 36127 9503
rect 2421 9401 2455 9435
rect 2973 9401 3007 9435
rect 8769 9401 8803 9435
rect 10470 9401 10504 9435
rect 12633 9401 12667 9435
rect 14933 9401 14967 9435
rect 15387 9401 15421 9435
rect 19619 9401 19653 9435
rect 20913 9401 20947 9435
rect 21326 9401 21360 9435
rect 23994 9401 24028 9435
rect 25605 9401 25639 9435
rect 27537 9401 27571 9435
rect 29101 9401 29135 9435
rect 29647 9401 29681 9435
rect 32229 9401 32263 9435
rect 32683 9401 32717 9435
rect 34713 9401 34747 9435
rect 35081 9401 35115 9435
rect 36553 9401 36587 9435
rect 36645 9401 36679 9435
rect 1685 9333 1719 9367
rect 4261 9333 4295 9367
rect 6193 9333 6227 9367
rect 6929 9333 6963 9367
rect 7849 9333 7883 9367
rect 8401 9333 8435 9367
rect 9965 9333 9999 9367
rect 14151 9333 14185 9367
rect 17095 9333 17129 9367
rect 18383 9333 18417 9367
rect 19165 9333 19199 9367
rect 20545 9333 20579 9367
rect 23489 9333 23523 9367
rect 26525 9333 26559 9367
rect 34345 9333 34379 9367
rect 7573 9129 7607 9163
rect 8125 9129 8159 9163
rect 10149 9129 10183 9163
rect 10885 9129 10919 9163
rect 11989 9129 12023 9163
rect 12541 9129 12575 9163
rect 15025 9129 15059 9163
rect 16681 9129 16715 9163
rect 17601 9129 17635 9163
rect 18705 9129 18739 9163
rect 20729 9129 20763 9163
rect 21833 9129 21867 9163
rect 25053 9129 25087 9163
rect 26617 9129 26651 9163
rect 28549 9129 28583 9163
rect 29561 9129 29595 9163
rect 35265 9129 35299 9163
rect 36369 9129 36403 9163
rect 36737 9129 36771 9163
rect 2605 9061 2639 9095
rect 5089 9061 5123 9095
rect 6561 9061 6595 9095
rect 6653 9061 6687 9095
rect 9827 9061 9861 9095
rect 11390 9061 11424 9095
rect 13829 9061 13863 9095
rect 14381 9061 14415 9095
rect 16082 9061 16116 9095
rect 18981 9061 19015 9095
rect 19073 9061 19107 9095
rect 23029 9061 23063 9095
rect 24178 9061 24212 9095
rect 25513 9061 25547 9095
rect 29003 9061 29037 9095
rect 31217 9061 31251 9095
rect 33149 9061 33183 9095
rect 34063 9061 34097 9095
rect 35811 9061 35845 9095
rect 1476 8993 1510 9027
rect 8125 8993 8159 9027
rect 8493 8993 8527 9027
rect 9724 8993 9758 9027
rect 11069 8993 11103 9027
rect 15761 8993 15795 9027
rect 17912 8993 17946 9027
rect 20948 8993 20982 9027
rect 22569 8993 22603 9027
rect 22753 8993 22787 9027
rect 24777 8993 24811 9027
rect 26525 8993 26559 9027
rect 26985 8993 27019 9027
rect 28641 8993 28675 9027
rect 30481 8993 30515 9027
rect 30941 8993 30975 9027
rect 32137 8993 32171 9027
rect 32597 8993 32631 9027
rect 34621 8993 34655 9027
rect 2513 8925 2547 8959
rect 2881 8925 2915 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 6837 8925 6871 8959
rect 13737 8925 13771 8959
rect 19993 8925 20027 8959
rect 23857 8925 23891 8959
rect 26341 8925 26375 8959
rect 32873 8925 32907 8959
rect 33517 8925 33551 8959
rect 33701 8925 33735 8959
rect 35449 8925 35483 8959
rect 18015 8857 18049 8891
rect 19533 8857 19567 8891
rect 1547 8789 1581 8823
rect 1869 8789 1903 8823
rect 2329 8789 2363 8823
rect 9137 8789 9171 8823
rect 10609 8789 10643 8823
rect 12817 8789 12851 8823
rect 13553 8789 13587 8823
rect 18429 8789 18463 8823
rect 21051 8789 21085 8823
rect 21557 8789 21591 8823
rect 23673 8789 23707 8823
rect 27721 8789 27755 8823
rect 30113 8789 30147 8823
rect 34897 8789 34931 8823
rect 1593 8585 1627 8619
rect 3249 8585 3283 8619
rect 3985 8585 4019 8619
rect 6285 8585 6319 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 9183 8585 9217 8619
rect 9873 8585 9907 8619
rect 10977 8585 11011 8619
rect 11713 8585 11747 8619
rect 13737 8585 13771 8619
rect 14013 8585 14047 8619
rect 17325 8585 17359 8619
rect 17877 8585 17911 8619
rect 19257 8585 19291 8619
rect 20637 8585 20671 8619
rect 21373 8585 21407 8619
rect 22845 8585 22879 8619
rect 24593 8585 24627 8619
rect 24961 8585 24995 8619
rect 25513 8585 25547 8619
rect 27077 8585 27111 8619
rect 29009 8585 29043 8619
rect 31723 8585 31757 8619
rect 32137 8585 32171 8619
rect 34069 8585 34103 8619
rect 35909 8585 35943 8619
rect 36277 8585 36311 8619
rect 36645 8585 36679 8619
rect 2881 8517 2915 8551
rect 15485 8517 15519 8551
rect 16129 8517 16163 8551
rect 21005 8517 21039 8551
rect 27445 8517 27479 8551
rect 2329 8449 2363 8483
rect 3617 8449 3651 8483
rect 5089 8449 5123 8483
rect 5549 8449 5583 8483
rect 6929 8449 6963 8483
rect 10057 8449 10091 8483
rect 12817 8449 12851 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 19717 8449 19751 8483
rect 25789 8449 25823 8483
rect 26433 8449 26467 8483
rect 31033 8449 31067 8483
rect 32781 8449 32815 8483
rect 34989 8449 35023 8483
rect 35265 8449 35299 8483
rect 3801 8381 3835 8415
rect 4169 8381 4203 8415
rect 7849 8381 7883 8415
rect 9080 8381 9114 8415
rect 9505 8381 9539 8415
rect 14565 8381 14599 8415
rect 16313 8381 16347 8415
rect 16865 8381 16899 8415
rect 21465 8381 21499 8415
rect 21925 8381 21959 8415
rect 23673 8381 23707 8415
rect 27629 8381 27663 8415
rect 28089 8381 28123 8415
rect 28365 8381 28399 8415
rect 31620 8381 31654 8415
rect 33701 8381 33735 8415
rect 34621 8381 34655 8415
rect 36461 8381 36495 8415
rect 37013 8381 37047 8415
rect 2145 8313 2179 8347
rect 2421 8313 2455 8347
rect 5273 8313 5307 8347
rect 5365 8313 5399 8347
rect 6653 8313 6687 8347
rect 7250 8313 7284 8347
rect 10378 8313 10412 8347
rect 11253 8313 11287 8347
rect 12725 8313 12759 8347
rect 13179 8313 13213 8347
rect 14473 8313 14507 8347
rect 14927 8313 14961 8347
rect 17049 8313 17083 8347
rect 18337 8313 18371 8347
rect 20038 8313 20072 8347
rect 22569 8313 22603 8347
rect 23994 8313 24028 8347
rect 25881 8313 25915 8347
rect 26709 8313 26743 8347
rect 28733 8313 28767 8347
rect 29929 8313 29963 8347
rect 30113 8313 30147 8347
rect 30205 8313 30239 8347
rect 30757 8313 30791 8347
rect 31401 8313 31435 8347
rect 32689 8313 32723 8347
rect 33143 8313 33177 8347
rect 35081 8313 35115 8347
rect 4169 8245 4203 8279
rect 4445 8245 4479 8279
rect 15761 8245 15795 8279
rect 19625 8245 19659 8279
rect 21557 8245 21591 8279
rect 23489 8245 23523 8279
rect 2697 8041 2731 8075
rect 3893 8041 3927 8075
rect 5181 8041 5215 8075
rect 5549 8041 5583 8075
rect 5825 8041 5859 8075
rect 6561 8041 6595 8075
rect 7757 8041 7791 8075
rect 8723 8041 8757 8075
rect 10793 8041 10827 8075
rect 13185 8041 13219 8075
rect 16957 8041 16991 8075
rect 18521 8041 18555 8075
rect 20085 8041 20119 8075
rect 23857 8041 23891 8075
rect 25421 8041 25455 8075
rect 25789 8041 25823 8075
rect 29837 8041 29871 8075
rect 30481 8041 30515 8075
rect 30665 8041 30699 8075
rect 32413 8041 32447 8075
rect 34437 8041 34471 8075
rect 2139 7973 2173 8007
rect 4261 7973 4295 8007
rect 4813 7973 4847 8007
rect 7199 7973 7233 8007
rect 14381 7973 14415 8007
rect 14657 7973 14691 8007
rect 15663 7973 15697 8007
rect 17693 7973 17727 8007
rect 19266 7973 19300 8007
rect 21649 7973 21683 8007
rect 24822 7973 24856 8007
rect 26887 7973 26921 8007
rect 29238 7973 29272 8007
rect 33879 7973 33913 8007
rect 35449 7973 35483 8007
rect 36001 7973 36035 8007
rect 1777 7905 1811 7939
rect 5641 7905 5675 7939
rect 8652 7905 8686 7939
rect 10793 7905 10827 7939
rect 10977 7905 11011 7939
rect 12357 7905 12391 7939
rect 12633 7905 12667 7939
rect 13829 7905 13863 7939
rect 14105 7905 14139 7939
rect 16221 7905 16255 7939
rect 18889 7905 18923 7939
rect 23029 7905 23063 7939
rect 23213 7905 23247 7939
rect 30113 7905 30147 7939
rect 32572 7905 32606 7939
rect 3525 7837 3559 7871
rect 4169 7837 4203 7871
rect 6837 7837 6871 7871
rect 12817 7837 12851 7871
rect 15301 7837 15335 7871
rect 17601 7837 17635 7871
rect 18245 7837 18279 7871
rect 19165 7837 19199 7871
rect 19533 7837 19567 7871
rect 21281 7837 21315 7871
rect 21557 7837 21591 7871
rect 23581 7837 23615 7871
rect 24501 7837 24535 7871
rect 26525 7837 26559 7871
rect 28917 7837 28951 7871
rect 33517 7837 33551 7871
rect 35357 7837 35391 7871
rect 22109 7769 22143 7803
rect 33333 7769 33367 7803
rect 3065 7701 3099 7735
rect 10057 7701 10091 7735
rect 13553 7701 13587 7735
rect 16589 7701 16623 7735
rect 24225 7701 24259 7735
rect 27445 7701 27479 7735
rect 27721 7701 27755 7735
rect 32643 7701 32677 7735
rect 34897 7701 34931 7735
rect 3157 7497 3191 7531
rect 5733 7497 5767 7531
rect 8769 7497 8803 7531
rect 9689 7497 9723 7531
rect 11161 7497 11195 7531
rect 11805 7497 11839 7531
rect 13461 7497 13495 7531
rect 14565 7497 14599 7531
rect 15301 7497 15335 7531
rect 17601 7497 17635 7531
rect 20085 7497 20119 7531
rect 22385 7497 22419 7531
rect 29101 7497 29135 7531
rect 31033 7497 31067 7531
rect 32781 7497 32815 7531
rect 34253 7497 34287 7531
rect 35909 7497 35943 7531
rect 36645 7497 36679 7531
rect 9965 7429 9999 7463
rect 12173 7429 12207 7463
rect 19257 7429 19291 7463
rect 4169 7361 4203 7395
rect 10517 7361 10551 7395
rect 13921 7361 13955 7395
rect 16221 7361 16255 7395
rect 18705 7361 18739 7395
rect 20315 7361 20349 7395
rect 21465 7361 21499 7395
rect 24225 7361 24259 7395
rect 25881 7361 25915 7395
rect 27721 7361 27755 7395
rect 28089 7361 28123 7395
rect 2237 7293 2271 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 7849 7293 7883 7327
rect 12608 7293 12642 7327
rect 15117 7293 15151 7327
rect 17141 7293 17175 7327
rect 18429 7293 18463 7327
rect 20212 7293 20246 7327
rect 20637 7293 20671 7327
rect 23121 7293 23155 7327
rect 23489 7293 23523 7327
rect 23949 7293 23983 7327
rect 24133 7293 24167 7327
rect 26801 7293 26835 7327
rect 27445 7293 27479 7327
rect 2558 7225 2592 7259
rect 4490 7225 4524 7259
rect 8170 7225 8204 7259
rect 10241 7225 10275 7259
rect 10333 7225 10367 7259
rect 13645 7225 13679 7259
rect 13737 7225 13771 7259
rect 15669 7225 15703 7259
rect 16129 7225 16163 7259
rect 16583 7225 16617 7259
rect 18797 7225 18831 7259
rect 21373 7225 21407 7259
rect 21827 7225 21861 7259
rect 25697 7225 25731 7259
rect 26202 7225 26236 7259
rect 27077 7225 27111 7259
rect 27813 7225 27847 7259
rect 32367 7429 32401 7463
rect 30113 7361 30147 7395
rect 33333 7361 33367 7395
rect 34989 7361 35023 7395
rect 35357 7361 35391 7395
rect 32296 7293 32330 7327
rect 32505 7293 32539 7327
rect 33977 7293 34011 7327
rect 36461 7293 36495 7327
rect 37013 7293 37047 7327
rect 29469 7225 29503 7259
rect 30021 7225 30055 7259
rect 30475 7225 30509 7259
rect 1869 7157 1903 7191
rect 3525 7157 3559 7191
rect 3985 7157 4019 7191
rect 5089 7157 5123 7191
rect 6285 7157 6319 7191
rect 7021 7157 7055 7191
rect 7297 7157 7331 7191
rect 7665 7157 7699 7191
rect 9321 7157 9355 7191
rect 12679 7157 12713 7191
rect 13093 7157 13127 7191
rect 14933 7157 14967 7191
rect 19625 7157 19659 7191
rect 22661 7157 22695 7191
rect 24685 7157 24719 7191
rect 25053 7157 25087 7191
rect 29009 7157 29043 7191
rect 29101 7157 29135 7191
rect 33434 7225 33468 7259
rect 34621 7225 34655 7259
rect 35081 7225 35115 7259
rect 32505 7157 32539 7191
rect 33149 7157 33183 7191
rect 1777 6953 1811 6987
rect 10609 6953 10643 6987
rect 13737 6953 13771 6987
rect 17509 6953 17543 6987
rect 22017 6953 22051 6987
rect 25973 6953 26007 6987
rect 33885 6953 33919 6987
rect 35449 6953 35483 6987
rect 2558 6885 2592 6919
rect 4537 6885 4571 6919
rect 6923 6885 6957 6919
rect 10010 6885 10044 6919
rect 12351 6885 12385 6919
rect 15853 6885 15887 6919
rect 16129 6885 16163 6919
rect 19343 6885 19377 6919
rect 21097 6885 21131 6919
rect 24501 6885 24535 6919
rect 27261 6885 27295 6919
rect 27813 6885 27847 6919
rect 28825 6885 28859 6919
rect 32499 6885 32533 6919
rect 34621 6885 34655 6919
rect 35173 6885 35207 6919
rect 36185 6885 36219 6919
rect 3893 6817 3927 6851
rect 8585 6817 8619 6851
rect 14197 6817 14231 6851
rect 16681 6817 16715 6851
rect 17601 6817 17635 6851
rect 17785 6817 17819 6851
rect 18521 6817 18555 6851
rect 19901 6817 19935 6851
rect 22512 6817 22546 6851
rect 24041 6817 24075 6851
rect 24317 6817 24351 6851
rect 25329 6817 25363 6851
rect 30389 6817 30423 6851
rect 30757 6817 30791 6851
rect 30941 6817 30975 6851
rect 2237 6749 2271 6783
rect 4445 6749 4479 6783
rect 6561 6749 6595 6783
rect 9689 6749 9723 6783
rect 11989 6749 12023 6783
rect 16037 6749 16071 6783
rect 18153 6749 18187 6783
rect 18981 6749 19015 6783
rect 20729 6749 20763 6783
rect 21005 6749 21039 6783
rect 21649 6749 21683 6783
rect 27169 6749 27203 6783
rect 28549 6749 28583 6783
rect 28733 6749 28767 6783
rect 29101 6749 29135 6783
rect 31217 6749 31251 6783
rect 32137 6749 32171 6783
rect 34529 6749 34563 6783
rect 36093 6749 36127 6783
rect 36369 6749 36403 6783
rect 4997 6681 5031 6715
rect 8769 6681 8803 6715
rect 14381 6681 14415 6715
rect 25513 6681 25547 6715
rect 3157 6613 3191 6647
rect 3433 6613 3467 6647
rect 7481 6613 7515 6647
rect 7941 6613 7975 6647
rect 9045 6613 9079 6647
rect 12909 6613 12943 6647
rect 14013 6613 14047 6647
rect 16957 6613 16991 6647
rect 18889 6613 18923 6647
rect 22293 6613 22327 6647
rect 22615 6613 22649 6647
rect 26709 6613 26743 6647
rect 33057 6613 33091 6647
rect 33517 6613 33551 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 4169 6409 4203 6443
rect 5273 6409 5307 6443
rect 6561 6409 6595 6443
rect 8309 6409 8343 6443
rect 12081 6409 12115 6443
rect 13369 6409 13403 6443
rect 16313 6409 16347 6443
rect 16589 6409 16623 6443
rect 16957 6409 16991 6443
rect 17693 6409 17727 6443
rect 21189 6409 21223 6443
rect 21833 6409 21867 6443
rect 23121 6409 23155 6443
rect 24961 6409 24995 6443
rect 25329 6409 25363 6443
rect 27169 6409 27203 6443
rect 28733 6409 28767 6443
rect 30573 6409 30607 6443
rect 32229 6409 32263 6443
rect 32505 6409 32539 6443
rect 33885 6409 33919 6443
rect 36599 6409 36633 6443
rect 3341 6341 3375 6375
rect 24593 6341 24627 6375
rect 34253 6341 34287 6375
rect 36001 6341 36035 6375
rect 2789 6273 2823 6307
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 6285 6273 6319 6307
rect 7573 6273 7607 6307
rect 11069 6273 11103 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 27721 6273 27755 6307
rect 27997 6273 28031 6307
rect 29653 6273 29687 6307
rect 35357 6273 35391 6307
rect 1409 6205 1443 6239
rect 8677 6205 8711 6239
rect 8861 6205 8895 6239
rect 12449 6205 12483 6239
rect 13645 6205 13679 6239
rect 14105 6205 14139 6239
rect 14197 6205 14231 6239
rect 15393 6205 15427 6239
rect 19993 6205 20027 6239
rect 22017 6205 22051 6239
rect 22569 6205 22603 6239
rect 23673 6205 23707 6239
rect 25881 6205 25915 6239
rect 31033 6205 31067 6239
rect 31401 6205 31435 6239
rect 31585 6205 31619 6239
rect 31861 6205 31895 6239
rect 32689 6205 32723 6239
rect 33609 6205 33643 6239
rect 34621 6205 34655 6239
rect 36496 6205 36530 6239
rect 36921 6205 36955 6239
rect 2329 6137 2363 6171
rect 2881 6137 2915 6171
rect 4445 6137 4479 6171
rect 6929 6137 6963 6171
rect 7021 6137 7055 6171
rect 10793 6137 10827 6171
rect 10885 6137 10919 6171
rect 12811 6137 12845 6171
rect 15301 6137 15335 6171
rect 15755 6137 15789 6171
rect 18613 6137 18647 6171
rect 19533 6137 19567 6171
rect 19901 6137 19935 6171
rect 20355 6137 20389 6171
rect 23994 6137 24028 6171
rect 26202 6137 26236 6171
rect 27813 6137 27847 6171
rect 29377 6137 29411 6171
rect 29469 6137 29503 6171
rect 33010 6137 33044 6171
rect 34989 6137 35023 6171
rect 35081 6137 35115 6171
rect 3709 6069 3743 6103
rect 7849 6069 7883 6103
rect 8493 6069 8527 6103
rect 9781 6069 9815 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 14381 6069 14415 6103
rect 14749 6069 14783 6103
rect 18337 6069 18371 6103
rect 20913 6069 20947 6103
rect 22293 6069 22327 6103
rect 23397 6069 23431 6103
rect 25697 6069 25731 6103
rect 26801 6069 26835 6103
rect 27537 6069 27571 6103
rect 29101 6069 29135 6103
rect 2973 5865 3007 5899
rect 5089 5865 5123 5899
rect 6745 5865 6779 5899
rect 7297 5865 7331 5899
rect 8493 5865 8527 5899
rect 10609 5865 10643 5899
rect 11989 5865 12023 5899
rect 13185 5865 13219 5899
rect 13553 5865 13587 5899
rect 16497 5865 16531 5899
rect 18521 5865 18555 5899
rect 19901 5865 19935 5899
rect 22109 5865 22143 5899
rect 24409 5865 24443 5899
rect 26341 5865 26375 5899
rect 31125 5865 31159 5899
rect 32689 5865 32723 5899
rect 33563 5865 33597 5899
rect 34253 5865 34287 5899
rect 35449 5865 35483 5899
rect 36461 5865 36495 5899
rect 2053 5797 2087 5831
rect 4261 5797 4295 5831
rect 5825 5797 5859 5831
rect 7113 5797 7147 5831
rect 10010 5797 10044 5831
rect 12265 5797 12299 5831
rect 13737 5797 13771 5831
rect 13829 5797 13863 5831
rect 15485 5797 15519 5831
rect 16957 5797 16991 5831
rect 17049 5797 17083 5831
rect 18975 5797 19009 5831
rect 21097 5797 21131 5831
rect 21649 5797 21683 5831
rect 22477 5797 22511 5831
rect 23534 5797 23568 5831
rect 27169 5797 27203 5831
rect 27721 5797 27755 5831
rect 28733 5797 28767 5831
rect 30849 5797 30883 5831
rect 34621 5797 34655 5831
rect 35173 5797 35207 5831
rect 7481 5729 7515 5763
rect 7757 5729 7791 5763
rect 18613 5729 18647 5763
rect 24961 5729 24995 5763
rect 25145 5729 25179 5763
rect 30113 5729 30147 5763
rect 30665 5729 30699 5763
rect 32204 5729 32238 5763
rect 33460 5729 33494 5763
rect 36036 5729 36070 5763
rect 1961 5661 1995 5695
rect 3525 5661 3559 5695
rect 4169 5661 4203 5695
rect 4445 5661 4479 5695
rect 5733 5661 5767 5695
rect 6009 5661 6043 5695
rect 9689 5661 9723 5695
rect 12173 5661 12207 5695
rect 14381 5661 14415 5695
rect 15393 5661 15427 5695
rect 15669 5661 15703 5695
rect 17233 5661 17267 5695
rect 21005 5661 21039 5695
rect 23213 5661 23247 5695
rect 25513 5661 25547 5695
rect 26893 5661 26927 5695
rect 27077 5661 27111 5695
rect 28641 5661 28675 5695
rect 29101 5661 29135 5695
rect 34529 5661 34563 5695
rect 36139 5661 36173 5695
rect 2513 5593 2547 5627
rect 10885 5593 10919 5627
rect 12725 5593 12759 5627
rect 17969 5593 18003 5627
rect 19533 5593 19567 5627
rect 24133 5593 24167 5627
rect 29653 5593 29687 5627
rect 32275 5593 32309 5627
rect 1685 5525 1719 5559
rect 3249 5525 3283 5559
rect 3525 5525 3559 5559
rect 3709 5525 3743 5559
rect 8769 5525 8803 5559
rect 14749 5525 14783 5559
rect 15117 5525 15151 5559
rect 20177 5525 20211 5559
rect 20729 5525 20763 5559
rect 25881 5525 25915 5559
rect 28089 5525 28123 5559
rect 2513 5321 2547 5355
rect 4629 5321 4663 5355
rect 4997 5321 5031 5355
rect 5641 5321 5675 5355
rect 5917 5321 5951 5355
rect 6653 5321 6687 5355
rect 7297 5321 7331 5355
rect 9137 5321 9171 5355
rect 10425 5321 10459 5355
rect 12173 5321 12207 5355
rect 14105 5321 14139 5355
rect 14473 5321 14507 5355
rect 17325 5321 17359 5355
rect 18337 5321 18371 5355
rect 19349 5321 19383 5355
rect 20545 5321 20579 5355
rect 20913 5321 20947 5355
rect 22477 5321 22511 5355
rect 24777 5321 24811 5355
rect 25145 5321 25179 5355
rect 26249 5321 26283 5355
rect 26893 5321 26927 5355
rect 29423 5321 29457 5355
rect 29745 5321 29779 5355
rect 30113 5321 30147 5355
rect 30435 5321 30469 5355
rect 32229 5321 32263 5355
rect 33425 5321 33459 5355
rect 34161 5321 34195 5355
rect 34529 5321 34563 5355
rect 35035 5321 35069 5355
rect 8033 5253 8067 5287
rect 13737 5253 13771 5287
rect 30573 5253 30607 5287
rect 30849 5253 30883 5287
rect 14749 5185 14783 5219
rect 15393 5185 15427 5219
rect 16773 5185 16807 5219
rect 20177 5185 20211 5219
rect 25881 5185 25915 5219
rect 27813 5185 27847 5219
rect 29009 5185 29043 5219
rect 31447 5185 31481 5219
rect 1593 5117 1627 5151
rect 2789 5117 2823 5151
rect 3709 5117 3743 5151
rect 5733 5117 5767 5151
rect 7113 5117 7147 5151
rect 7573 5117 7607 5151
rect 8217 5117 8251 5151
rect 10609 5117 10643 5151
rect 16221 5117 16255 5151
rect 16681 5117 16715 5151
rect 18245 5117 18279 5151
rect 19717 5117 19751 5151
rect 19993 5117 20027 5151
rect 21741 5117 21775 5151
rect 23673 5117 23707 5151
rect 24225 5117 24259 5151
rect 25237 5117 25271 5151
rect 25789 5117 25823 5151
rect 29352 5117 29386 5151
rect 30364 5117 30398 5151
rect 30573 5117 30607 5151
rect 31344 5117 31378 5151
rect 34964 5117 34998 5151
rect 1914 5049 1948 5083
rect 4071 5049 4105 5083
rect 6285 5049 6319 5083
rect 8538 5049 8572 5083
rect 9689 5049 9723 5083
rect 10930 5049 10964 5083
rect 13185 5049 13219 5083
rect 13277 5049 13311 5083
rect 14841 5049 14875 5083
rect 16129 5049 16163 5083
rect 18061 5049 18095 5083
rect 21281 5049 21315 5083
rect 22937 5049 22971 5083
rect 27169 5049 27203 5083
rect 27261 5049 27295 5083
rect 3249 4981 3283 5015
rect 3617 4981 3651 5015
rect 10057 4981 10091 5015
rect 11529 4981 11563 5015
rect 13001 4981 13035 5015
rect 15669 4981 15703 5015
rect 17785 4981 17819 5015
rect 18981 4981 19015 5015
rect 23305 4981 23339 5015
rect 23765 4981 23799 5015
rect 28181 4981 28215 5015
rect 28549 4981 28583 5015
rect 31769 4981 31803 5015
rect 35449 4981 35483 5015
rect 36001 4981 36035 5015
rect 1961 4777 1995 4811
rect 2237 4777 2271 4811
rect 3801 4777 3835 4811
rect 4169 4777 4203 4811
rect 7665 4777 7699 4811
rect 10701 4777 10735 4811
rect 12357 4777 12391 4811
rect 13461 4777 13495 4811
rect 14749 4777 14783 4811
rect 17785 4777 17819 4811
rect 19349 4777 19383 4811
rect 19993 4777 20027 4811
rect 20729 4777 20763 4811
rect 20913 4777 20947 4811
rect 23673 4777 23707 4811
rect 25789 4777 25823 4811
rect 27629 4777 27663 4811
rect 29791 4777 29825 4811
rect 30205 4777 30239 4811
rect 2605 4709 2639 4743
rect 6377 4709 6411 4743
rect 8861 4709 8895 4743
rect 13829 4709 13863 4743
rect 14381 4709 14415 4743
rect 15117 4709 15151 4743
rect 16681 4709 16715 4743
rect 18981 4709 19015 4743
rect 25513 4709 25547 4743
rect 28825 4709 28859 4743
rect 1476 4641 1510 4675
rect 4353 4641 4387 4675
rect 4537 4641 4571 4675
rect 5549 4641 5583 4675
rect 5641 4641 5675 4675
rect 5887 4641 5921 4675
rect 7205 4641 7239 4675
rect 7481 4641 7515 4675
rect 9689 4641 9723 4675
rect 9965 4641 9999 4675
rect 12265 4641 12299 4675
rect 12633 4641 12667 4675
rect 15301 4641 15335 4675
rect 15485 4641 15519 4675
rect 15853 4641 15887 4675
rect 16828 4641 16862 4675
rect 18061 4641 18095 4675
rect 18245 4641 18279 4675
rect 18797 4641 18831 4675
rect 19809 4641 19843 4675
rect 20269 4641 20303 4675
rect 22385 4641 22419 4675
rect 22937 4641 22971 4675
rect 25053 4641 25087 4675
rect 25329 4641 25363 4675
rect 27169 4641 27203 4675
rect 28089 4641 28123 4675
rect 28641 4641 28675 4675
rect 29720 4641 29754 4675
rect 2513 4573 2547 4607
rect 2973 4573 3007 4607
rect 10149 4573 10183 4607
rect 13737 4573 13771 4607
rect 17049 4573 17083 4607
rect 17141 4573 17175 4607
rect 22845 4573 22879 4607
rect 26525 4573 26559 4607
rect 5733 4505 5767 4539
rect 7021 4505 7055 4539
rect 7297 4505 7331 4539
rect 9781 4505 9815 4539
rect 1547 4437 1581 4471
rect 8401 4437 8435 4471
rect 9505 4437 9539 4471
rect 11897 4437 11931 4471
rect 13093 4437 13127 4471
rect 16497 4437 16531 4471
rect 16957 4437 16991 4471
rect 19717 4437 19751 4471
rect 21741 4437 21775 4471
rect 23213 4437 23247 4471
rect 24501 4437 24535 4471
rect 1685 4233 1719 4267
rect 4813 4233 4847 4267
rect 5273 4233 5307 4267
rect 7113 4233 7147 4267
rect 11897 4233 11931 4267
rect 13737 4233 13771 4267
rect 16313 4233 16347 4267
rect 19901 4233 19935 4267
rect 24041 4233 24075 4267
rect 25789 4233 25823 4267
rect 27261 4233 27295 4267
rect 27721 4233 27755 4267
rect 27997 4233 28031 4267
rect 30205 4233 30239 4267
rect 5641 4165 5675 4199
rect 16681 4165 16715 4199
rect 17601 4165 17635 4199
rect 19533 4165 19567 4199
rect 19763 4165 19797 4199
rect 1961 4097 1995 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 11345 4097 11379 4131
rect 12173 4097 12207 4131
rect 13001 4097 13035 4131
rect 15577 4097 15611 4131
rect 16773 4097 16807 4131
rect 17049 4097 17083 4131
rect 3341 4029 3375 4063
rect 3709 4029 3743 4063
rect 3985 4029 4019 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 7481 4029 7515 4063
rect 8401 4029 8435 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9781 4029 9815 4063
rect 10149 4029 10183 4063
rect 10517 4029 10551 4063
rect 12449 4029 12483 4063
rect 12909 4029 12943 4063
rect 14749 4029 14783 4063
rect 15393 4029 15427 4063
rect 16405 4029 16439 4063
rect 16552 4029 16586 4063
rect 17877 4097 17911 4131
rect 18153 4097 18187 4131
rect 19993 4097 20027 4131
rect 20085 4097 20119 4131
rect 23489 4097 23523 4131
rect 26157 4097 26191 4131
rect 28273 4097 28307 4131
rect 29423 4097 29457 4131
rect 18061 4029 18095 4063
rect 18291 4029 18325 4063
rect 19073 4029 19107 4063
rect 21465 4029 21499 4063
rect 21649 4029 21683 4063
rect 22293 4029 22327 4063
rect 22477 4029 22511 4063
rect 23029 4029 23063 4063
rect 24501 4029 24535 4063
rect 25421 4029 25455 4063
rect 27813 4029 27847 4063
rect 28641 4029 28675 4063
rect 29336 4029 29370 4063
rect 29837 4029 29871 4063
rect 30297 4029 30331 4063
rect 30757 4029 30791 4063
rect 2053 3961 2087 3995
rect 6193 3961 6227 3995
rect 17417 3961 17451 3995
rect 17601 3961 17635 3995
rect 18797 3961 18831 3995
rect 19625 3961 19659 3995
rect 20637 3961 20671 3995
rect 24409 3961 24443 3995
rect 24863 3961 24897 3995
rect 26341 3961 26375 3995
rect 26433 3961 26467 3995
rect 26985 3961 27019 3995
rect 3525 3893 3559 3927
rect 4445 3893 4479 3927
rect 5917 3893 5951 3927
rect 7849 3893 7883 3927
rect 8217 3893 8251 3927
rect 8861 3893 8895 3927
rect 10241 3893 10275 3927
rect 11069 3893 11103 3927
rect 14013 3893 14047 3927
rect 15853 3893 15887 3927
rect 21097 3893 21131 3927
rect 22753 3893 22787 3927
rect 30481 3893 30515 3927
rect 1777 3689 1811 3723
rect 2697 3689 2731 3723
rect 3065 3689 3099 3723
rect 3525 3689 3559 3723
rect 4215 3689 4249 3723
rect 5733 3689 5767 3723
rect 6561 3689 6595 3723
rect 8493 3689 8527 3723
rect 9229 3689 9263 3723
rect 9781 3689 9815 3723
rect 10701 3689 10735 3723
rect 12909 3689 12943 3723
rect 15853 3689 15887 3723
rect 16497 3689 16531 3723
rect 17049 3689 17083 3723
rect 17601 3689 17635 3723
rect 18429 3689 18463 3723
rect 20729 3689 20763 3723
rect 21005 3689 21039 3723
rect 23949 3689 23983 3723
rect 28641 3689 28675 3723
rect 5227 3621 5261 3655
rect 7297 3621 7331 3655
rect 12265 3621 12299 3655
rect 15577 3621 15611 3655
rect 17785 3621 17819 3655
rect 19901 3621 19935 3655
rect 24225 3621 24259 3655
rect 28083 3621 28117 3655
rect 29653 3621 29687 3655
rect 1961 3553 1995 3587
rect 2237 3553 2271 3587
rect 4144 3553 4178 3587
rect 5124 3553 5158 3587
rect 6377 3553 6411 3587
rect 7389 3553 7423 3587
rect 7665 3553 7699 3587
rect 9689 3553 9723 3587
rect 10287 3553 10321 3587
rect 11621 3553 11655 3587
rect 12633 3553 12667 3587
rect 13921 3553 13955 3587
rect 14013 3553 14047 3587
rect 14381 3553 14415 3587
rect 16313 3553 16347 3587
rect 17932 3553 17966 3587
rect 18797 3553 18831 3587
rect 19349 3553 19383 3587
rect 19533 3553 19567 3587
rect 20913 3553 20947 3587
rect 21373 3553 21407 3587
rect 21741 3553 21775 3587
rect 22753 3553 22787 3587
rect 22845 3553 22879 3587
rect 23673 3553 23707 3587
rect 23857 3553 23891 3587
rect 24869 3553 24903 3587
rect 26560 3553 26594 3587
rect 8125 3485 8159 3519
rect 18153 3485 18187 3519
rect 27721 3485 27755 3519
rect 29561 3485 29595 3519
rect 7481 3417 7515 3451
rect 18061 3417 18095 3451
rect 20177 3417 20211 3451
rect 30113 3417 30147 3451
rect 14933 3349 14967 3383
rect 19165 3349 19199 3383
rect 22293 3349 22327 3383
rect 24593 3349 24627 3383
rect 25237 3349 25271 3383
rect 26249 3349 26283 3383
rect 26663 3349 26697 3383
rect 26985 3349 27019 3383
rect 3847 3145 3881 3179
rect 4169 3145 4203 3179
rect 5089 3145 5123 3179
rect 5641 3145 5675 3179
rect 8769 3145 8803 3179
rect 10057 3145 10091 3179
rect 10333 3145 10367 3179
rect 11483 3145 11517 3179
rect 13185 3145 13219 3179
rect 13415 3145 13449 3179
rect 15117 3145 15151 3179
rect 15485 3145 15519 3179
rect 17785 3145 17819 3179
rect 18521 3145 18555 3179
rect 20269 3145 20303 3179
rect 23121 3145 23155 3179
rect 23213 3145 23247 3179
rect 23489 3145 23523 3179
rect 27261 3145 27295 3179
rect 27721 3145 27755 3179
rect 30757 3145 30791 3179
rect 3433 3077 3467 3111
rect 5917 3077 5951 3111
rect 6285 3077 6319 3111
rect 6653 3077 6687 3111
rect 7757 3077 7791 3111
rect 2605 3009 2639 3043
rect 4537 3009 4571 3043
rect 8125 3009 8159 3043
rect 9137 3009 9171 3043
rect 9781 3009 9815 3043
rect 10609 3077 10643 3111
rect 11805 3077 11839 3111
rect 12173 3077 12207 3111
rect 13829 3077 13863 3111
rect 16497 3077 16531 3111
rect 22477 3077 22511 3111
rect 14197 3009 14231 3043
rect 15209 3009 15243 3043
rect 17509 3009 17543 3043
rect 19349 3009 19383 3043
rect 22707 3009 22741 3043
rect 25605 3009 25639 3043
rect 26341 3009 26375 3043
rect 26985 3009 27019 3043
rect 29469 3009 29503 3043
rect 30113 3009 30147 3043
rect 30941 3009 30975 3043
rect 1777 2941 1811 2975
rect 1961 2941 1995 2975
rect 2513 2941 2547 2975
rect 2973 2941 3007 2975
rect 3776 2941 3810 2975
rect 5733 2941 5767 2975
rect 7389 2941 7423 2975
rect 7665 2941 7699 2975
rect 7941 2941 7975 2975
rect 9229 2941 9263 2975
rect 9689 2941 9723 2975
rect 10057 2941 10091 2975
rect 11412 2941 11446 2975
rect 13344 2941 13378 2975
rect 14749 2941 14783 2975
rect 14988 2941 15022 2975
rect 16037 2941 16071 2975
rect 16405 2941 16439 2975
rect 16681 2941 16715 2975
rect 17141 2941 17175 2975
rect 18061 2941 18095 2975
rect 19993 2941 20027 2975
rect 20821 2941 20855 2975
rect 21741 2941 21775 2975
rect 22017 2941 22051 2975
rect 22620 2941 22654 2975
rect 23213 2941 23247 2975
rect 23673 2941 23707 2975
rect 27813 2941 27847 2975
rect 28641 2941 28675 2975
rect 14841 2873 14875 2907
rect 19441 2873 19475 2907
rect 21142 2873 21176 2907
rect 24035 2873 24069 2907
rect 26157 2873 26191 2907
rect 26433 2873 26467 2907
rect 29101 2873 29135 2907
rect 29561 2873 29595 2907
rect 7113 2805 7147 2839
rect 18245 2805 18279 2839
rect 19165 2805 19199 2839
rect 20729 2805 20763 2839
rect 24593 2805 24627 2839
rect 24869 2805 24903 2839
rect 25237 2805 25271 2839
rect 27997 2805 28031 2839
rect 28365 2805 28399 2839
rect 30389 2805 30423 2839
rect 1961 2601 1995 2635
rect 2375 2601 2409 2635
rect 8125 2601 8159 2635
rect 8493 2601 8527 2635
rect 8861 2601 8895 2635
rect 9597 2601 9631 2635
rect 10057 2601 10091 2635
rect 11667 2601 11701 2635
rect 12955 2601 12989 2635
rect 14933 2601 14967 2635
rect 16589 2601 16623 2635
rect 17325 2601 17359 2635
rect 17969 2601 18003 2635
rect 18705 2601 18739 2635
rect 19073 2601 19107 2635
rect 22109 2601 22143 2635
rect 23765 2601 23799 2635
rect 25237 2601 25271 2635
rect 27031 2601 27065 2635
rect 29101 2601 29135 2635
rect 29469 2601 29503 2635
rect 7849 2533 7883 2567
rect 10793 2533 10827 2567
rect 14565 2533 14599 2567
rect 19441 2533 19475 2567
rect 19717 2533 19751 2567
rect 20913 2533 20947 2567
rect 22569 2533 22603 2567
rect 24317 2533 24351 2567
rect 29745 2533 29779 2567
rect 2272 2465 2306 2499
rect 2697 2465 2731 2499
rect 6745 2465 6779 2499
rect 7757 2465 7791 2499
rect 8677 2465 8711 2499
rect 9137 2465 9171 2499
rect 9781 2465 9815 2499
rect 10241 2465 10275 2499
rect 11564 2465 11598 2499
rect 11989 2465 12023 2499
rect 12868 2465 12902 2499
rect 13369 2465 13403 2499
rect 13737 2465 13771 2499
rect 14473 2465 14507 2499
rect 15669 2465 15703 2499
rect 17141 2465 17175 2499
rect 18521 2465 18555 2499
rect 21256 2465 21290 2499
rect 21649 2465 21683 2499
rect 26960 2465 26994 2499
rect 27940 2465 27974 2499
rect 28365 2465 28399 2499
rect 29837 2465 29871 2499
rect 31344 2465 31378 2499
rect 31769 2465 31803 2499
rect 15209 2397 15243 2431
rect 16313 2397 16347 2431
rect 16957 2397 16991 2431
rect 17601 2397 17635 2431
rect 19625 2397 19659 2431
rect 22477 2397 22511 2431
rect 24225 2397 24259 2431
rect 25513 2397 25547 2431
rect 25697 2397 25731 2431
rect 20177 2329 20211 2363
rect 21327 2329 21361 2363
rect 23029 2329 23063 2363
rect 24777 2329 24811 2363
rect 26249 2329 26283 2363
rect 26525 2261 26559 2295
rect 27445 2261 27479 2295
rect 28043 2261 28077 2295
rect 31447 2261 31481 2295
<< metal1 >>
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1581 12971 1639 12977
rect 1581 12968 1593 12971
rect 1544 12940 1593 12968
rect 1544 12928 1550 12940
rect 1581 12937 1593 12940
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 1728 12940 2421 12968
rect 1728 12928 1734 12940
rect 2409 12937 2421 12940
rect 2455 12968 2467 12971
rect 9122 12968 9128 12980
rect 2455 12940 9128 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 9122 12928 9128 12940
rect 9180 12928 9186 12980
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 24280 12767 24338 12773
rect 1443 12736 2084 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2056 12637 2084 12736
rect 24280 12733 24292 12767
rect 24326 12764 24338 12767
rect 24326 12736 24808 12764
rect 24326 12733 24338 12736
rect 24280 12727 24338 12733
rect 2041 12631 2099 12637
rect 2041 12597 2053 12631
rect 2087 12628 2099 12631
rect 2130 12628 2136 12640
rect 2087 12600 2136 12628
rect 2087 12597 2099 12600
rect 2041 12591 2099 12597
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 3786 12588 3792 12640
rect 3844 12628 3850 12640
rect 5810 12628 5816 12640
rect 3844 12600 5816 12628
rect 3844 12588 3850 12600
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 24351 12631 24409 12637
rect 24351 12597 24363 12631
rect 24397 12628 24409 12631
rect 24578 12628 24584 12640
rect 24397 12600 24584 12628
rect 24397 12597 24409 12600
rect 24351 12591 24409 12597
rect 24578 12588 24584 12600
rect 24636 12588 24642 12640
rect 24780 12637 24808 12736
rect 24765 12631 24823 12637
rect 24765 12597 24777 12631
rect 24811 12628 24823 12631
rect 24946 12628 24952 12640
rect 24811 12600 24952 12628
rect 24811 12597 24823 12600
rect 24765 12591 24823 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 35618 12424 35624 12436
rect 35579 12396 35624 12424
rect 35618 12384 35624 12396
rect 35676 12384 35682 12436
rect 1740 12291 1798 12297
rect 1740 12257 1752 12291
rect 1786 12288 1798 12291
rect 2038 12288 2044 12300
rect 1786 12260 2044 12288
rect 1786 12257 1798 12260
rect 1740 12251 1798 12257
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 2752 12291 2810 12297
rect 2752 12257 2764 12291
rect 2798 12288 2810 12291
rect 3142 12288 3148 12300
rect 2798 12260 3148 12288
rect 2798 12257 2810 12260
rect 2752 12251 2810 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 11032 12291 11090 12297
rect 11032 12257 11044 12291
rect 11078 12288 11090 12291
rect 11330 12288 11336 12300
rect 11078 12260 11336 12288
rect 11078 12257 11090 12260
rect 11032 12251 11090 12257
rect 11330 12248 11336 12260
rect 11388 12248 11394 12300
rect 19153 12291 19211 12297
rect 19153 12257 19165 12291
rect 19199 12288 19211 12291
rect 19426 12288 19432 12300
rect 19199 12260 19432 12288
rect 19199 12257 19211 12260
rect 19153 12251 19211 12257
rect 19426 12248 19432 12260
rect 19484 12248 19490 12300
rect 24118 12297 24124 12300
rect 24096 12291 24124 12297
rect 24096 12257 24108 12291
rect 24096 12251 24124 12257
rect 24118 12248 24124 12251
rect 24176 12248 24182 12300
rect 25108 12291 25166 12297
rect 25108 12257 25120 12291
rect 25154 12288 25166 12291
rect 25222 12288 25228 12300
rect 25154 12260 25228 12288
rect 25154 12257 25166 12260
rect 25108 12251 25166 12257
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 34400 12291 34458 12297
rect 34400 12257 34412 12291
rect 34446 12288 34458 12291
rect 34606 12288 34612 12300
rect 34446 12260 34612 12288
rect 34446 12257 34458 12260
rect 34400 12251 34458 12257
rect 34606 12248 34612 12260
rect 34664 12248 34670 12300
rect 35434 12288 35440 12300
rect 35395 12260 35440 12288
rect 35434 12248 35440 12260
rect 35492 12248 35498 12300
rect 29546 12220 29552 12232
rect 29507 12192 29552 12220
rect 29546 12180 29552 12192
rect 29604 12180 29610 12232
rect 1811 12087 1869 12093
rect 1811 12053 1823 12087
rect 1857 12084 1869 12087
rect 2314 12084 2320 12096
rect 1857 12056 2320 12084
rect 1857 12053 1869 12056
rect 1811 12047 1869 12053
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2774 12044 2780 12096
rect 2832 12093 2838 12096
rect 2832 12087 2881 12093
rect 2832 12053 2835 12087
rect 2869 12053 2881 12087
rect 10134 12084 10140 12096
rect 10095 12056 10140 12084
rect 2832 12047 2881 12053
rect 2832 12044 2838 12047
rect 10134 12044 10140 12056
rect 10192 12044 10198 12096
rect 11103 12087 11161 12093
rect 11103 12053 11115 12087
rect 11149 12084 11161 12087
rect 11422 12084 11428 12096
rect 11149 12056 11428 12084
rect 11149 12053 11161 12056
rect 11103 12047 11161 12053
rect 11422 12044 11428 12056
rect 11480 12044 11486 12096
rect 19334 12084 19340 12096
rect 19295 12056 19340 12084
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 24167 12087 24225 12093
rect 24167 12053 24179 12087
rect 24213 12084 24225 12087
rect 24394 12084 24400 12096
rect 24213 12056 24400 12084
rect 24213 12053 24225 12056
rect 24167 12047 24225 12053
rect 24394 12044 24400 12056
rect 24452 12044 24458 12096
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 25179 12087 25237 12093
rect 25179 12084 25191 12087
rect 24912 12056 25191 12084
rect 24912 12044 24918 12056
rect 25179 12053 25191 12056
rect 25225 12053 25237 12087
rect 25179 12047 25237 12053
rect 34146 12044 34152 12096
rect 34204 12084 34210 12096
rect 34471 12087 34529 12093
rect 34471 12084 34483 12087
rect 34204 12056 34483 12084
rect 34204 12044 34210 12056
rect 34471 12053 34483 12056
rect 34517 12053 34529 12087
rect 34471 12047 34529 12053
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 20855 11883 20913 11889
rect 20855 11849 20867 11883
rect 20901 11880 20913 11883
rect 22462 11880 22468 11892
rect 20901 11852 22468 11880
rect 20901 11849 20913 11852
rect 20855 11843 20913 11849
rect 22462 11840 22468 11852
rect 22520 11840 22526 11892
rect 31757 11883 31815 11889
rect 31757 11849 31769 11883
rect 31803 11880 31815 11883
rect 35345 11883 35403 11889
rect 35345 11880 35357 11883
rect 31803 11852 35357 11880
rect 31803 11849 31815 11852
rect 31757 11843 31815 11849
rect 2038 11812 2044 11824
rect 1999 11784 2044 11812
rect 2038 11772 2044 11784
rect 2096 11772 2102 11824
rect 18785 11815 18843 11821
rect 18785 11781 18797 11815
rect 18831 11812 18843 11815
rect 19518 11812 19524 11824
rect 18831 11784 19524 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 19518 11772 19524 11784
rect 19576 11772 19582 11824
rect 2222 11704 2228 11756
rect 2280 11744 2286 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 2280 11716 3341 11744
rect 2280 11704 2286 11716
rect 2608 11685 2636 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 10134 11744 10140 11756
rect 9732 11716 10140 11744
rect 9732 11704 9738 11716
rect 10134 11704 10140 11716
rect 10192 11744 10198 11756
rect 10962 11744 10968 11756
rect 10192 11716 10968 11744
rect 10192 11704 10198 11716
rect 10336 11685 10364 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2568 11679 2636 11685
rect 1443 11648 2452 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 2424 11552 2452 11648
rect 2568 11645 2580 11679
rect 2614 11648 2636 11679
rect 10321 11679 10379 11685
rect 2614 11645 2626 11648
rect 2568 11639 2626 11645
rect 10321 11645 10333 11679
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10597 11679 10655 11685
rect 10597 11645 10609 11679
rect 10643 11645 10655 11679
rect 18598 11676 18604 11688
rect 18559 11648 18604 11676
rect 10597 11639 10655 11645
rect 2406 11540 2412 11552
rect 2367 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 2590 11500 2596 11552
rect 2648 11549 2654 11552
rect 2648 11543 2697 11549
rect 2648 11509 2651 11543
rect 2685 11509 2697 11543
rect 2648 11503 2697 11509
rect 3053 11543 3111 11549
rect 3053 11509 3065 11543
rect 3099 11540 3111 11543
rect 3142 11540 3148 11552
rect 3099 11512 3148 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 2648 11500 2654 11503
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10612 11540 10640 11639
rect 18598 11636 18604 11648
rect 18656 11676 18662 11688
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 18656 11648 19073 11676
rect 18656 11636 18662 11648
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 20784 11679 20842 11685
rect 20784 11645 20796 11679
rect 20830 11676 20842 11679
rect 20830 11648 21312 11676
rect 20830 11645 20842 11648
rect 20784 11639 20842 11645
rect 10778 11608 10784 11620
rect 10739 11580 10784 11608
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 10686 11540 10692 11552
rect 9999 11512 10692 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 11330 11540 11336 11552
rect 11195 11512 11336 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11330 11500 11336 11512
rect 11388 11500 11394 11552
rect 15654 11540 15660 11552
rect 15615 11512 15660 11540
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 19426 11540 19432 11552
rect 19387 11512 19432 11540
rect 19426 11500 19432 11512
rect 19484 11500 19490 11552
rect 19702 11540 19708 11552
rect 19663 11512 19708 11540
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 21284 11549 21312 11648
rect 24302 11636 24308 11688
rect 24360 11676 24366 11688
rect 30098 11685 30104 11688
rect 24432 11679 24490 11685
rect 24432 11676 24444 11679
rect 24360 11648 24444 11676
rect 24360 11636 24366 11648
rect 24432 11645 24444 11648
rect 24478 11676 24490 11679
rect 24857 11679 24915 11685
rect 24857 11676 24869 11679
rect 24478 11648 24869 11676
rect 24478 11645 24490 11648
rect 24432 11639 24490 11645
rect 24857 11645 24869 11648
rect 24903 11645 24915 11679
rect 24857 11639 24915 11645
rect 30076 11679 30104 11685
rect 30076 11645 30088 11679
rect 30156 11676 30162 11688
rect 31272 11679 31330 11685
rect 30156 11648 30604 11676
rect 30076 11639 30104 11645
rect 30098 11636 30104 11639
rect 30156 11636 30162 11648
rect 30576 11617 30604 11648
rect 31272 11645 31284 11679
rect 31318 11676 31330 11679
rect 31772 11676 31800 11843
rect 33428 11824 33456 11852
rect 35345 11849 35357 11852
rect 35391 11880 35403 11883
rect 35434 11880 35440 11892
rect 35391 11852 35440 11880
rect 35391 11849 35403 11852
rect 35345 11843 35403 11849
rect 35434 11840 35440 11852
rect 35492 11840 35498 11892
rect 35621 11883 35679 11889
rect 35621 11849 35633 11883
rect 35667 11880 35679 11883
rect 35710 11880 35716 11892
rect 35667 11852 35716 11880
rect 35667 11849 35679 11852
rect 35621 11843 35679 11849
rect 35710 11840 35716 11852
rect 35768 11840 35774 11892
rect 36679 11883 36737 11889
rect 36679 11849 36691 11883
rect 36725 11880 36737 11883
rect 37182 11880 37188 11892
rect 36725 11852 37188 11880
rect 36725 11849 36737 11852
rect 36679 11843 36737 11849
rect 37182 11840 37188 11852
rect 37240 11840 37246 11892
rect 33410 11772 33416 11824
rect 33468 11772 33474 11824
rect 33870 11685 33876 11688
rect 31318 11648 31800 11676
rect 33848 11679 33876 11685
rect 31318 11645 31330 11648
rect 31272 11639 31330 11645
rect 33848 11645 33860 11679
rect 33928 11676 33934 11688
rect 34241 11679 34299 11685
rect 34241 11676 34253 11679
rect 33928 11648 34253 11676
rect 33848 11639 33876 11645
rect 33870 11636 33876 11639
rect 33928 11636 33934 11648
rect 34241 11645 34253 11648
rect 34287 11645 34299 11679
rect 34241 11639 34299 11645
rect 35342 11636 35348 11688
rect 35400 11676 35406 11688
rect 35437 11679 35495 11685
rect 35437 11676 35449 11679
rect 35400 11648 35449 11676
rect 35400 11636 35406 11648
rect 35437 11645 35449 11648
rect 35483 11676 35495 11679
rect 35989 11679 36047 11685
rect 35989 11676 36001 11679
rect 35483 11648 36001 11676
rect 35483 11645 35495 11648
rect 35437 11639 35495 11645
rect 35989 11645 36001 11648
rect 36035 11645 36047 11679
rect 35989 11639 36047 11645
rect 36538 11636 36544 11688
rect 36596 11685 36602 11688
rect 36596 11679 36634 11685
rect 36622 11676 36634 11679
rect 37001 11679 37059 11685
rect 37001 11676 37013 11679
rect 36622 11648 37013 11676
rect 36622 11645 36634 11648
rect 36596 11639 36634 11645
rect 37001 11645 37013 11648
rect 37047 11645 37059 11679
rect 37001 11639 37059 11645
rect 36596 11636 36602 11639
rect 30561 11611 30619 11617
rect 30561 11577 30573 11611
rect 30607 11608 30619 11611
rect 30607 11580 31616 11608
rect 30607 11577 30619 11580
rect 30561 11571 30619 11577
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21634 11540 21640 11552
rect 21315 11512 21640 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 24118 11540 24124 11552
rect 24079 11512 24124 11540
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24535 11543 24593 11549
rect 24535 11509 24547 11543
rect 24581 11540 24593 11543
rect 24670 11540 24676 11552
rect 24581 11512 24676 11540
rect 24581 11509 24593 11512
rect 24535 11503 24593 11509
rect 24670 11500 24676 11512
rect 24728 11500 24734 11552
rect 25222 11540 25228 11552
rect 25183 11512 25228 11540
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 25406 11540 25412 11552
rect 25367 11512 25412 11540
rect 25406 11500 25412 11512
rect 25464 11500 25470 11552
rect 30147 11543 30205 11549
rect 30147 11509 30159 11543
rect 30193 11540 30205 11543
rect 30282 11540 30288 11552
rect 30193 11512 30288 11540
rect 30193 11509 30205 11512
rect 30147 11503 30205 11509
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 31343 11543 31401 11549
rect 31343 11509 31355 11543
rect 31389 11540 31401 11543
rect 31478 11540 31484 11552
rect 31389 11512 31484 11540
rect 31389 11509 31401 11512
rect 31343 11503 31401 11509
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 31588 11540 31616 11580
rect 32030 11568 32036 11620
rect 32088 11608 32094 11620
rect 34606 11608 34612 11620
rect 32088 11580 34612 11608
rect 32088 11568 32094 11580
rect 34606 11568 34612 11580
rect 34664 11568 34670 11620
rect 33778 11540 33784 11552
rect 31588 11512 33784 11540
rect 33778 11500 33784 11512
rect 33836 11500 33842 11552
rect 33919 11543 33977 11549
rect 33919 11509 33931 11543
rect 33965 11540 33977 11543
rect 34054 11540 34060 11552
rect 33965 11512 34060 11540
rect 33965 11509 33977 11512
rect 33919 11503 33977 11509
rect 34054 11500 34060 11512
rect 34112 11500 34118 11552
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 10134 11336 10140 11348
rect 10095 11308 10140 11336
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 26651 11339 26709 11345
rect 26651 11305 26663 11339
rect 26697 11336 26709 11339
rect 27430 11336 27436 11348
rect 26697 11308 27436 11336
rect 26697 11305 26709 11308
rect 26651 11299 26709 11305
rect 27430 11296 27436 11308
rect 27488 11296 27494 11348
rect 31478 11336 31484 11348
rect 31439 11308 31484 11336
rect 31478 11296 31484 11308
rect 31536 11296 31542 11348
rect 35618 11336 35624 11348
rect 35579 11308 35624 11336
rect 35618 11296 35624 11308
rect 35676 11296 35682 11348
rect 11606 11268 11612 11280
rect 11567 11240 11612 11268
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 20806 11228 20812 11280
rect 20864 11268 20870 11280
rect 21085 11271 21143 11277
rect 21085 11268 21097 11271
rect 20864 11240 21097 11268
rect 20864 11228 20870 11240
rect 21085 11237 21097 11240
rect 21131 11237 21143 11271
rect 24394 11268 24400 11280
rect 24355 11240 24400 11268
rect 21085 11231 21143 11237
rect 24394 11228 24400 11240
rect 24452 11228 24458 11280
rect 24486 11228 24492 11280
rect 24544 11268 24550 11280
rect 24544 11240 24589 11268
rect 24544 11228 24550 11240
rect 29546 11228 29552 11280
rect 29604 11268 29610 11280
rect 29825 11271 29883 11277
rect 29825 11268 29837 11271
rect 29604 11240 29837 11268
rect 29604 11228 29610 11240
rect 29825 11237 29837 11240
rect 29871 11237 29883 11271
rect 29825 11231 29883 11237
rect 29914 11228 29920 11280
rect 29972 11268 29978 11280
rect 30466 11268 30472 11280
rect 29972 11240 30017 11268
rect 30427 11240 30472 11268
rect 29972 11228 29978 11240
rect 30466 11228 30472 11240
rect 30524 11228 30530 11280
rect 33502 11228 33508 11280
rect 33560 11268 33566 11280
rect 33560 11240 36584 11268
rect 33560 11228 33566 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1670 11200 1676 11212
rect 1443 11172 1676 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 2507 11203 2565 11209
rect 2507 11169 2519 11203
rect 2553 11169 2565 11203
rect 2507 11163 2565 11169
rect 4132 11203 4190 11209
rect 4132 11169 4144 11203
rect 4178 11200 4190 11203
rect 4798 11200 4804 11212
rect 4178 11172 4804 11200
rect 4178 11169 4190 11172
rect 4132 11163 4190 11169
rect 2516 11132 2544 11163
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 8570 11200 8576 11212
rect 8531 11172 8576 11200
rect 8570 11160 8576 11172
rect 8628 11160 8634 11212
rect 10042 11200 10048 11212
rect 10003 11172 10048 11200
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10686 11200 10692 11212
rect 10459 11172 10692 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11200 13047 11203
rect 13446 11200 13452 11212
rect 13035 11172 13452 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 13446 11160 13452 11172
rect 13504 11160 13510 11212
rect 15473 11203 15531 11209
rect 15473 11169 15485 11203
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 11514 11132 11520 11144
rect 2516 11104 2728 11132
rect 11475 11104 11520 11132
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 2700 10996 2728 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 15488 11132 15516 11163
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 18230 11209 18236 11212
rect 15933 11203 15991 11209
rect 15933 11200 15945 11203
rect 15620 11172 15945 11200
rect 15620 11160 15626 11172
rect 15933 11169 15945 11172
rect 15979 11169 15991 11203
rect 15933 11163 15991 11169
rect 18208 11203 18236 11209
rect 18208 11169 18220 11203
rect 18208 11163 18236 11169
rect 18230 11160 18236 11163
rect 18288 11160 18294 11212
rect 19334 11200 19340 11212
rect 19295 11172 19340 11200
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 23382 11209 23388 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19576 11172 19625 11200
rect 19576 11160 19582 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 23360 11203 23388 11209
rect 23360 11169 23372 11203
rect 23360 11163 23388 11169
rect 23382 11160 23388 11163
rect 23440 11160 23446 11212
rect 26580 11203 26638 11209
rect 26580 11169 26592 11203
rect 26626 11200 26638 11203
rect 27062 11200 27068 11212
rect 26626 11172 27068 11200
rect 26626 11169 26638 11172
rect 26580 11163 26638 11169
rect 27062 11160 27068 11172
rect 27120 11160 27126 11212
rect 28074 11200 28080 11212
rect 28035 11172 28080 11200
rect 28074 11160 28080 11172
rect 28132 11160 28138 11212
rect 28261 11203 28319 11209
rect 28261 11169 28273 11203
rect 28307 11169 28319 11203
rect 28261 11163 28319 11169
rect 16114 11132 16120 11144
rect 15488 11104 16120 11132
rect 11793 11095 11851 11101
rect 4246 11073 4252 11076
rect 4203 11067 4252 11073
rect 4203 11033 4215 11067
rect 4249 11033 4252 11067
rect 4203 11027 4252 11033
rect 4246 11024 4252 11027
rect 4304 11024 4310 11076
rect 8757 11067 8815 11073
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 10042 11064 10048 11076
rect 8803 11036 10048 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11808 11064 11836 11095
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11132 21051 11135
rect 21450 11132 21456 11144
rect 21039 11104 21456 11132
rect 21039 11101 21051 11104
rect 20993 11095 21051 11101
rect 13170 11064 13176 11076
rect 11204 11036 11836 11064
rect 13131 11036 13176 11064
rect 11204 11024 11210 11036
rect 13170 11024 13176 11036
rect 13228 11024 13234 11076
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 18279 11067 18337 11073
rect 18279 11064 18291 11067
rect 18012 11036 18291 11064
rect 18012 11024 18018 11036
rect 18279 11033 18291 11036
rect 18325 11033 18337 11067
rect 19904 11064 19932 11095
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21634 11132 21640 11144
rect 21595 11104 21640 11132
rect 21634 11092 21640 11104
rect 21692 11092 21698 11144
rect 25038 11132 25044 11144
rect 24999 11104 25044 11132
rect 25038 11092 25044 11104
rect 25096 11092 25102 11144
rect 28276 11132 28304 11163
rect 31754 11160 31760 11212
rect 31812 11200 31818 11212
rect 32125 11203 32183 11209
rect 32125 11200 32137 11203
rect 31812 11172 32137 11200
rect 31812 11160 31818 11172
rect 32125 11169 32137 11172
rect 32171 11169 32183 11203
rect 32125 11163 32183 11169
rect 32398 11160 32404 11212
rect 32456 11200 32462 11212
rect 32585 11203 32643 11209
rect 32585 11200 32597 11203
rect 32456 11172 32597 11200
rect 32456 11160 32462 11172
rect 32585 11169 32597 11172
rect 32631 11169 32643 11203
rect 32585 11163 32643 11169
rect 33962 11160 33968 11212
rect 34020 11200 34026 11212
rect 34333 11203 34391 11209
rect 34333 11200 34345 11203
rect 34020 11172 34345 11200
rect 34020 11160 34026 11172
rect 34333 11169 34345 11172
rect 34379 11169 34391 11203
rect 35434 11200 35440 11212
rect 35395 11172 35440 11200
rect 34333 11163 34391 11169
rect 35434 11160 35440 11172
rect 35492 11200 35498 11212
rect 35894 11200 35900 11212
rect 35492 11172 35900 11200
rect 35492 11160 35498 11172
rect 35894 11160 35900 11172
rect 35952 11160 35958 11212
rect 36556 11209 36584 11240
rect 36541 11203 36599 11209
rect 36541 11169 36553 11203
rect 36587 11200 36599 11203
rect 36998 11200 37004 11212
rect 36587 11172 37004 11200
rect 36587 11169 36599 11172
rect 36541 11163 36599 11169
rect 36998 11160 37004 11172
rect 37056 11160 37062 11212
rect 27632 11104 28304 11132
rect 28537 11135 28595 11141
rect 21266 11064 21272 11076
rect 19904 11036 21272 11064
rect 18279 11027 18337 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 27632 11008 27660 11104
rect 28537 11101 28549 11135
rect 28583 11132 28595 11135
rect 28902 11132 28908 11144
rect 28583 11104 28908 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 28902 11092 28908 11104
rect 28960 11092 28966 11144
rect 32674 11132 32680 11144
rect 32635 11104 32680 11132
rect 32674 11092 32680 11104
rect 32732 11092 32738 11144
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11132 35035 11135
rect 35066 11132 35072 11144
rect 35023 11104 35072 11132
rect 35023 11101 35035 11104
rect 34977 11095 35035 11101
rect 35066 11092 35072 11104
rect 35124 11092 35130 11144
rect 36722 11064 36728 11076
rect 36683 11036 36728 11064
rect 36722 11024 36728 11036
rect 36780 11024 36786 11076
rect 3418 10996 3424 11008
rect 2700 10968 3424 10996
rect 3418 10956 3424 10968
rect 3476 10956 3482 11008
rect 10226 10956 10232 11008
rect 10284 10996 10290 11008
rect 10873 10999 10931 11005
rect 10873 10996 10885 10999
rect 10284 10968 10885 10996
rect 10284 10956 10290 10968
rect 10873 10965 10885 10968
rect 10919 10965 10931 10999
rect 10873 10959 10931 10965
rect 12529 10999 12587 11005
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12710 10996 12716 11008
rect 12575 10968 12716 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 20162 10996 20168 11008
rect 20123 10968 20168 10996
rect 20162 10956 20168 10968
rect 20220 10956 20226 11008
rect 23198 10956 23204 11008
rect 23256 10996 23262 11008
rect 23431 10999 23489 11005
rect 23431 10996 23443 10999
rect 23256 10968 23443 10996
rect 23256 10956 23262 10968
rect 23431 10965 23443 10968
rect 23477 10965 23489 10999
rect 27614 10996 27620 11008
rect 27575 10968 27620 10996
rect 23431 10959 23489 10965
rect 27614 10956 27620 10968
rect 27672 10956 27678 11008
rect 34517 10999 34575 11005
rect 34517 10965 34529 10999
rect 34563 10996 34575 10999
rect 34790 10996 34796 11008
rect 34563 10968 34796 10996
rect 34563 10965 34575 10968
rect 34517 10959 34575 10965
rect 34790 10956 34796 10968
rect 34848 10956 34854 11008
rect 34974 10956 34980 11008
rect 35032 10996 35038 11008
rect 35253 10999 35311 11005
rect 35253 10996 35265 10999
rect 35032 10968 35265 10996
rect 35032 10956 35038 10968
rect 35253 10965 35265 10968
rect 35299 10965 35311 10999
rect 35253 10959 35311 10965
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 4798 10792 4804 10804
rect 4759 10764 4804 10792
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8628 10764 8953 10792
rect 8628 10752 8634 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 11517 10795 11575 10801
rect 11517 10761 11529 10795
rect 11563 10792 11575 10795
rect 11606 10792 11612 10804
rect 11563 10764 11612 10792
rect 11563 10761 11575 10764
rect 11517 10755 11575 10761
rect 11606 10752 11612 10764
rect 11664 10752 11670 10804
rect 16715 10795 16773 10801
rect 16715 10761 16727 10795
rect 16761 10792 16773 10795
rect 17494 10792 17500 10804
rect 16761 10764 17500 10792
rect 16761 10761 16773 10764
rect 16715 10755 16773 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19392 10764 19809 10792
rect 19392 10752 19398 10764
rect 19797 10761 19809 10764
rect 19843 10792 19855 10795
rect 21358 10792 21364 10804
rect 19843 10764 21364 10792
rect 19843 10761 19855 10764
rect 19797 10755 19855 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 21726 10792 21732 10804
rect 21687 10764 21732 10792
rect 21726 10752 21732 10764
rect 21784 10752 21790 10804
rect 23106 10792 23112 10804
rect 23067 10764 23112 10792
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 24029 10795 24087 10801
rect 24029 10761 24041 10795
rect 24075 10792 24087 10795
rect 24394 10792 24400 10804
rect 24075 10764 24400 10792
rect 24075 10761 24087 10764
rect 24029 10755 24087 10761
rect 24394 10752 24400 10764
rect 24452 10752 24458 10804
rect 27062 10792 27068 10804
rect 27023 10764 27068 10792
rect 27062 10752 27068 10764
rect 27120 10752 27126 10804
rect 29546 10752 29552 10804
rect 29604 10792 29610 10804
rect 29733 10795 29791 10801
rect 29733 10792 29745 10795
rect 29604 10764 29745 10792
rect 29604 10752 29610 10764
rect 29733 10761 29745 10764
rect 29779 10761 29791 10795
rect 29733 10755 29791 10761
rect 33226 10752 33232 10804
rect 33284 10792 33290 10804
rect 33962 10792 33968 10804
rect 33284 10764 33968 10792
rect 33284 10752 33290 10764
rect 33962 10752 33968 10764
rect 34020 10792 34026 10804
rect 34333 10795 34391 10801
rect 34333 10792 34345 10795
rect 34020 10764 34345 10792
rect 34020 10752 34026 10764
rect 34333 10761 34345 10764
rect 34379 10761 34391 10795
rect 35894 10792 35900 10804
rect 35855 10764 35900 10792
rect 34333 10755 34391 10761
rect 35894 10752 35900 10764
rect 35952 10752 35958 10804
rect 36630 10792 36636 10804
rect 36591 10764 36636 10792
rect 36630 10752 36636 10764
rect 36688 10752 36694 10804
rect 36998 10792 37004 10804
rect 36959 10764 37004 10792
rect 36998 10752 37004 10764
rect 37056 10752 37062 10804
rect 8297 10727 8355 10733
rect 8297 10693 8309 10727
rect 8343 10724 8355 10727
rect 9582 10724 9588 10736
rect 8343 10696 9588 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 9582 10684 9588 10696
rect 9640 10684 9646 10736
rect 29089 10727 29147 10733
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 29454 10724 29460 10736
rect 29135 10696 29460 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 29454 10684 29460 10696
rect 29512 10724 29518 10736
rect 29914 10724 29920 10736
rect 29512 10696 29920 10724
rect 29512 10684 29518 10696
rect 29914 10684 29920 10696
rect 29972 10684 29978 10736
rect 31478 10684 31484 10736
rect 31536 10684 31542 10736
rect 34054 10684 34060 10736
rect 34112 10724 34118 10736
rect 36265 10727 36323 10733
rect 36265 10724 36277 10727
rect 34112 10696 36277 10724
rect 34112 10684 34118 10696
rect 36265 10693 36277 10696
rect 36311 10693 36323 10727
rect 36265 10687 36323 10693
rect 9263 10659 9321 10665
rect 9263 10625 9275 10659
rect 9309 10656 9321 10659
rect 11514 10656 11520 10668
rect 9309 10628 11520 10656
rect 9309 10625 9321 10628
rect 9263 10619 9321 10625
rect 11514 10616 11520 10628
rect 11572 10656 11578 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 11572 10628 11805 10656
rect 11572 10616 11578 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 14918 10616 14924 10668
rect 14976 10656 14982 10668
rect 15381 10659 15439 10665
rect 15381 10656 15393 10659
rect 14976 10628 15393 10656
rect 14976 10616 14982 10628
rect 15381 10625 15393 10628
rect 15427 10656 15439 10659
rect 16206 10656 16212 10668
rect 15427 10628 16212 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 19702 10616 19708 10668
rect 19760 10656 19766 10668
rect 20070 10656 20076 10668
rect 19760 10628 20076 10656
rect 19760 10616 19766 10628
rect 20070 10616 20076 10628
rect 20128 10616 20134 10668
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10656 20775 10659
rect 21634 10656 21640 10668
rect 20763 10628 21640 10656
rect 20763 10625 20775 10628
rect 20717 10619 20775 10625
rect 21634 10616 21640 10628
rect 21692 10616 21698 10668
rect 24578 10656 24584 10668
rect 24539 10628 24584 10656
rect 24578 10616 24584 10628
rect 24636 10656 24642 10668
rect 25501 10659 25559 10665
rect 25501 10656 25513 10659
rect 24636 10628 25513 10656
rect 24636 10616 24642 10628
rect 25501 10625 25513 10628
rect 25547 10625 25559 10659
rect 29270 10656 29276 10668
rect 25501 10619 25559 10625
rect 26068 10628 29276 10656
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2056 10464 2084 10560
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2568 10591 2626 10597
rect 2568 10588 2580 10591
rect 2188 10560 2580 10588
rect 2188 10548 2194 10560
rect 2568 10557 2580 10560
rect 2614 10557 2626 10591
rect 3050 10588 3056 10600
rect 3011 10560 3056 10588
rect 2568 10551 2626 10557
rect 2583 10520 2611 10551
rect 3050 10548 3056 10560
rect 3108 10548 3114 10600
rect 3948 10591 4006 10597
rect 3948 10557 3960 10591
rect 3994 10588 4006 10591
rect 8113 10591 8171 10597
rect 3994 10560 4476 10588
rect 3994 10557 4006 10560
rect 3948 10551 4006 10557
rect 3068 10520 3096 10548
rect 2583 10492 3096 10520
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2682 10461 2688 10464
rect 2639 10455 2688 10461
rect 2639 10421 2651 10455
rect 2685 10421 2688 10455
rect 2639 10415 2688 10421
rect 2682 10412 2688 10415
rect 2740 10412 2746 10464
rect 3418 10452 3424 10464
rect 3379 10424 3424 10452
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4062 10461 4068 10464
rect 4019 10455 4068 10461
rect 4019 10421 4031 10455
rect 4065 10421 4068 10455
rect 4019 10415 4068 10421
rect 4062 10412 4068 10415
rect 4120 10412 4126 10464
rect 4448 10461 4476 10560
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8159 10560 8585 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 9122 10588 9128 10600
rect 9086 10560 9128 10588
rect 8573 10551 8631 10557
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4706 10452 4712 10464
rect 4479 10424 4712 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6604 10424 6837 10452
rect 6604 10412 6610 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 8588 10452 8616 10551
rect 9122 10548 9128 10560
rect 9180 10597 9186 10600
rect 9180 10591 9234 10597
rect 9180 10557 9188 10591
rect 9222 10588 9234 10591
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9222 10560 9689 10588
rect 9222 10557 9234 10560
rect 9180 10551 9234 10557
rect 9677 10557 9689 10560
rect 9723 10588 9735 10591
rect 9950 10588 9956 10600
rect 9723 10560 9956 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 9180 10548 9186 10551
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 12710 10588 12716 10600
rect 12671 10560 12716 10588
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 14182 10588 14188 10600
rect 13035 10560 14188 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 10226 10520 10232 10532
rect 10187 10492 10232 10520
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10873 10523 10931 10529
rect 10376 10492 10421 10520
rect 10376 10480 10382 10492
rect 10873 10489 10885 10523
rect 10919 10520 10931 10523
rect 11146 10520 11152 10532
rect 10919 10492 11152 10520
rect 10919 10489 10931 10492
rect 10873 10483 10931 10489
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 13004 10520 13032 10551
rect 14182 10548 14188 10560
rect 14240 10548 14246 10600
rect 16224 10588 16252 10616
rect 16612 10591 16670 10597
rect 16612 10588 16624 10591
rect 16224 10560 16624 10588
rect 16612 10557 16624 10560
rect 16658 10588 16670 10591
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 16658 10560 17049 10588
rect 16658 10557 16670 10560
rect 16612 10551 16670 10557
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 17678 10548 17684 10600
rect 17736 10588 17742 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17736 10560 17877 10588
rect 17736 10548 17742 10560
rect 17865 10557 17877 10560
rect 17911 10588 17923 10591
rect 18417 10591 18475 10597
rect 18417 10588 18429 10591
rect 17911 10560 18429 10588
rect 17911 10557 17923 10560
rect 17865 10551 17923 10557
rect 18417 10557 18429 10560
rect 18463 10557 18475 10591
rect 18417 10551 18475 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10557 19027 10591
rect 21542 10588 21548 10600
rect 21503 10560 21548 10588
rect 18969 10551 19027 10557
rect 15102 10520 15108 10532
rect 12176 10492 13032 10520
rect 15063 10492 15108 10520
rect 9214 10452 9220 10464
rect 8588 10424 9220 10452
rect 6825 10415 6883 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10452 10103 10455
rect 10686 10452 10692 10464
rect 10091 10424 10692 10452
rect 10091 10421 10103 10424
rect 10045 10415 10103 10421
rect 10686 10412 10692 10424
rect 10744 10452 10750 10464
rect 12176 10461 12204 10492
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 15194 10480 15200 10532
rect 15252 10520 15258 10532
rect 16114 10520 16120 10532
rect 15252 10492 15297 10520
rect 16027 10492 16120 10520
rect 15252 10480 15258 10492
rect 16114 10480 16120 10492
rect 16172 10520 16178 10532
rect 17696 10520 17724 10548
rect 16172 10492 17724 10520
rect 16172 10480 16178 10492
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 10744 10424 12173 10452
rect 10744 10412 10750 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 12342 10412 12348 10464
rect 12400 10452 12406 10464
rect 12529 10455 12587 10461
rect 12529 10452 12541 10455
rect 12400 10424 12541 10452
rect 12400 10412 12406 10424
rect 12529 10421 12541 10424
rect 12575 10421 12587 10455
rect 13446 10452 13452 10464
rect 13407 10424 13452 10452
rect 12529 10415 12587 10421
rect 13446 10412 13452 10424
rect 13504 10412 13510 10464
rect 14001 10455 14059 10461
rect 14001 10421 14013 10455
rect 14047 10452 14059 10455
rect 14826 10452 14832 10464
rect 14047 10424 14832 10452
rect 14047 10421 14059 10424
rect 14001 10415 14059 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14921 10455 14979 10461
rect 14921 10421 14933 10455
rect 14967 10452 14979 10455
rect 15212 10452 15240 10480
rect 18230 10452 18236 10464
rect 14967 10424 15240 10452
rect 18191 10424 18236 10452
rect 14967 10421 14979 10424
rect 14921 10415 14979 10421
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 18984 10452 19012 10551
rect 21542 10548 21548 10560
rect 21600 10588 21606 10600
rect 22005 10591 22063 10597
rect 22005 10588 22017 10591
rect 21600 10560 22017 10588
rect 21600 10548 21606 10560
rect 22005 10557 22017 10560
rect 22051 10557 22063 10591
rect 22005 10551 22063 10557
rect 22186 10548 22192 10600
rect 22244 10588 22250 10600
rect 22624 10591 22682 10597
rect 22624 10588 22636 10591
rect 22244 10560 22636 10588
rect 22244 10548 22250 10560
rect 22624 10557 22636 10560
rect 22670 10588 22682 10591
rect 23106 10588 23112 10600
rect 22670 10560 23112 10588
rect 22670 10557 22682 10560
rect 22624 10551 22682 10557
rect 23106 10548 23112 10560
rect 23164 10548 23170 10600
rect 25958 10588 25964 10600
rect 25871 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10588 26022 10600
rect 26068 10597 26096 10628
rect 26053 10591 26111 10597
rect 26053 10588 26065 10591
rect 26016 10560 26065 10588
rect 26016 10548 26022 10560
rect 26053 10557 26065 10560
rect 26099 10557 26111 10591
rect 26053 10551 26111 10557
rect 26142 10548 26148 10600
rect 26200 10588 26206 10600
rect 27632 10597 27660 10628
rect 29270 10616 29276 10628
rect 29328 10616 29334 10668
rect 30466 10656 30472 10668
rect 30427 10628 30472 10656
rect 30466 10616 30472 10628
rect 30524 10616 30530 10668
rect 31496 10656 31524 10684
rect 31573 10659 31631 10665
rect 31573 10656 31585 10659
rect 31496 10628 31585 10656
rect 31573 10625 31585 10628
rect 31619 10625 31631 10659
rect 31573 10619 31631 10625
rect 32398 10616 32404 10668
rect 32456 10656 32462 10668
rect 32456 10628 33548 10656
rect 32456 10616 32462 10628
rect 26513 10591 26571 10597
rect 26513 10588 26525 10591
rect 26200 10560 26525 10588
rect 26200 10548 26206 10560
rect 26513 10557 26525 10560
rect 26559 10557 26571 10591
rect 26513 10551 26571 10557
rect 27525 10591 27583 10597
rect 27525 10557 27537 10591
rect 27571 10588 27583 10591
rect 27617 10591 27675 10597
rect 27617 10588 27629 10591
rect 27571 10560 27629 10588
rect 27571 10557 27583 10560
rect 27525 10551 27583 10557
rect 27617 10557 27629 10560
rect 27663 10557 27675 10591
rect 27617 10551 27675 10557
rect 27706 10548 27712 10600
rect 27764 10588 27770 10600
rect 27982 10588 27988 10600
rect 27764 10560 27988 10588
rect 27764 10548 27770 10560
rect 27982 10548 27988 10560
rect 28040 10588 28046 10600
rect 33520 10597 33548 10628
rect 28077 10591 28135 10597
rect 28077 10588 28089 10591
rect 28040 10560 28089 10588
rect 28040 10548 28046 10560
rect 28077 10557 28089 10560
rect 28123 10557 28135 10591
rect 33045 10591 33103 10597
rect 33045 10588 33057 10591
rect 28077 10551 28135 10557
rect 32876 10560 33057 10588
rect 19150 10520 19156 10532
rect 19111 10492 19156 10520
rect 19150 10480 19156 10492
rect 19208 10480 19214 10532
rect 20162 10480 20168 10532
rect 20220 10520 20226 10532
rect 20220 10492 20265 10520
rect 20220 10480 20226 10492
rect 24578 10480 24584 10532
rect 24636 10520 24642 10532
rect 24673 10523 24731 10529
rect 24673 10520 24685 10523
rect 24636 10492 24685 10520
rect 24636 10480 24642 10492
rect 24673 10489 24685 10492
rect 24719 10489 24731 10523
rect 24673 10483 24731 10489
rect 25038 10480 25044 10532
rect 25096 10520 25102 10532
rect 25225 10523 25283 10529
rect 25225 10520 25237 10523
rect 25096 10492 25237 10520
rect 25096 10480 25102 10492
rect 25225 10489 25237 10492
rect 25271 10489 25283 10523
rect 28350 10520 28356 10532
rect 28311 10492 28356 10520
rect 25225 10483 25283 10489
rect 28350 10480 28356 10492
rect 28408 10480 28414 10532
rect 30009 10523 30067 10529
rect 30009 10489 30021 10523
rect 30055 10489 30067 10523
rect 30009 10483 30067 10489
rect 19518 10452 19524 10464
rect 18984 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 20806 10412 20812 10464
rect 20864 10452 20870 10464
rect 20993 10455 21051 10461
rect 20993 10452 21005 10455
rect 20864 10424 21005 10452
rect 20864 10412 20870 10424
rect 20993 10421 21005 10424
rect 21039 10421 21051 10455
rect 21450 10452 21456 10464
rect 21411 10424 21456 10452
rect 20993 10415 21051 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 22695 10455 22753 10461
rect 22695 10421 22707 10455
rect 22741 10452 22753 10455
rect 22922 10452 22928 10464
rect 22741 10424 22928 10452
rect 22741 10421 22753 10424
rect 22695 10415 22753 10421
rect 22922 10412 22928 10424
rect 22980 10412 22986 10464
rect 23477 10455 23535 10461
rect 23477 10421 23489 10455
rect 23523 10452 23535 10455
rect 23566 10452 23572 10464
rect 23523 10424 23572 10452
rect 23523 10421 23535 10424
rect 23477 10415 23535 10421
rect 23566 10412 23572 10424
rect 23624 10412 23630 10464
rect 24394 10452 24400 10464
rect 24355 10424 24400 10452
rect 24394 10412 24400 10424
rect 24452 10412 24458 10464
rect 26234 10412 26240 10464
rect 26292 10452 26298 10464
rect 26329 10455 26387 10461
rect 26329 10452 26341 10455
rect 26292 10424 26341 10452
rect 26292 10412 26298 10424
rect 26329 10421 26341 10424
rect 26375 10421 26387 10455
rect 26329 10415 26387 10421
rect 28074 10412 28080 10464
rect 28132 10452 28138 10464
rect 28629 10455 28687 10461
rect 28629 10452 28641 10455
rect 28132 10424 28641 10452
rect 28132 10412 28138 10424
rect 28629 10421 28641 10424
rect 28675 10421 28687 10455
rect 30024 10452 30052 10483
rect 30098 10480 30104 10532
rect 30156 10520 30162 10532
rect 30156 10492 30201 10520
rect 30156 10480 30162 10492
rect 30466 10480 30472 10532
rect 30524 10520 30530 10532
rect 31297 10523 31355 10529
rect 31297 10520 31309 10523
rect 30524 10492 31309 10520
rect 30524 10480 30530 10492
rect 31297 10489 31309 10492
rect 31343 10489 31355 10523
rect 31297 10483 31355 10489
rect 31021 10455 31079 10461
rect 31021 10452 31033 10455
rect 30024 10424 31033 10452
rect 28629 10415 28687 10421
rect 31021 10421 31033 10424
rect 31067 10452 31079 10455
rect 31110 10452 31116 10464
rect 31067 10424 31116 10452
rect 31067 10421 31079 10424
rect 31021 10415 31079 10421
rect 31110 10412 31116 10424
rect 31168 10412 31174 10464
rect 31312 10452 31340 10483
rect 31570 10480 31576 10532
rect 31628 10520 31634 10532
rect 31665 10523 31723 10529
rect 31665 10520 31677 10523
rect 31628 10492 31677 10520
rect 31628 10480 31634 10492
rect 31665 10489 31677 10492
rect 31711 10489 31723 10523
rect 32214 10520 32220 10532
rect 32175 10492 32220 10520
rect 31665 10483 31723 10489
rect 32214 10480 32220 10492
rect 32272 10480 32278 10532
rect 32876 10464 32904 10560
rect 33045 10557 33057 10560
rect 33091 10557 33103 10591
rect 33045 10551 33103 10557
rect 33505 10591 33563 10597
rect 33505 10557 33517 10591
rect 33551 10557 33563 10591
rect 36280 10588 36308 10687
rect 36449 10591 36507 10597
rect 36449 10588 36461 10591
rect 36280 10560 36461 10588
rect 33505 10551 33563 10557
rect 36449 10557 36461 10560
rect 36495 10557 36507 10591
rect 37588 10591 37646 10597
rect 37588 10588 37600 10591
rect 36449 10551 36507 10557
rect 36740 10560 37600 10588
rect 33781 10523 33839 10529
rect 33781 10489 33793 10523
rect 33827 10520 33839 10523
rect 34054 10520 34060 10532
rect 33827 10492 34060 10520
rect 33827 10489 33839 10492
rect 33781 10483 33839 10489
rect 34054 10480 34060 10492
rect 34112 10480 34118 10532
rect 34974 10520 34980 10532
rect 34935 10492 34980 10520
rect 34974 10480 34980 10492
rect 35032 10480 35038 10532
rect 35066 10480 35072 10532
rect 35124 10520 35130 10532
rect 35621 10523 35679 10529
rect 35124 10492 35169 10520
rect 35124 10480 35130 10492
rect 35621 10489 35633 10523
rect 35667 10520 35679 10523
rect 35802 10520 35808 10532
rect 35667 10492 35808 10520
rect 35667 10489 35679 10492
rect 35621 10483 35679 10489
rect 35802 10480 35808 10492
rect 35860 10480 35866 10532
rect 31754 10452 31760 10464
rect 31312 10424 31760 10452
rect 31754 10412 31760 10424
rect 31812 10412 31818 10464
rect 32398 10412 32404 10464
rect 32456 10452 32462 10464
rect 32493 10455 32551 10461
rect 32493 10452 32505 10455
rect 32456 10424 32505 10452
rect 32456 10412 32462 10424
rect 32493 10421 32505 10424
rect 32539 10421 32551 10455
rect 32858 10452 32864 10464
rect 32819 10424 32864 10452
rect 32493 10415 32551 10421
rect 32858 10412 32864 10424
rect 32916 10412 32922 10464
rect 36078 10412 36084 10464
rect 36136 10452 36142 10464
rect 36740 10452 36768 10560
rect 37588 10557 37600 10560
rect 37634 10588 37646 10591
rect 38013 10591 38071 10597
rect 38013 10588 38025 10591
rect 37634 10560 38025 10588
rect 37634 10557 37646 10560
rect 37588 10551 37646 10557
rect 38013 10557 38025 10560
rect 38059 10557 38071 10591
rect 38013 10551 38071 10557
rect 36136 10424 36768 10452
rect 36136 10412 36142 10424
rect 37274 10412 37280 10464
rect 37332 10452 37338 10464
rect 37691 10455 37749 10461
rect 37691 10452 37703 10455
rect 37332 10424 37703 10452
rect 37332 10412 37338 10424
rect 37691 10421 37703 10424
rect 37737 10421 37749 10455
rect 37691 10415 37749 10421
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 1820 10220 2053 10248
rect 1820 10208 1826 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 2041 10211 2099 10217
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4939 10251 4997 10257
rect 4939 10248 4951 10251
rect 4212 10220 4951 10248
rect 4212 10208 4218 10220
rect 4939 10217 4951 10220
rect 4985 10217 4997 10251
rect 4939 10211 4997 10217
rect 9953 10251 10011 10257
rect 9953 10217 9965 10251
rect 9999 10248 10011 10251
rect 10042 10248 10048 10260
rect 9999 10220 10048 10248
rect 9999 10217 10011 10220
rect 9953 10211 10011 10217
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 10318 10208 10324 10220
rect 10376 10248 10382 10260
rect 10962 10248 10968 10260
rect 10376 10220 10968 10248
rect 10376 10208 10382 10220
rect 10962 10208 10968 10220
rect 11020 10208 11026 10260
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 13078 10248 13084 10260
rect 11664 10220 12204 10248
rect 11664 10208 11670 10220
rect 10594 10180 10600 10192
rect 10555 10152 10600 10180
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 12176 10189 12204 10220
rect 12728 10220 13084 10248
rect 12728 10189 12756 10220
rect 13078 10208 13084 10220
rect 13136 10248 13142 10260
rect 15102 10248 15108 10260
rect 13136 10220 15108 10248
rect 13136 10208 13142 10220
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15562 10248 15568 10260
rect 15523 10220 15568 10248
rect 15562 10208 15568 10220
rect 15620 10208 15626 10260
rect 19061 10251 19119 10257
rect 19061 10217 19073 10251
rect 19107 10248 19119 10251
rect 19150 10248 19156 10260
rect 19107 10220 19156 10248
rect 19107 10217 19119 10220
rect 19061 10211 19119 10217
rect 19150 10208 19156 10220
rect 19208 10208 19214 10260
rect 19426 10248 19432 10260
rect 19387 10220 19432 10248
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 20070 10208 20076 10260
rect 20128 10248 20134 10260
rect 20165 10251 20223 10257
rect 20165 10248 20177 10251
rect 20128 10220 20177 10248
rect 20128 10208 20134 10220
rect 20165 10217 20177 10220
rect 20211 10217 20223 10251
rect 26142 10248 26148 10260
rect 26103 10220 26148 10248
rect 20165 10211 20223 10217
rect 26142 10208 26148 10220
rect 26200 10208 26206 10260
rect 26510 10208 26516 10260
rect 26568 10248 26574 10260
rect 27893 10251 27951 10257
rect 26568 10220 26740 10248
rect 26568 10208 26574 10220
rect 12069 10183 12127 10189
rect 12069 10180 12081 10183
rect 11480 10152 12081 10180
rect 11480 10140 11486 10152
rect 12069 10149 12081 10152
rect 12115 10149 12127 10183
rect 12069 10143 12127 10149
rect 12161 10183 12219 10189
rect 12161 10149 12173 10183
rect 12207 10149 12219 10183
rect 12161 10143 12219 10149
rect 12713 10183 12771 10189
rect 12713 10149 12725 10183
rect 12759 10149 12771 10183
rect 12713 10143 12771 10149
rect 2130 10112 2136 10124
rect 2091 10084 2136 10112
rect 2130 10072 2136 10084
rect 2188 10072 2194 10124
rect 2406 10112 2412 10124
rect 2367 10084 2412 10112
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 4868 10115 4926 10121
rect 4868 10081 4880 10115
rect 4914 10112 4926 10115
rect 5166 10112 5172 10124
rect 4914 10084 5172 10112
rect 4914 10081 4926 10084
rect 4868 10075 4926 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 7374 10072 7380 10124
rect 7432 10112 7438 10124
rect 7596 10115 7654 10121
rect 7596 10112 7608 10115
rect 7432 10084 7608 10112
rect 7432 10072 7438 10084
rect 7596 10081 7608 10084
rect 7642 10081 7654 10115
rect 7596 10075 7654 10081
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8608 10115 8666 10121
rect 8608 10112 8620 10115
rect 8444 10084 8620 10112
rect 8444 10072 8450 10084
rect 8608 10081 8620 10084
rect 8654 10081 8666 10115
rect 8608 10075 8666 10081
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10081 13967 10115
rect 14182 10112 14188 10124
rect 14095 10084 14188 10112
rect 13909 10075 13967 10081
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6730 10044 6736 10056
rect 6595 10016 6736 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 10502 10044 10508 10056
rect 10463 10016 10508 10044
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 13924 10044 13952 10075
rect 14182 10072 14188 10084
rect 14240 10112 14246 10124
rect 15580 10112 15608 10208
rect 15654 10140 15660 10192
rect 15712 10180 15718 10192
rect 15933 10183 15991 10189
rect 15933 10180 15945 10183
rect 15712 10152 15945 10180
rect 15712 10140 15718 10152
rect 15933 10149 15945 10152
rect 15979 10149 15991 10183
rect 15933 10143 15991 10149
rect 16025 10183 16083 10189
rect 16025 10149 16037 10183
rect 16071 10180 16083 10183
rect 16574 10180 16580 10192
rect 16071 10152 16580 10180
rect 16071 10149 16083 10152
rect 16025 10143 16083 10149
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 18693 10183 18751 10189
rect 18693 10149 18705 10183
rect 18739 10180 18751 10183
rect 21085 10183 21143 10189
rect 18739 10152 19564 10180
rect 18739 10149 18751 10152
rect 18693 10143 18751 10149
rect 19536 10124 19564 10152
rect 21085 10149 21097 10183
rect 21131 10180 21143 10183
rect 21910 10180 21916 10192
rect 21131 10152 21916 10180
rect 21131 10149 21143 10152
rect 21085 10143 21143 10149
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 23198 10180 23204 10192
rect 23159 10152 23204 10180
rect 23198 10140 23204 10152
rect 23256 10140 23262 10192
rect 23290 10140 23296 10192
rect 23348 10180 23354 10192
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 23348 10152 24501 10180
rect 23348 10140 23354 10152
rect 24489 10149 24501 10152
rect 24535 10180 24547 10183
rect 24578 10180 24584 10192
rect 24535 10152 24584 10180
rect 24535 10149 24547 10152
rect 24489 10143 24547 10149
rect 24578 10140 24584 10152
rect 24636 10140 24642 10192
rect 24762 10180 24768 10192
rect 24723 10152 24768 10180
rect 24762 10140 24768 10152
rect 24820 10140 24826 10192
rect 24857 10183 24915 10189
rect 24857 10149 24869 10183
rect 24903 10180 24915 10183
rect 24946 10180 24952 10192
rect 24903 10152 24952 10180
rect 24903 10149 24915 10152
rect 24857 10143 24915 10149
rect 24946 10140 24952 10152
rect 25004 10140 25010 10192
rect 26602 10180 26608 10192
rect 26563 10152 26608 10180
rect 26602 10140 26608 10152
rect 26660 10140 26666 10192
rect 26712 10189 26740 10220
rect 27893 10217 27905 10251
rect 27939 10248 27951 10251
rect 27982 10248 27988 10260
rect 27939 10220 27988 10248
rect 27939 10217 27951 10220
rect 27893 10211 27951 10217
rect 27982 10208 27988 10220
rect 28040 10208 28046 10260
rect 29454 10248 29460 10260
rect 29415 10220 29460 10248
rect 29454 10208 29460 10220
rect 29512 10208 29518 10260
rect 30374 10208 30380 10260
rect 30432 10248 30438 10260
rect 31570 10248 31576 10260
rect 30432 10220 30512 10248
rect 30432 10208 30438 10220
rect 26697 10183 26755 10189
rect 26697 10149 26709 10183
rect 26743 10149 26755 10183
rect 26697 10143 26755 10149
rect 28810 10140 28816 10192
rect 28868 10189 28874 10192
rect 28868 10183 28916 10189
rect 28868 10149 28870 10183
rect 28904 10149 28916 10183
rect 28868 10143 28916 10149
rect 28868 10140 28874 10143
rect 28994 10140 29000 10192
rect 29052 10180 29058 10192
rect 30484 10189 30512 10220
rect 30576 10220 31576 10248
rect 30576 10192 30604 10220
rect 31570 10208 31576 10220
rect 31628 10208 31634 10260
rect 32674 10248 32680 10260
rect 32635 10220 32680 10248
rect 32674 10208 32680 10220
rect 32732 10208 32738 10260
rect 34057 10251 34115 10257
rect 34057 10217 34069 10251
rect 34103 10248 34115 10251
rect 35802 10248 35808 10260
rect 34103 10220 35808 10248
rect 34103 10217 34115 10220
rect 34057 10211 34115 10217
rect 29733 10183 29791 10189
rect 29733 10180 29745 10183
rect 29052 10152 29745 10180
rect 29052 10140 29058 10152
rect 29733 10149 29745 10152
rect 29779 10149 29791 10183
rect 29733 10143 29791 10149
rect 30469 10183 30527 10189
rect 30469 10149 30481 10183
rect 30515 10149 30527 10183
rect 30469 10143 30527 10149
rect 30558 10140 30564 10192
rect 30616 10180 30622 10192
rect 33134 10180 33140 10192
rect 30616 10152 30709 10180
rect 33095 10152 33140 10180
rect 30616 10140 30622 10152
rect 33134 10140 33140 10152
rect 33192 10140 33198 10192
rect 33686 10180 33692 10192
rect 33647 10152 33692 10180
rect 33686 10140 33692 10152
rect 33744 10140 33750 10192
rect 17586 10112 17592 10124
rect 14240 10084 15608 10112
rect 17547 10084 17592 10112
rect 14240 10072 14246 10084
rect 17586 10072 17592 10084
rect 17644 10072 17650 10124
rect 17862 10072 17868 10124
rect 17920 10112 17926 10124
rect 18141 10115 18199 10121
rect 18141 10112 18153 10115
rect 17920 10084 18153 10112
rect 17920 10072 17926 10084
rect 18141 10081 18153 10084
rect 18187 10112 18199 10115
rect 19334 10112 19340 10124
rect 18187 10084 18460 10112
rect 19295 10084 19340 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 14090 10044 14096 10056
rect 13924 10016 14096 10044
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 16206 10044 16212 10056
rect 16167 10016 16212 10044
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 18322 10044 18328 10056
rect 18283 10016 18328 10044
rect 18322 10004 18328 10016
rect 18380 10004 18386 10056
rect 18432 10044 18460 10084
rect 19334 10072 19340 10084
rect 19392 10072 19398 10124
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 19705 10115 19763 10121
rect 19705 10112 19717 10115
rect 19576 10084 19717 10112
rect 19576 10072 19582 10084
rect 19705 10081 19717 10084
rect 19751 10112 19763 10115
rect 19978 10112 19984 10124
rect 19751 10084 19984 10112
rect 19751 10081 19763 10084
rect 19705 10075 19763 10081
rect 19978 10072 19984 10084
rect 20036 10072 20042 10124
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 21692 10084 21737 10112
rect 21692 10072 21698 10084
rect 19242 10044 19248 10056
rect 18432 10016 19248 10044
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20990 10044 20996 10056
rect 20772 10016 20996 10044
rect 20772 10004 20778 10016
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 23474 10044 23480 10056
rect 23435 10016 23480 10044
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 25038 10044 25044 10056
rect 24999 10016 25044 10044
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 26878 10044 26884 10056
rect 26839 10016 26884 10044
rect 26878 10004 26884 10016
rect 26936 10004 26942 10056
rect 28534 10044 28540 10056
rect 28495 10016 28540 10044
rect 28534 10004 28540 10016
rect 28592 10004 28598 10056
rect 31110 10044 31116 10056
rect 31071 10016 31116 10044
rect 31110 10004 31116 10016
rect 31168 10004 31174 10056
rect 32214 10004 32220 10056
rect 32272 10044 32278 10056
rect 33045 10047 33103 10053
rect 33045 10044 33057 10047
rect 32272 10016 33057 10044
rect 32272 10004 32278 10016
rect 33045 10013 33057 10016
rect 33091 10044 33103 10047
rect 34072 10044 34100 10211
rect 35802 10208 35808 10220
rect 35860 10208 35866 10260
rect 36265 10251 36323 10257
rect 36265 10217 36277 10251
rect 36311 10248 36323 10251
rect 36354 10248 36360 10260
rect 36311 10220 36360 10248
rect 36311 10217 36323 10220
rect 36265 10211 36323 10217
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 36446 10208 36452 10260
rect 36504 10248 36510 10260
rect 36633 10251 36691 10257
rect 36633 10248 36645 10251
rect 36504 10220 36645 10248
rect 36504 10208 36510 10220
rect 36633 10217 36645 10220
rect 36679 10217 36691 10251
rect 36633 10211 36691 10217
rect 34698 10180 34704 10192
rect 34659 10152 34704 10180
rect 34698 10140 34704 10152
rect 34756 10140 34762 10192
rect 36078 10112 36084 10124
rect 36039 10084 36084 10112
rect 36078 10072 36084 10084
rect 36136 10072 36142 10124
rect 34606 10044 34612 10056
rect 33091 10016 34100 10044
rect 34567 10016 34612 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 34606 10004 34612 10016
rect 34664 10004 34670 10056
rect 34882 10044 34888 10056
rect 34843 10016 34888 10044
rect 34882 10004 34888 10016
rect 34940 10004 34946 10056
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 18782 9976 18788 9988
rect 9732 9948 18788 9976
rect 9732 9936 9738 9948
rect 18782 9936 18788 9948
rect 18840 9936 18846 9988
rect 7699 9911 7757 9917
rect 7699 9877 7711 9911
rect 7745 9908 7757 9911
rect 8202 9908 8208 9920
rect 7745 9880 8208 9908
rect 7745 9877 7757 9880
rect 7699 9871 7757 9877
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 8711 9911 8769 9917
rect 8711 9877 8723 9911
rect 8757 9908 8769 9911
rect 8846 9908 8852 9920
rect 8757 9880 8852 9908
rect 8757 9877 8769 9880
rect 8711 9871 8769 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 24118 9908 24124 9920
rect 24079 9880 24124 9908
rect 24118 9868 24124 9880
rect 24176 9868 24182 9920
rect 30098 9908 30104 9920
rect 30059 9880 30104 9908
rect 30098 9868 30104 9880
rect 30156 9868 30162 9920
rect 32398 9908 32404 9920
rect 32359 9880 32404 9908
rect 32398 9868 32404 9880
rect 32456 9868 32462 9920
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 5166 9704 5172 9716
rect 5127 9676 5172 9704
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 8904 9676 9597 9704
rect 8904 9664 8910 9676
rect 9585 9673 9597 9676
rect 9631 9704 9643 9707
rect 10502 9704 10508 9716
rect 9631 9676 10508 9704
rect 9631 9673 9643 9676
rect 9585 9667 9643 9673
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 11422 9704 11428 9716
rect 11383 9676 11428 9704
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11606 9664 11612 9716
rect 11664 9704 11670 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11664 9676 11805 9704
rect 11664 9664 11670 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 13725 9707 13783 9713
rect 13725 9673 13737 9707
rect 13771 9704 13783 9707
rect 14182 9704 14188 9716
rect 13771 9676 14188 9704
rect 13771 9673 13783 9676
rect 13725 9667 13783 9673
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 16209 9707 16267 9713
rect 16209 9704 16221 9707
rect 15712 9676 16221 9704
rect 15712 9664 15718 9676
rect 16209 9673 16221 9676
rect 16255 9673 16267 9707
rect 18782 9704 18788 9716
rect 18743 9676 18788 9704
rect 16209 9667 16267 9673
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 20162 9704 20168 9716
rect 20123 9676 20168 9704
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21910 9704 21916 9716
rect 21871 9676 21916 9704
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22741 9707 22799 9713
rect 22741 9673 22753 9707
rect 22787 9704 22799 9707
rect 23198 9704 23204 9716
rect 22787 9676 23204 9704
rect 22787 9673 22799 9676
rect 22741 9667 22799 9673
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 23474 9664 23480 9716
rect 23532 9704 23538 9716
rect 24946 9704 24952 9716
rect 23532 9676 24808 9704
rect 24907 9676 24952 9704
rect 23532 9664 23538 9676
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 2406 9636 2412 9648
rect 2087 9608 2412 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 2406 9596 2412 9608
rect 2464 9636 2470 9648
rect 5902 9645 5908 9648
rect 3973 9639 4031 9645
rect 3973 9636 3985 9639
rect 2464 9608 3985 9636
rect 2464 9596 2470 9608
rect 3973 9605 3985 9608
rect 4019 9605 4031 9639
rect 3973 9599 4031 9605
rect 5859 9639 5908 9645
rect 5859 9605 5871 9639
rect 5905 9605 5908 9639
rect 5859 9599 5908 9605
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9568 2378 9580
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2372 9540 3249 9568
rect 2372 9528 2378 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3988 9568 4016 9599
rect 5902 9596 5908 9599
rect 5960 9596 5966 9648
rect 11054 9636 11060 9648
rect 11015 9608 11060 9636
rect 11054 9596 11060 9608
rect 11112 9636 11118 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 11112 9608 12173 9636
rect 11112 9596 11118 9608
rect 12161 9605 12173 9608
rect 12207 9636 12219 9639
rect 12618 9636 12624 9648
rect 12207 9608 12624 9636
rect 12207 9605 12219 9608
rect 12161 9599 12219 9605
rect 12618 9596 12624 9608
rect 12676 9596 12682 9648
rect 13078 9636 13084 9648
rect 13039 9608 13084 9636
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15252 9608 15945 9636
rect 15252 9596 15258 9608
rect 15933 9605 15945 9608
rect 15979 9605 15991 9639
rect 16574 9636 16580 9648
rect 16535 9608 16580 9636
rect 15933 9599 15991 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 17126 9596 17132 9648
rect 17184 9636 17190 9648
rect 17862 9636 17868 9648
rect 17184 9608 17868 9636
rect 17184 9596 17190 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 6641 9571 6699 9577
rect 3988 9540 4660 9568
rect 3237 9531 3295 9537
rect 4632 9512 4660 9540
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 8665 9571 8723 9577
rect 6687 9540 7328 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 7300 9512 7328 9540
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 9030 9568 9036 9580
rect 8711 9540 9036 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 9030 9528 9036 9540
rect 9088 9528 9094 9580
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 10134 9568 10140 9580
rect 10095 9540 10140 9568
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 15010 9568 15016 9580
rect 14424 9540 15016 9568
rect 14424 9528 14430 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 19150 9528 19156 9580
rect 19208 9568 19214 9580
rect 19245 9571 19303 9577
rect 19245 9568 19257 9571
rect 19208 9540 19257 9568
rect 19208 9528 19214 9540
rect 19245 9537 19257 9540
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 20993 9571 21051 9577
rect 20993 9537 21005 9571
rect 21039 9568 21051 9571
rect 21266 9568 21272 9580
rect 21039 9540 21272 9568
rect 21039 9537 21051 9540
rect 20993 9531 21051 9537
rect 21266 9528 21272 9540
rect 21324 9528 21330 9580
rect 21928 9568 21956 9664
rect 23109 9639 23167 9645
rect 23109 9605 23121 9639
rect 23155 9636 23167 9639
rect 23290 9636 23296 9648
rect 23155 9608 23296 9636
rect 23155 9605 23167 9608
rect 23109 9599 23167 9605
rect 23290 9596 23296 9608
rect 23348 9636 23354 9648
rect 24581 9639 24639 9645
rect 24581 9636 24593 9639
rect 23348 9608 24593 9636
rect 23348 9596 23354 9608
rect 24581 9605 24593 9608
rect 24627 9605 24639 9639
rect 24780 9636 24808 9676
rect 24946 9664 24952 9676
rect 25004 9704 25010 9716
rect 25225 9707 25283 9713
rect 25225 9704 25237 9707
rect 25004 9676 25237 9704
rect 25004 9664 25010 9676
rect 25225 9673 25237 9676
rect 25271 9673 25283 9707
rect 26878 9704 26884 9716
rect 25225 9667 25283 9673
rect 26252 9676 26884 9704
rect 26252 9636 26280 9676
rect 26878 9664 26884 9676
rect 26936 9664 26942 9716
rect 30374 9664 30380 9716
rect 30432 9704 30438 9716
rect 30837 9707 30895 9713
rect 30837 9704 30849 9707
rect 30432 9676 30849 9704
rect 30432 9664 30438 9676
rect 30837 9673 30849 9676
rect 30883 9673 30895 9707
rect 30837 9667 30895 9673
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33229 9707 33287 9713
rect 33229 9704 33241 9707
rect 33192 9676 33241 9704
rect 33192 9664 33198 9676
rect 33229 9673 33241 9676
rect 33275 9704 33287 9707
rect 33505 9707 33563 9713
rect 33505 9704 33517 9707
rect 33275 9676 33517 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33505 9673 33517 9676
rect 33551 9673 33563 9707
rect 34606 9704 34612 9716
rect 33505 9667 33563 9673
rect 34440 9676 34612 9704
rect 24780 9608 26280 9636
rect 27157 9639 27215 9645
rect 24581 9599 24639 9605
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 21928 9540 22201 9568
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 25498 9568 25504 9580
rect 24728 9540 25504 9568
rect 24728 9528 24734 9540
rect 25498 9528 25504 9540
rect 25556 9528 25562 9580
rect 25792 9577 25820 9608
rect 27157 9605 27169 9639
rect 27203 9636 27215 9639
rect 27982 9636 27988 9648
rect 27203 9608 27988 9636
rect 27203 9605 27215 9608
rect 27157 9599 27215 9605
rect 27982 9596 27988 9608
rect 28040 9596 28046 9648
rect 28721 9639 28779 9645
rect 28721 9605 28733 9639
rect 28767 9636 28779 9639
rect 28810 9636 28816 9648
rect 28767 9608 28816 9636
rect 28767 9605 28779 9608
rect 28721 9599 28779 9605
rect 28810 9596 28816 9608
rect 28868 9636 28874 9648
rect 30193 9639 30251 9645
rect 28868 9608 28948 9636
rect 28868 9596 28874 9608
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 3697 9503 3755 9509
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 4433 9503 4491 9509
rect 4433 9500 4445 9503
rect 3743 9472 4445 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 4433 9469 4445 9472
rect 4479 9500 4491 9503
rect 4522 9500 4528 9512
rect 4479 9472 4528 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 4522 9460 4528 9472
rect 4580 9460 4586 9512
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5626 9500 5632 9512
rect 4672 9472 4765 9500
rect 5587 9472 5632 9500
rect 4672 9460 4678 9472
rect 5626 9460 5632 9472
rect 5684 9500 5690 9512
rect 5756 9503 5814 9509
rect 5756 9500 5768 9503
rect 5684 9472 5768 9500
rect 5684 9460 5690 9472
rect 5756 9469 5768 9472
rect 5802 9469 5814 9503
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 5756 9463 5814 9469
rect 6196 9472 6837 9500
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 2961 9435 3019 9441
rect 2464 9404 2509 9432
rect 2464 9392 2470 9404
rect 2961 9401 2973 9435
rect 3007 9432 3019 9435
rect 3326 9432 3332 9444
rect 3007 9404 3332 9432
rect 3007 9401 3019 9404
rect 2961 9395 3019 9401
rect 3326 9392 3332 9404
rect 3384 9392 3390 9444
rect 6196 9376 6224 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 7282 9500 7288 9512
rect 7195 9472 7288 9500
rect 6825 9463 6883 9469
rect 7282 9460 7288 9472
rect 7340 9460 7346 9512
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 14036 9503 14094 9509
rect 14036 9500 14048 9503
rect 13596 9472 14048 9500
rect 13596 9460 13602 9472
rect 14036 9469 14048 9472
rect 14082 9500 14094 9503
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14082 9472 14473 9500
rect 14082 9469 14094 9472
rect 14036 9463 14094 9469
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 16942 9460 16948 9512
rect 17000 9509 17006 9512
rect 17000 9503 17038 9509
rect 17026 9500 17038 9503
rect 17402 9500 17408 9512
rect 17026 9472 17408 9500
rect 17026 9469 17038 9472
rect 17000 9463 17038 9469
rect 17000 9460 17006 9463
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 18300 9503 18358 9509
rect 18300 9469 18312 9503
rect 18346 9500 18358 9503
rect 18782 9500 18788 9512
rect 18346 9472 18788 9500
rect 18346 9469 18358 9472
rect 18300 9463 18358 9469
rect 18782 9460 18788 9472
rect 18840 9460 18846 9512
rect 23014 9460 23020 9512
rect 23072 9500 23078 9512
rect 23661 9503 23719 9509
rect 23661 9500 23673 9503
rect 23072 9472 23673 9500
rect 23072 9460 23078 9472
rect 23661 9469 23673 9472
rect 23707 9500 23719 9503
rect 24118 9500 24124 9512
rect 23707 9472 24124 9500
rect 23707 9469 23719 9472
rect 23661 9463 23719 9469
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 27893 9503 27951 9509
rect 27893 9469 27905 9503
rect 27939 9469 27951 9503
rect 28000 9500 28028 9596
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9568 28411 9571
rect 28534 9568 28540 9580
rect 28399 9540 28540 9568
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 28534 9528 28540 9540
rect 28592 9528 28598 9580
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 28000 9472 28089 9500
rect 27893 9463 27951 9469
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 8754 9432 8760 9444
rect 8715 9404 8760 9432
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 10458 9435 10516 9441
rect 10458 9432 10470 9435
rect 9968 9404 10470 9432
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 2130 9364 2136 9376
rect 1719 9336 2136 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 4212 9336 4261 9364
rect 4212 9324 4218 9336
rect 4249 9333 4261 9336
rect 4295 9333 4307 9367
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 4249 9327 4307 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6880 9336 6929 9364
rect 6880 9324 6886 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7834 9364 7840 9376
rect 7432 9336 7840 9364
rect 7432 9324 7438 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8386 9364 8392 9376
rect 8347 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 9968 9373 9996 9404
rect 10458 9401 10470 9404
rect 10504 9401 10516 9435
rect 10458 9395 10516 9401
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 14921 9435 14979 9441
rect 12676 9404 12721 9432
rect 12676 9392 12682 9404
rect 14921 9401 14933 9435
rect 14967 9432 14979 9435
rect 15375 9435 15433 9441
rect 15375 9432 15387 9435
rect 14967 9404 15387 9432
rect 14967 9401 14979 9404
rect 14921 9395 14979 9401
rect 15375 9401 15387 9404
rect 15421 9432 15433 9435
rect 15930 9432 15936 9444
rect 15421 9404 15936 9432
rect 15421 9401 15433 9404
rect 15375 9395 15433 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 19607 9435 19665 9441
rect 19607 9432 19619 9435
rect 19168 9404 19619 9432
rect 19168 9376 19196 9404
rect 19607 9401 19619 9404
rect 19653 9432 19665 9435
rect 20901 9435 20959 9441
rect 20901 9432 20913 9435
rect 19653 9404 20913 9432
rect 19653 9401 19665 9404
rect 19607 9395 19665 9401
rect 20901 9401 20913 9404
rect 20947 9432 20959 9435
rect 21314 9435 21372 9441
rect 21314 9432 21326 9435
rect 20947 9404 21326 9432
rect 20947 9401 20959 9404
rect 20901 9395 20959 9401
rect 21314 9401 21326 9404
rect 21360 9401 21372 9435
rect 21314 9395 21372 9401
rect 23982 9435 24040 9441
rect 23982 9401 23994 9435
rect 24028 9401 24040 9435
rect 23982 9395 24040 9401
rect 25593 9435 25651 9441
rect 25593 9401 25605 9435
rect 25639 9401 25651 9435
rect 25593 9395 25651 9401
rect 27525 9435 27583 9441
rect 27525 9401 27537 9435
rect 27571 9432 27583 9435
rect 27908 9432 27936 9463
rect 28166 9432 28172 9444
rect 27571 9404 28172 9432
rect 27571 9401 27583 9404
rect 27525 9395 27583 9401
rect 9953 9367 10011 9373
rect 9953 9364 9965 9367
rect 9824 9336 9965 9364
rect 9824 9324 9830 9336
rect 9953 9333 9965 9336
rect 9999 9333 10011 9367
rect 9953 9327 10011 9333
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14139 9367 14197 9373
rect 14139 9364 14151 9367
rect 13964 9336 14151 9364
rect 13964 9324 13970 9336
rect 14139 9333 14151 9336
rect 14185 9333 14197 9367
rect 14139 9327 14197 9333
rect 17083 9367 17141 9373
rect 17083 9333 17095 9367
rect 17129 9364 17141 9367
rect 17310 9364 17316 9376
rect 17129 9336 17316 9364
rect 17129 9333 17141 9336
rect 17083 9327 17141 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 18371 9367 18429 9373
rect 18371 9333 18383 9367
rect 18417 9364 18429 9367
rect 18690 9364 18696 9376
rect 18417 9336 18696 9364
rect 18417 9333 18429 9336
rect 18371 9327 18429 9333
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 19150 9364 19156 9376
rect 19111 9336 19156 9364
rect 19150 9324 19156 9336
rect 19208 9324 19214 9376
rect 19334 9324 19340 9376
rect 19392 9364 19398 9376
rect 19794 9364 19800 9376
rect 19392 9336 19800 9364
rect 19392 9324 19398 9336
rect 19794 9324 19800 9336
rect 19852 9364 19858 9376
rect 20533 9367 20591 9373
rect 20533 9364 20545 9367
rect 19852 9336 20545 9364
rect 19852 9324 19858 9336
rect 20533 9333 20545 9336
rect 20579 9364 20591 9367
rect 21450 9364 21456 9376
rect 20579 9336 21456 9364
rect 20579 9333 20591 9336
rect 20533 9327 20591 9333
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23658 9364 23664 9376
rect 23523 9336 23664 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23658 9324 23664 9336
rect 23716 9364 23722 9376
rect 23997 9364 24025 9395
rect 23716 9336 24025 9364
rect 23716 9324 23722 9336
rect 24946 9324 24952 9376
rect 25004 9364 25010 9376
rect 25608 9364 25636 9395
rect 28166 9392 28172 9404
rect 28224 9392 28230 9444
rect 28920 9432 28948 9608
rect 30193 9605 30205 9639
rect 30239 9636 30251 9639
rect 30558 9636 30564 9648
rect 30239 9608 30564 9636
rect 30239 9605 30251 9608
rect 30193 9599 30251 9605
rect 30558 9596 30564 9608
rect 30616 9596 30622 9648
rect 31478 9645 31484 9648
rect 31435 9639 31484 9645
rect 31435 9605 31447 9639
rect 31481 9605 31484 9639
rect 31435 9599 31484 9605
rect 31478 9596 31484 9599
rect 31536 9596 31542 9648
rect 33965 9639 34023 9645
rect 33965 9605 33977 9639
rect 34011 9636 34023 9639
rect 34440 9636 34468 9676
rect 34606 9664 34612 9676
rect 34664 9664 34670 9716
rect 34011 9608 34468 9636
rect 34011 9605 34023 9608
rect 33965 9599 34023 9605
rect 34882 9596 34888 9648
rect 34940 9636 34946 9648
rect 34940 9608 35296 9636
rect 34940 9596 34946 9608
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29273 9571 29331 9577
rect 29273 9568 29285 9571
rect 29052 9540 29285 9568
rect 29052 9528 29058 9540
rect 29273 9537 29285 9540
rect 29319 9537 29331 9571
rect 29273 9531 29331 9537
rect 32309 9571 32367 9577
rect 32309 9537 32321 9571
rect 32355 9568 32367 9571
rect 32674 9568 32680 9580
rect 32355 9540 32680 9568
rect 32355 9537 32367 9540
rect 32309 9531 32367 9537
rect 32674 9528 32680 9540
rect 32732 9528 32738 9580
rect 34146 9528 34152 9580
rect 34204 9568 34210 9580
rect 34977 9571 35035 9577
rect 34977 9568 34989 9571
rect 34204 9540 34989 9568
rect 34204 9528 34210 9540
rect 34977 9537 34989 9540
rect 35023 9568 35035 9571
rect 35158 9568 35164 9580
rect 35023 9540 35164 9568
rect 35023 9537 35035 9540
rect 34977 9531 35035 9537
rect 35158 9528 35164 9540
rect 35216 9528 35222 9580
rect 35268 9577 35296 9608
rect 35253 9571 35311 9577
rect 35253 9537 35265 9571
rect 35299 9537 35311 9571
rect 35253 9531 35311 9537
rect 35894 9528 35900 9580
rect 35952 9568 35958 9580
rect 36817 9571 36875 9577
rect 36817 9568 36829 9571
rect 35952 9540 36829 9568
rect 35952 9528 35958 9540
rect 36817 9537 36829 9540
rect 36863 9537 36875 9571
rect 36817 9531 36875 9537
rect 30742 9460 30748 9512
rect 30800 9500 30806 9512
rect 31332 9503 31390 9509
rect 31332 9500 31344 9503
rect 30800 9472 31344 9500
rect 30800 9460 30806 9472
rect 31332 9469 31344 9472
rect 31378 9500 31390 9503
rect 31849 9503 31907 9509
rect 31849 9500 31861 9503
rect 31378 9472 31861 9500
rect 31378 9469 31390 9472
rect 31332 9463 31390 9469
rect 31849 9469 31861 9472
rect 31895 9500 31907 9503
rect 33042 9500 33048 9512
rect 31895 9472 33048 9500
rect 31895 9469 31907 9472
rect 31849 9463 31907 9469
rect 33042 9460 33048 9472
rect 33100 9460 33106 9512
rect 36078 9500 36084 9512
rect 36039 9472 36084 9500
rect 36078 9460 36084 9472
rect 36136 9460 36142 9512
rect 29089 9435 29147 9441
rect 29089 9432 29101 9435
rect 28920 9404 29101 9432
rect 29089 9401 29101 9404
rect 29135 9432 29147 9435
rect 29178 9432 29184 9444
rect 29135 9404 29184 9432
rect 29135 9401 29147 9404
rect 29089 9395 29147 9401
rect 29178 9392 29184 9404
rect 29236 9432 29242 9444
rect 32674 9441 32680 9444
rect 29635 9435 29693 9441
rect 29635 9432 29647 9435
rect 29236 9404 29647 9432
rect 29236 9392 29242 9404
rect 29635 9401 29647 9404
rect 29681 9432 29693 9435
rect 32217 9435 32275 9441
rect 32217 9432 32229 9435
rect 29681 9404 32229 9432
rect 29681 9401 29693 9404
rect 29635 9395 29693 9401
rect 32217 9401 32229 9404
rect 32263 9432 32275 9435
rect 32671 9432 32680 9441
rect 32263 9404 32680 9432
rect 32263 9401 32275 9404
rect 32217 9395 32275 9401
rect 32671 9395 32680 9404
rect 32674 9392 32680 9395
rect 32732 9392 32738 9444
rect 34701 9435 34759 9441
rect 34701 9401 34713 9435
rect 34747 9432 34759 9435
rect 35066 9432 35072 9444
rect 34747 9404 35072 9432
rect 34747 9401 34759 9404
rect 34701 9395 34759 9401
rect 35066 9392 35072 9404
rect 35124 9432 35130 9444
rect 36354 9432 36360 9444
rect 35124 9404 36360 9432
rect 35124 9392 35130 9404
rect 36354 9392 36360 9404
rect 36412 9392 36418 9444
rect 36538 9432 36544 9444
rect 36499 9404 36544 9432
rect 36538 9392 36544 9404
rect 36596 9392 36602 9444
rect 36633 9435 36691 9441
rect 36633 9401 36645 9435
rect 36679 9432 36691 9435
rect 36722 9432 36728 9444
rect 36679 9404 36728 9432
rect 36679 9401 36691 9404
rect 36633 9395 36691 9401
rect 36722 9392 36728 9404
rect 36780 9392 36786 9444
rect 26510 9364 26516 9376
rect 25004 9336 25636 9364
rect 26471 9336 26516 9364
rect 25004 9324 25010 9336
rect 26510 9324 26516 9336
rect 26568 9324 26574 9376
rect 34330 9364 34336 9376
rect 34291 9336 34336 9364
rect 34330 9324 34336 9336
rect 34388 9324 34394 9376
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 6972 9132 7573 9160
rect 6972 9120 6978 9132
rect 7561 9129 7573 9132
rect 7607 9160 7619 9163
rect 8113 9163 8171 9169
rect 8113 9160 8125 9163
rect 7607 9132 8125 9160
rect 7607 9129 7619 9132
rect 7561 9123 7619 9129
rect 8113 9129 8125 9132
rect 8159 9129 8171 9163
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 8113 9123 8171 9129
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 10873 9163 10931 9169
rect 10873 9160 10885 9163
rect 10836 9132 10885 9160
rect 10836 9120 10842 9132
rect 10873 9129 10885 9132
rect 10919 9129 10931 9163
rect 10873 9123 10931 9129
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11664 9132 11989 9160
rect 11664 9120 11670 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 11977 9123 12035 9129
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 15010 9160 15016 9172
rect 14971 9132 15016 9160
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16632 9132 16681 9160
rect 16632 9120 16638 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 17586 9160 17592 9172
rect 17547 9132 17592 9160
rect 16669 9123 16727 9129
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 18690 9160 18696 9172
rect 18651 9132 18696 9160
rect 18690 9120 18696 9132
rect 18748 9160 18754 9172
rect 20714 9160 20720 9172
rect 18748 9132 19012 9160
rect 20675 9132 20720 9160
rect 18748 9120 18754 9132
rect 2590 9092 2596 9104
rect 2551 9064 2596 9092
rect 2590 9052 2596 9064
rect 2648 9052 2654 9104
rect 5074 9092 5080 9104
rect 5035 9064 5080 9092
rect 5074 9052 5080 9064
rect 5132 9052 5138 9104
rect 6546 9092 6552 9104
rect 6507 9064 6552 9092
rect 6546 9052 6552 9064
rect 6604 9052 6610 9104
rect 6638 9052 6644 9104
rect 6696 9092 6702 9104
rect 9815 9095 9873 9101
rect 6696 9064 6741 9092
rect 6696 9052 6702 9064
rect 9815 9061 9827 9095
rect 9861 9092 9873 9095
rect 10226 9092 10232 9104
rect 9861 9064 10232 9092
rect 9861 9061 9873 9064
rect 9815 9055 9873 9061
rect 10226 9052 10232 9064
rect 10284 9052 10290 9104
rect 11238 9052 11244 9104
rect 11296 9092 11302 9104
rect 11378 9095 11436 9101
rect 11378 9092 11390 9095
rect 11296 9064 11390 9092
rect 11296 9052 11302 9064
rect 11378 9061 11390 9064
rect 11424 9061 11436 9095
rect 13814 9092 13820 9104
rect 13775 9064 13820 9092
rect 11378 9055 11436 9061
rect 13814 9052 13820 9064
rect 13872 9052 13878 9104
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 14918 9092 14924 9104
rect 14415 9064 14924 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 15930 9052 15936 9104
rect 15988 9092 15994 9104
rect 18984 9101 19012 9132
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 21266 9120 21272 9172
rect 21324 9160 21330 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21324 9132 21833 9160
rect 21324 9120 21330 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 24854 9120 24860 9172
rect 24912 9160 24918 9172
rect 25041 9163 25099 9169
rect 25041 9160 25053 9163
rect 24912 9132 25053 9160
rect 24912 9120 24918 9132
rect 25041 9129 25053 9132
rect 25087 9129 25099 9163
rect 25041 9123 25099 9129
rect 25130 9120 25136 9172
rect 25188 9160 25194 9172
rect 26605 9163 26663 9169
rect 26605 9160 26617 9163
rect 25188 9132 26617 9160
rect 25188 9120 25194 9132
rect 26605 9129 26617 9132
rect 26651 9129 26663 9163
rect 28534 9160 28540 9172
rect 28495 9132 28540 9160
rect 26605 9123 26663 9129
rect 28534 9120 28540 9132
rect 28592 9120 28598 9172
rect 29549 9163 29607 9169
rect 29549 9129 29561 9163
rect 29595 9160 29607 9163
rect 30098 9160 30104 9172
rect 29595 9132 30104 9160
rect 29595 9129 29607 9132
rect 29549 9123 29607 9129
rect 30098 9120 30104 9132
rect 30156 9120 30162 9172
rect 35158 9120 35164 9172
rect 35216 9160 35222 9172
rect 35253 9163 35311 9169
rect 35253 9160 35265 9163
rect 35216 9132 35265 9160
rect 35216 9120 35222 9132
rect 35253 9129 35265 9132
rect 35299 9129 35311 9163
rect 36354 9160 36360 9172
rect 36315 9132 36360 9160
rect 35253 9123 35311 9129
rect 36354 9120 36360 9132
rect 36412 9120 36418 9172
rect 36722 9160 36728 9172
rect 36683 9132 36728 9160
rect 36722 9120 36728 9132
rect 36780 9120 36786 9172
rect 16070 9095 16128 9101
rect 16070 9092 16082 9095
rect 15988 9064 16082 9092
rect 15988 9052 15994 9064
rect 16070 9061 16082 9064
rect 16116 9061 16128 9095
rect 16070 9055 16128 9061
rect 18969 9095 19027 9101
rect 18969 9061 18981 9095
rect 19015 9061 19027 9095
rect 18969 9055 19027 9061
rect 19058 9052 19064 9104
rect 19116 9092 19122 9104
rect 23014 9092 23020 9104
rect 19116 9064 19161 9092
rect 22975 9064 23020 9092
rect 19116 9052 19122 9064
rect 23014 9052 23020 9064
rect 23072 9052 23078 9104
rect 23658 9052 23664 9104
rect 23716 9092 23722 9104
rect 24166 9095 24224 9101
rect 24166 9092 24178 9095
rect 23716 9064 24178 9092
rect 23716 9052 23722 9064
rect 24166 9061 24178 9064
rect 24212 9061 24224 9095
rect 25498 9092 25504 9104
rect 25459 9064 25504 9092
rect 24166 9055 24224 9061
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 28991 9095 29049 9101
rect 28991 9061 29003 9095
rect 29037 9092 29049 9095
rect 29178 9092 29184 9104
rect 29037 9064 29184 9092
rect 29037 9061 29049 9064
rect 28991 9055 29049 9061
rect 29178 9052 29184 9064
rect 29236 9052 29242 9104
rect 31205 9095 31263 9101
rect 31205 9061 31217 9095
rect 31251 9092 31263 9095
rect 32766 9092 32772 9104
rect 31251 9064 32772 9092
rect 31251 9061 31263 9064
rect 31205 9055 31263 9061
rect 32766 9052 32772 9064
rect 32824 9092 32830 9104
rect 33137 9095 33195 9101
rect 33137 9092 33149 9095
rect 32824 9064 33149 9092
rect 32824 9052 32830 9064
rect 33137 9061 33149 9064
rect 33183 9061 33195 9095
rect 33137 9055 33195 9061
rect 34051 9095 34109 9101
rect 34051 9061 34063 9095
rect 34097 9092 34109 9095
rect 34146 9092 34152 9104
rect 34097 9064 34152 9092
rect 34097 9061 34109 9064
rect 34051 9055 34109 9061
rect 34146 9052 34152 9064
rect 34204 9052 34210 9104
rect 35799 9095 35857 9101
rect 35799 9061 35811 9095
rect 35845 9092 35857 9095
rect 35894 9092 35900 9104
rect 35845 9064 35900 9092
rect 35845 9061 35857 9064
rect 35799 9055 35857 9061
rect 35894 9052 35900 9064
rect 35952 9052 35958 9104
rect 1486 9033 1492 9036
rect 1464 9027 1492 9033
rect 1464 8993 1476 9027
rect 1464 8987 1492 8993
rect 1486 8984 1492 8987
rect 1544 8984 1550 9036
rect 8110 9024 8116 9036
rect 8071 8996 8116 9024
rect 8110 8984 8116 8996
rect 8168 8984 8174 9036
rect 8294 8984 8300 9036
rect 8352 9024 8358 9036
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8352 8996 8493 9024
rect 8352 8984 8358 8996
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 9674 8984 9680 9036
rect 9732 9033 9738 9036
rect 9732 9027 9770 9033
rect 9758 8993 9770 9027
rect 9732 8987 9770 8993
rect 11057 9027 11115 9033
rect 11057 8993 11069 9027
rect 11103 9024 11115 9027
rect 12342 9024 12348 9036
rect 11103 8996 12348 9024
rect 11103 8993 11115 8996
rect 11057 8987 11115 8993
rect 9732 8984 9738 8987
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 15746 9024 15752 9036
rect 15707 8996 15752 9024
rect 15746 8984 15752 8996
rect 15804 8984 15810 9036
rect 17862 8984 17868 9036
rect 17920 9033 17926 9036
rect 17920 9027 17958 9033
rect 17946 8993 17958 9027
rect 17920 8987 17958 8993
rect 17920 8984 17926 8987
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 20936 9027 20994 9033
rect 20936 9024 20948 9027
rect 20772 8996 20948 9024
rect 20772 8984 20778 8996
rect 20936 8993 20948 8996
rect 20982 9024 20994 9027
rect 21266 9024 21272 9036
rect 20982 8996 21272 9024
rect 20982 8993 20994 8996
rect 20936 8987 20994 8993
rect 21266 8984 21272 8996
rect 21324 8984 21330 9036
rect 22554 9024 22560 9036
rect 22515 8996 22560 9024
rect 22554 8984 22560 8996
rect 22612 8984 22618 9036
rect 22738 9024 22744 9036
rect 22699 8996 22744 9024
rect 22738 8984 22744 8996
rect 22796 8984 22802 9036
rect 24765 9027 24823 9033
rect 24765 8993 24777 9027
rect 24811 9024 24823 9027
rect 24946 9024 24952 9036
rect 24811 8996 24952 9024
rect 24811 8993 24823 8996
rect 24765 8987 24823 8993
rect 24946 8984 24952 8996
rect 25004 8984 25010 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 26970 9024 26976 9036
rect 26931 8996 26976 9024
rect 26970 8984 26976 8996
rect 27028 8984 27034 9036
rect 28350 8984 28356 9036
rect 28408 9024 28414 9036
rect 28629 9027 28687 9033
rect 28629 9024 28641 9027
rect 28408 8996 28641 9024
rect 28408 8984 28414 8996
rect 28629 8993 28641 8996
rect 28675 8993 28687 9027
rect 30466 9024 30472 9036
rect 30427 8996 30472 9024
rect 28629 8987 28687 8993
rect 30466 8984 30472 8996
rect 30524 8984 30530 9036
rect 30926 9024 30932 9036
rect 30887 8996 30932 9024
rect 30926 8984 30932 8996
rect 30984 8984 30990 9036
rect 32122 9024 32128 9036
rect 32083 8996 32128 9024
rect 32122 8984 32128 8996
rect 32180 8984 32186 9036
rect 32398 8984 32404 9036
rect 32456 9024 32462 9036
rect 32585 9027 32643 9033
rect 32585 9024 32597 9027
rect 32456 8996 32597 9024
rect 32456 8984 32462 8996
rect 32585 8993 32597 8996
rect 32631 8993 32643 9027
rect 32585 8987 32643 8993
rect 34330 8984 34336 9036
rect 34388 9024 34394 9036
rect 34609 9027 34667 9033
rect 34609 9024 34621 9027
rect 34388 8996 34621 9024
rect 34388 8984 34394 8996
rect 34609 8993 34621 8996
rect 34655 9024 34667 9027
rect 34698 9024 34704 9036
rect 34655 8996 34704 9024
rect 34655 8993 34667 8996
rect 34609 8987 34667 8993
rect 34698 8984 34704 8996
rect 34756 9024 34762 9036
rect 36740 9024 36768 9120
rect 34756 8996 36768 9024
rect 34756 8984 34762 8996
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2682 8956 2688 8968
rect 2547 8928 2688 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8956 2930 8968
rect 4709 8959 4767 8965
rect 4709 8956 4721 8959
rect 2924 8928 4721 8956
rect 2924 8916 2930 8928
rect 4709 8925 4721 8928
rect 4755 8956 4767 8959
rect 4798 8956 4804 8968
rect 4755 8928 4804 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4798 8916 4804 8928
rect 4856 8956 4862 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5166 8916 5172 8968
rect 5224 8956 5230 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5224 8928 5273 8956
rect 5224 8916 5230 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 5307 8928 6837 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 13722 8956 13728 8968
rect 13683 8928 13728 8956
rect 6825 8919 6883 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 19978 8956 19984 8968
rect 19939 8928 19984 8956
rect 19978 8916 19984 8928
rect 20036 8916 20042 8968
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 25130 8956 25136 8968
rect 23891 8928 25136 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 25130 8916 25136 8928
rect 25188 8916 25194 8968
rect 26329 8959 26387 8965
rect 26329 8925 26341 8959
rect 26375 8956 26387 8959
rect 26602 8956 26608 8968
rect 26375 8928 26608 8956
rect 26375 8925 26387 8928
rect 26329 8919 26387 8925
rect 26602 8916 26608 8928
rect 26660 8916 26666 8968
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 33505 8959 33563 8965
rect 33505 8956 33517 8959
rect 32907 8928 33517 8956
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33505 8925 33517 8928
rect 33551 8956 33563 8959
rect 33689 8959 33747 8965
rect 33689 8956 33701 8959
rect 33551 8928 33701 8956
rect 33551 8925 33563 8928
rect 33505 8919 33563 8925
rect 33689 8925 33701 8928
rect 33735 8925 33747 8959
rect 33689 8919 33747 8925
rect 34054 8916 34060 8968
rect 34112 8956 34118 8968
rect 35437 8959 35495 8965
rect 35437 8956 35449 8959
rect 34112 8928 35449 8956
rect 34112 8916 34118 8928
rect 35437 8925 35449 8928
rect 35483 8956 35495 8959
rect 36262 8956 36268 8968
rect 35483 8928 36268 8956
rect 35483 8925 35495 8928
rect 35437 8919 35495 8925
rect 36262 8916 36268 8928
rect 36320 8916 36326 8968
rect 18003 8891 18061 8897
rect 18003 8857 18015 8891
rect 18049 8888 18061 8891
rect 18966 8888 18972 8900
rect 18049 8860 18972 8888
rect 18049 8857 18061 8860
rect 18003 8851 18061 8857
rect 18966 8848 18972 8860
rect 19024 8848 19030 8900
rect 19518 8888 19524 8900
rect 19479 8860 19524 8888
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 1535 8823 1593 8829
rect 1535 8789 1547 8823
rect 1581 8820 1593 8823
rect 1854 8820 1860 8832
rect 1581 8792 1860 8820
rect 1581 8789 1593 8792
rect 1535 8783 1593 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2314 8820 2320 8832
rect 2275 8792 2320 8820
rect 2314 8780 2320 8792
rect 2372 8780 2378 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8812 8792 9137 8820
rect 8812 8780 8818 8792
rect 9125 8789 9137 8792
rect 9171 8820 9183 8823
rect 10594 8820 10600 8832
rect 9171 8792 10600 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 12802 8820 12808 8832
rect 12763 8792 12808 8820
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 14090 8820 14096 8832
rect 13587 8792 14096 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 18414 8820 18420 8832
rect 18375 8792 18420 8820
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21039 8823 21097 8829
rect 21039 8820 21051 8823
rect 20772 8792 21051 8820
rect 20772 8780 20778 8792
rect 21039 8789 21051 8792
rect 21085 8789 21097 8823
rect 21542 8820 21548 8832
rect 21503 8792 21548 8820
rect 21039 8783 21097 8789
rect 21542 8780 21548 8792
rect 21600 8780 21606 8832
rect 23658 8820 23664 8832
rect 23619 8792 23664 8820
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 27706 8820 27712 8832
rect 27667 8792 27712 8820
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 30101 8823 30159 8829
rect 30101 8789 30113 8823
rect 30147 8820 30159 8823
rect 30190 8820 30196 8832
rect 30147 8792 30196 8820
rect 30147 8789 30159 8792
rect 30101 8783 30159 8789
rect 30190 8780 30196 8792
rect 30248 8780 30254 8832
rect 34698 8780 34704 8832
rect 34756 8820 34762 8832
rect 34885 8823 34943 8829
rect 34885 8820 34897 8823
rect 34756 8792 34897 8820
rect 34756 8780 34762 8792
rect 34885 8789 34897 8792
rect 34931 8789 34943 8823
rect 34885 8783 34943 8789
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 3142 8616 3148 8628
rect 2648 8588 3148 8616
rect 2648 8576 2654 8588
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3200 8588 3249 8616
rect 3200 8576 3206 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3237 8579 3295 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 6273 8619 6331 8625
rect 6273 8585 6285 8619
rect 6319 8616 6331 8619
rect 6546 8616 6552 8628
rect 6319 8588 6552 8616
rect 6319 8585 6331 8588
rect 6273 8579 6331 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8352 8588 8493 8616
rect 8352 8576 8358 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 9030 8576 9036 8628
rect 9088 8616 9094 8628
rect 9171 8619 9229 8625
rect 9171 8616 9183 8619
rect 9088 8588 9183 8616
rect 9088 8576 9094 8588
rect 9171 8585 9183 8588
rect 9217 8585 9229 8619
rect 9171 8579 9229 8585
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9732 8588 9873 8616
rect 9732 8576 9738 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 10965 8619 11023 8625
rect 10965 8616 10977 8619
rect 10652 8588 10977 8616
rect 10652 8576 10658 8588
rect 10965 8585 10977 8588
rect 11011 8585 11023 8619
rect 10965 8579 11023 8585
rect 11701 8619 11759 8625
rect 11701 8585 11713 8619
rect 11747 8616 11759 8619
rect 12342 8616 12348 8628
rect 11747 8588 12348 8616
rect 11747 8585 11759 8588
rect 11701 8579 11759 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13814 8616 13820 8628
rect 13771 8588 13820 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13814 8576 13820 8588
rect 13872 8616 13878 8628
rect 14001 8619 14059 8625
rect 14001 8616 14013 8619
rect 13872 8588 14013 8616
rect 13872 8576 13878 8588
rect 14001 8585 14013 8588
rect 14047 8585 14059 8619
rect 14001 8579 14059 8585
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 15804 8588 17325 8616
rect 15804 8576 15810 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17313 8579 17371 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 19245 8619 19303 8625
rect 19245 8585 19257 8619
rect 19291 8616 19303 8619
rect 19426 8616 19432 8628
rect 19291 8588 19432 8616
rect 19291 8585 19303 8588
rect 19245 8579 19303 8585
rect 19426 8576 19432 8588
rect 19484 8576 19490 8628
rect 20625 8619 20683 8625
rect 20625 8585 20637 8619
rect 20671 8616 20683 8619
rect 20806 8616 20812 8628
rect 20671 8588 20812 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 21358 8616 21364 8628
rect 21319 8588 21364 8616
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22796 8588 22845 8616
rect 22796 8576 22802 8588
rect 22833 8585 22845 8588
rect 22879 8616 22891 8619
rect 23474 8616 23480 8628
rect 22879 8588 23480 8616
rect 22879 8585 22891 8588
rect 22833 8579 22891 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 24394 8576 24400 8628
rect 24452 8616 24458 8628
rect 24581 8619 24639 8625
rect 24581 8616 24593 8619
rect 24452 8588 24593 8616
rect 24452 8576 24458 8588
rect 24581 8585 24593 8588
rect 24627 8585 24639 8619
rect 24581 8579 24639 8585
rect 24949 8619 25007 8625
rect 24949 8585 24961 8619
rect 24995 8616 25007 8619
rect 25130 8616 25136 8628
rect 24995 8588 25136 8616
rect 24995 8585 25007 8588
rect 24949 8579 25007 8585
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25406 8576 25412 8628
rect 25464 8616 25470 8628
rect 25501 8619 25559 8625
rect 25501 8616 25513 8619
rect 25464 8588 25513 8616
rect 25464 8576 25470 8588
rect 25501 8585 25513 8588
rect 25547 8585 25559 8619
rect 25501 8579 25559 8585
rect 2866 8548 2872 8560
rect 2827 8520 2872 8548
rect 2866 8508 2872 8520
rect 2924 8508 2930 8560
rect 5166 8508 5172 8560
rect 5224 8548 5230 8560
rect 15473 8551 15531 8557
rect 5224 8520 5580 8548
rect 5224 8508 5230 8520
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1912 8452 2329 8480
rect 1912 8440 1918 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 2740 8452 3617 8480
rect 2740 8440 2746 8452
rect 3605 8449 3617 8452
rect 3651 8449 3663 8483
rect 3605 8443 3663 8449
rect 5077 8483 5135 8489
rect 5077 8449 5089 8483
rect 5123 8480 5135 8483
rect 5350 8480 5356 8492
rect 5123 8452 5356 8480
rect 5123 8449 5135 8452
rect 5077 8443 5135 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5552 8489 5580 8520
rect 15473 8517 15485 8551
rect 15519 8517 15531 8551
rect 15473 8511 15531 8517
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 5537 8443 5595 8449
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 10778 8480 10784 8492
rect 10091 8452 10784 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 12802 8480 12808 8492
rect 12763 8452 12808 8480
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 15488 8480 15516 8511
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16117 8551 16175 8557
rect 16117 8548 16129 8551
rect 16080 8520 16129 8548
rect 16080 8508 16086 8520
rect 16117 8517 16129 8520
rect 16163 8517 16175 8551
rect 16117 8511 16175 8517
rect 15488 8452 17264 8480
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 3835 8384 4169 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 7834 8412 7840 8424
rect 7795 8384 7840 8412
rect 4157 8375 4215 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 9068 8415 9126 8421
rect 9068 8412 9080 8415
rect 8904 8384 9080 8412
rect 8904 8372 8910 8384
rect 9068 8381 9080 8384
rect 9114 8412 9126 8415
rect 9490 8412 9496 8424
rect 9114 8384 9496 8412
rect 9114 8381 9126 8384
rect 9068 8375 9126 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 14642 8412 14648 8424
rect 14599 8384 14648 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 14642 8372 14648 8384
rect 14700 8372 14706 8424
rect 16022 8372 16028 8424
rect 16080 8412 16086 8424
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 16080 8384 16313 8412
rect 16080 8372 16086 8384
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 16942 8412 16948 8424
rect 16899 8384 16948 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 2314 8344 2320 8356
rect 2179 8316 2320 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 2314 8304 2320 8316
rect 2372 8344 2378 8356
rect 2409 8347 2467 8353
rect 2409 8344 2421 8347
rect 2372 8316 2421 8344
rect 2372 8304 2378 8316
rect 2409 8313 2421 8316
rect 2455 8344 2467 8347
rect 2682 8344 2688 8356
rect 2455 8316 2688 8344
rect 2455 8313 2467 8316
rect 2409 8307 2467 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 3384 8316 5273 8344
rect 3384 8304 3390 8316
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4433 8279 4491 8285
rect 4433 8276 4445 8279
rect 4203 8248 4445 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4433 8245 4445 8248
rect 4479 8276 4491 8279
rect 4890 8276 4896 8288
rect 4479 8248 4896 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4890 8236 4896 8248
rect 4948 8236 4954 8288
rect 5276 8276 5304 8307
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 6641 8347 6699 8353
rect 5408 8316 5453 8344
rect 5408 8304 5414 8316
rect 6641 8313 6653 8347
rect 6687 8344 6699 8347
rect 7190 8344 7196 8356
rect 6687 8316 7196 8344
rect 6687 8313 6699 8316
rect 6641 8307 6699 8313
rect 7190 8304 7196 8316
rect 7248 8353 7254 8356
rect 7248 8347 7296 8353
rect 7248 8313 7250 8347
rect 7284 8344 7296 8347
rect 7284 8316 7341 8344
rect 7284 8313 7296 8316
rect 7248 8307 7296 8313
rect 7248 8304 7254 8307
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10366 8347 10424 8353
rect 10366 8344 10378 8347
rect 9824 8316 10378 8344
rect 9824 8304 9830 8316
rect 10366 8313 10378 8316
rect 10412 8344 10424 8347
rect 11238 8344 11244 8356
rect 10412 8316 11244 8344
rect 10412 8313 10424 8316
rect 10366 8307 10424 8313
rect 11238 8304 11244 8316
rect 11296 8344 11302 8356
rect 12713 8347 12771 8353
rect 12713 8344 12725 8347
rect 11296 8316 12725 8344
rect 11296 8304 11302 8316
rect 12713 8313 12725 8316
rect 12759 8344 12771 8347
rect 13167 8347 13225 8353
rect 13167 8344 13179 8347
rect 12759 8316 13179 8344
rect 12759 8313 12771 8316
rect 12713 8307 12771 8313
rect 13167 8313 13179 8316
rect 13213 8344 13225 8347
rect 14461 8347 14519 8353
rect 14461 8344 14473 8347
rect 13213 8316 14473 8344
rect 13213 8313 13225 8316
rect 13167 8307 13225 8313
rect 14461 8313 14473 8316
rect 14507 8344 14519 8347
rect 14915 8347 14973 8353
rect 14915 8344 14927 8347
rect 14507 8316 14927 8344
rect 14507 8313 14519 8316
rect 14461 8307 14519 8313
rect 14915 8313 14927 8316
rect 14961 8344 14973 8347
rect 17034 8344 17040 8356
rect 14961 8316 15792 8344
rect 16995 8316 17040 8344
rect 14961 8313 14973 8316
rect 14915 8307 14973 8313
rect 15764 8288 15792 8316
rect 17034 8304 17040 8316
rect 17092 8304 17098 8356
rect 17236 8344 17264 8452
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 17368 8452 18245 8480
rect 17368 8440 17374 8452
rect 18233 8449 18245 8452
rect 18279 8480 18291 8483
rect 18506 8480 18512 8492
rect 18279 8452 18512 8480
rect 18279 8449 18291 8452
rect 18233 8443 18291 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18598 8440 18604 8492
rect 18656 8480 18662 8492
rect 19444 8480 19472 8576
rect 20993 8551 21051 8557
rect 20993 8517 21005 8551
rect 21039 8548 21051 8551
rect 21266 8548 21272 8560
rect 21039 8520 21272 8548
rect 21039 8517 21051 8520
rect 20993 8511 21051 8517
rect 21266 8508 21272 8520
rect 21324 8508 21330 8560
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 18656 8452 18701 8480
rect 19444 8452 19717 8480
rect 18656 8440 18662 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 25516 8480 25544 8579
rect 26970 8576 26976 8628
rect 27028 8616 27034 8628
rect 27065 8619 27123 8625
rect 27065 8616 27077 8619
rect 27028 8588 27077 8616
rect 27028 8576 27034 8588
rect 27065 8585 27077 8588
rect 27111 8585 27123 8619
rect 27065 8579 27123 8585
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 28997 8619 29055 8625
rect 28997 8616 29009 8619
rect 28408 8588 29009 8616
rect 28408 8576 28414 8588
rect 28997 8585 29009 8588
rect 29043 8585 29055 8619
rect 28997 8579 29055 8585
rect 31662 8576 31668 8628
rect 31720 8625 31726 8628
rect 31720 8619 31769 8625
rect 31720 8585 31723 8619
rect 31757 8616 31769 8619
rect 31757 8588 31813 8616
rect 31757 8585 31769 8588
rect 31720 8579 31769 8585
rect 31720 8576 31726 8579
rect 31846 8576 31852 8628
rect 31904 8616 31910 8628
rect 32122 8616 32128 8628
rect 31904 8588 32128 8616
rect 31904 8576 31910 8588
rect 32122 8576 32128 8588
rect 32180 8576 32186 8628
rect 34057 8619 34115 8625
rect 34057 8585 34069 8619
rect 34103 8616 34115 8619
rect 34146 8616 34152 8628
rect 34103 8588 34152 8616
rect 34103 8585 34115 8588
rect 34057 8579 34115 8585
rect 34146 8576 34152 8588
rect 34204 8616 34210 8628
rect 35894 8616 35900 8628
rect 34204 8588 35900 8616
rect 34204 8576 34210 8588
rect 35894 8576 35900 8588
rect 35952 8576 35958 8628
rect 36262 8616 36268 8628
rect 36223 8588 36268 8616
rect 36262 8576 36268 8588
rect 36320 8576 36326 8628
rect 36630 8616 36636 8628
rect 36591 8588 36636 8616
rect 36630 8576 36636 8588
rect 36688 8576 36694 8628
rect 26510 8508 26516 8560
rect 26568 8548 26574 8560
rect 27433 8551 27491 8557
rect 27433 8548 27445 8551
rect 26568 8520 27445 8548
rect 26568 8508 26574 8520
rect 27433 8517 27445 8520
rect 27479 8548 27491 8551
rect 28074 8548 28080 8560
rect 27479 8520 28080 8548
rect 27479 8517 27491 8520
rect 27433 8511 27491 8517
rect 25777 8483 25835 8489
rect 25777 8480 25789 8483
rect 25516 8452 25789 8480
rect 19705 8443 19763 8449
rect 25777 8449 25789 8452
rect 25823 8449 25835 8483
rect 25777 8443 25835 8449
rect 26421 8483 26479 8489
rect 26421 8449 26433 8483
rect 26467 8480 26479 8483
rect 27062 8480 27068 8492
rect 26467 8452 27068 8480
rect 26467 8449 26479 8452
rect 26421 8443 26479 8449
rect 27062 8440 27068 8452
rect 27120 8440 27126 8492
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19208 8384 19656 8412
rect 19208 8372 19214 8384
rect 18325 8347 18383 8353
rect 18325 8344 18337 8347
rect 17236 8316 18337 8344
rect 18325 8313 18337 8316
rect 18371 8344 18383 8347
rect 18414 8344 18420 8356
rect 18371 8316 18420 8344
rect 18371 8313 18383 8316
rect 18325 8307 18383 8313
rect 18414 8304 18420 8316
rect 18472 8304 18478 8356
rect 18690 8304 18696 8356
rect 18748 8344 18754 8356
rect 19058 8344 19064 8356
rect 18748 8316 19064 8344
rect 18748 8304 18754 8316
rect 19058 8304 19064 8316
rect 19116 8304 19122 8356
rect 19628 8344 19656 8384
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 21416 8384 21465 8412
rect 21416 8372 21422 8384
rect 21453 8381 21465 8384
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 21600 8384 21925 8412
rect 21600 8372 21606 8384
rect 21913 8381 21925 8384
rect 21959 8381 21971 8415
rect 21913 8375 21971 8381
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8412 23719 8415
rect 24210 8412 24216 8424
rect 23707 8384 24216 8412
rect 23707 8381 23719 8384
rect 23661 8375 23719 8381
rect 24210 8372 24216 8384
rect 24268 8372 24274 8424
rect 20026 8347 20084 8353
rect 20026 8344 20038 8347
rect 19628 8316 20038 8344
rect 19628 8288 19656 8316
rect 20026 8313 20038 8316
rect 20072 8313 20084 8347
rect 20026 8307 20084 8313
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 21560 8344 21588 8372
rect 22554 8344 22560 8356
rect 20588 8316 21588 8344
rect 22515 8316 22560 8344
rect 20588 8304 20594 8316
rect 22554 8304 22560 8316
rect 22612 8304 22618 8356
rect 23982 8347 24040 8353
rect 23982 8313 23994 8347
rect 24028 8344 24040 8347
rect 24028 8316 24062 8344
rect 24028 8313 24040 8316
rect 23982 8307 24040 8313
rect 5534 8276 5540 8288
rect 5276 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 7374 8276 7380 8288
rect 6144 8248 7380 8276
rect 6144 8236 6150 8248
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 15746 8276 15752 8288
rect 15707 8248 15752 8276
rect 15746 8236 15752 8248
rect 15804 8276 15810 8288
rect 15930 8276 15936 8288
rect 15804 8248 15936 8276
rect 15804 8236 15810 8248
rect 15930 8236 15936 8248
rect 15988 8236 15994 8288
rect 18046 8236 18052 8288
rect 18104 8276 18110 8288
rect 19426 8276 19432 8288
rect 18104 8248 19432 8276
rect 18104 8236 18110 8248
rect 19426 8236 19432 8248
rect 19484 8236 19490 8288
rect 19610 8276 19616 8288
rect 19571 8248 19616 8276
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 21542 8276 21548 8288
rect 21503 8248 21548 8276
rect 21542 8236 21548 8248
rect 21600 8236 21606 8288
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23658 8276 23664 8288
rect 23523 8248 23664 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23658 8236 23664 8248
rect 23716 8276 23722 8288
rect 23997 8276 24025 8307
rect 25866 8304 25872 8356
rect 25924 8344 25930 8356
rect 25924 8316 25969 8344
rect 25924 8304 25930 8316
rect 26050 8304 26056 8356
rect 26108 8344 26114 8356
rect 26510 8344 26516 8356
rect 26108 8316 26516 8344
rect 26108 8304 26114 8316
rect 26510 8304 26516 8316
rect 26568 8344 26574 8356
rect 26697 8347 26755 8353
rect 26697 8344 26709 8347
rect 26568 8316 26709 8344
rect 26568 8304 26574 8316
rect 26697 8313 26709 8316
rect 26743 8313 26755 8347
rect 27080 8344 27108 8440
rect 27448 8412 27476 8511
rect 28074 8508 28080 8520
rect 28132 8508 28138 8560
rect 30374 8480 30380 8492
rect 28092 8452 30380 8480
rect 27617 8415 27675 8421
rect 27617 8412 27629 8415
rect 27448 8384 27629 8412
rect 27617 8381 27629 8384
rect 27663 8381 27675 8415
rect 27617 8375 27675 8381
rect 27706 8372 27712 8424
rect 27764 8412 27770 8424
rect 28092 8421 28120 8452
rect 30374 8440 30380 8452
rect 30432 8480 30438 8492
rect 30926 8480 30932 8492
rect 30432 8452 30932 8480
rect 30432 8440 30438 8452
rect 30926 8440 30932 8452
rect 30984 8480 30990 8492
rect 31021 8483 31079 8489
rect 31021 8480 31033 8483
rect 30984 8452 31033 8480
rect 30984 8440 30990 8452
rect 31021 8449 31033 8452
rect 31067 8449 31079 8483
rect 32766 8480 32772 8492
rect 32727 8452 32772 8480
rect 31021 8443 31079 8449
rect 32766 8440 32772 8452
rect 32824 8440 32830 8492
rect 34698 8440 34704 8492
rect 34756 8480 34762 8492
rect 34977 8483 35035 8489
rect 34977 8480 34989 8483
rect 34756 8452 34989 8480
rect 34756 8440 34762 8452
rect 34977 8449 34989 8452
rect 35023 8449 35035 8483
rect 35250 8480 35256 8492
rect 35211 8452 35256 8480
rect 34977 8443 35035 8449
rect 35250 8440 35256 8452
rect 35308 8440 35314 8492
rect 28077 8415 28135 8421
rect 28077 8412 28089 8415
rect 27764 8384 28089 8412
rect 27764 8372 27770 8384
rect 28077 8381 28089 8384
rect 28123 8381 28135 8415
rect 28077 8375 28135 8381
rect 28353 8415 28411 8421
rect 28353 8381 28365 8415
rect 28399 8412 28411 8415
rect 28994 8412 29000 8424
rect 28399 8384 29000 8412
rect 28399 8381 28411 8384
rect 28353 8375 28411 8381
rect 28994 8372 29000 8384
rect 29052 8372 29058 8424
rect 31570 8412 31576 8424
rect 31628 8421 31634 8424
rect 31628 8415 31666 8421
rect 31404 8384 31576 8412
rect 28721 8347 28779 8353
rect 27080 8316 27568 8344
rect 26697 8307 26755 8313
rect 24670 8276 24676 8288
rect 23716 8248 24676 8276
rect 23716 8236 23722 8248
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 27540 8276 27568 8316
rect 28721 8313 28733 8347
rect 28767 8344 28779 8347
rect 28902 8344 28908 8356
rect 28767 8316 28908 8344
rect 28767 8313 28779 8316
rect 28721 8307 28779 8313
rect 28902 8304 28908 8316
rect 28960 8304 28966 8356
rect 29917 8347 29975 8353
rect 29917 8313 29929 8347
rect 29963 8344 29975 8347
rect 30101 8347 30159 8353
rect 30101 8344 30113 8347
rect 29963 8316 30113 8344
rect 29963 8313 29975 8316
rect 29917 8307 29975 8313
rect 30101 8313 30113 8316
rect 30147 8313 30159 8347
rect 30101 8307 30159 8313
rect 28074 8276 28080 8288
rect 27540 8248 28080 8276
rect 28074 8236 28080 8248
rect 28132 8236 28138 8288
rect 30116 8276 30144 8307
rect 30190 8304 30196 8356
rect 30248 8344 30254 8356
rect 31404 8353 31432 8384
rect 31570 8372 31576 8384
rect 31654 8381 31666 8415
rect 31628 8375 31666 8381
rect 33689 8415 33747 8421
rect 33689 8381 33701 8415
rect 33735 8412 33747 8415
rect 34609 8415 34667 8421
rect 34609 8412 34621 8415
rect 33735 8384 34621 8412
rect 33735 8381 33747 8384
rect 33689 8375 33747 8381
rect 34609 8381 34621 8384
rect 34655 8381 34667 8415
rect 34609 8375 34667 8381
rect 31628 8372 31634 8375
rect 30745 8347 30803 8353
rect 30248 8316 30293 8344
rect 30248 8304 30254 8316
rect 30745 8313 30757 8347
rect 30791 8344 30803 8347
rect 31389 8347 31447 8353
rect 31389 8344 31401 8347
rect 30791 8316 31401 8344
rect 30791 8313 30803 8316
rect 30745 8307 30803 8313
rect 31389 8313 31401 8316
rect 31435 8313 31447 8347
rect 32674 8344 32680 8356
rect 32587 8316 32680 8344
rect 31389 8307 31447 8313
rect 32674 8304 32680 8316
rect 32732 8344 32738 8356
rect 33131 8347 33189 8353
rect 33131 8344 33143 8347
rect 32732 8316 33143 8344
rect 32732 8304 32738 8316
rect 33131 8313 33143 8316
rect 33177 8344 33189 8347
rect 34146 8344 34152 8356
rect 33177 8316 34152 8344
rect 33177 8313 33189 8316
rect 33131 8307 33189 8313
rect 34146 8304 34152 8316
rect 34204 8304 34210 8356
rect 34624 8344 34652 8375
rect 36078 8372 36084 8424
rect 36136 8412 36142 8424
rect 36449 8415 36507 8421
rect 36449 8412 36461 8415
rect 36136 8384 36461 8412
rect 36136 8372 36142 8384
rect 36449 8381 36461 8384
rect 36495 8412 36507 8415
rect 37001 8415 37059 8421
rect 37001 8412 37013 8415
rect 36495 8384 37013 8412
rect 36495 8381 36507 8384
rect 36449 8375 36507 8381
rect 37001 8381 37013 8384
rect 37047 8381 37059 8415
rect 37001 8375 37059 8381
rect 35069 8347 35127 8353
rect 34624 8316 34928 8344
rect 30650 8276 30656 8288
rect 30116 8248 30656 8276
rect 30650 8236 30656 8248
rect 30708 8236 30714 8288
rect 34900 8276 34928 8316
rect 35069 8313 35081 8347
rect 35115 8313 35127 8347
rect 35069 8307 35127 8313
rect 35084 8276 35112 8307
rect 34900 8248 35112 8276
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4154 8072 4160 8084
rect 3927 8044 4160 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 5166 8072 5172 8084
rect 5127 8044 5172 8072
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5534 8072 5540 8084
rect 5495 8044 5540 8072
rect 5534 8032 5540 8044
rect 5592 8032 5598 8084
rect 5810 8072 5816 8084
rect 5771 8044 5816 8072
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6549 8075 6607 8081
rect 6549 8041 6561 8075
rect 6595 8072 6607 8075
rect 6638 8072 6644 8084
rect 6595 8044 6644 8072
rect 6595 8041 6607 8044
rect 6549 8035 6607 8041
rect 6638 8032 6644 8044
rect 6696 8072 6702 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 6696 8044 7757 8072
rect 6696 8032 6702 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 8711 8075 8769 8081
rect 8711 8041 8723 8075
rect 8757 8072 8769 8075
rect 8938 8072 8944 8084
rect 8757 8044 8944 8072
rect 8757 8041 8769 8044
rect 8711 8035 8769 8041
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 10778 8072 10784 8084
rect 10739 8044 10784 8072
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 13173 8075 13231 8081
rect 13173 8041 13185 8075
rect 13219 8072 13231 8075
rect 13722 8072 13728 8084
rect 13219 8044 13728 8072
rect 13219 8041 13231 8044
rect 13173 8035 13231 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14734 8072 14740 8084
rect 13832 8044 14740 8072
rect 2127 8007 2185 8013
rect 2127 7973 2139 8007
rect 2173 8004 2185 8007
rect 2314 8004 2320 8016
rect 2173 7976 2320 8004
rect 2173 7973 2185 7976
rect 2127 7967 2185 7973
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 4249 8007 4307 8013
rect 4249 7973 4261 8007
rect 4295 8004 4307 8007
rect 4430 8004 4436 8016
rect 4295 7976 4436 8004
rect 4295 7973 4307 7976
rect 4249 7967 4307 7973
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 4798 8004 4804 8016
rect 4759 7976 4804 8004
rect 4798 7964 4804 7976
rect 4856 7964 4862 8016
rect 7190 8013 7196 8016
rect 7187 8004 7196 8013
rect 7151 7976 7196 8004
rect 7187 7967 7196 7976
rect 7190 7964 7196 7967
rect 7248 7964 7254 8016
rect 13832 8004 13860 8044
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 16945 8075 17003 8081
rect 16945 8041 16957 8075
rect 16991 8072 17003 8075
rect 17034 8072 17040 8084
rect 16991 8044 17040 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 19058 8032 19064 8084
rect 19116 8072 19122 8084
rect 20073 8075 20131 8081
rect 20073 8072 20085 8075
rect 19116 8044 20085 8072
rect 19116 8032 19122 8044
rect 20073 8041 20085 8044
rect 20119 8041 20131 8075
rect 20073 8035 20131 8041
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 23845 8075 23903 8081
rect 23845 8072 23857 8075
rect 23532 8044 23857 8072
rect 23532 8032 23538 8044
rect 23845 8041 23857 8044
rect 23891 8072 23903 8075
rect 24118 8072 24124 8084
rect 23891 8044 24124 8072
rect 23891 8041 23903 8044
rect 23845 8035 23903 8041
rect 24118 8032 24124 8044
rect 24176 8032 24182 8084
rect 25409 8075 25467 8081
rect 25409 8041 25421 8075
rect 25455 8072 25467 8075
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25455 8044 25789 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 25777 8041 25789 8044
rect 25823 8072 25835 8075
rect 25866 8072 25872 8084
rect 25823 8044 25872 8072
rect 25823 8041 25835 8044
rect 25777 8035 25835 8041
rect 25866 8032 25872 8044
rect 25924 8032 25930 8084
rect 29825 8075 29883 8081
rect 29825 8041 29837 8075
rect 29871 8072 29883 8075
rect 30190 8072 30196 8084
rect 29871 8044 30196 8072
rect 29871 8041 29883 8044
rect 29825 8035 29883 8041
rect 30190 8032 30196 8044
rect 30248 8032 30254 8084
rect 30466 8072 30472 8084
rect 30427 8044 30472 8072
rect 30466 8032 30472 8044
rect 30524 8032 30530 8084
rect 30650 8072 30656 8084
rect 30611 8044 30656 8072
rect 30650 8032 30656 8044
rect 30708 8032 30714 8084
rect 32398 8072 32404 8084
rect 32359 8044 32404 8072
rect 32398 8032 32404 8044
rect 32456 8032 32462 8084
rect 34425 8075 34483 8081
rect 34425 8041 34437 8075
rect 34471 8072 34483 8075
rect 34471 8044 35480 8072
rect 34471 8041 34483 8044
rect 34425 8035 34483 8041
rect 35452 8016 35480 8044
rect 12360 7976 13860 8004
rect 14369 8007 14427 8013
rect 1762 7936 1768 7948
rect 1723 7908 1768 7936
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5718 7936 5724 7948
rect 5675 7908 5724 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 8640 7939 8698 7945
rect 8640 7905 8652 7939
rect 8686 7936 8698 7939
rect 9030 7936 9036 7948
rect 8686 7908 9036 7936
rect 8686 7905 8698 7908
rect 8640 7899 8698 7905
rect 9030 7896 9036 7908
rect 9088 7896 9094 7948
rect 10778 7936 10784 7948
rect 10739 7908 10784 7936
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 10962 7896 10968 7948
rect 11020 7936 11026 7948
rect 11020 7908 11113 7936
rect 11020 7896 11026 7908
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 12158 7936 12164 7948
rect 11204 7908 12164 7936
rect 11204 7896 11210 7908
rect 12158 7896 12164 7908
rect 12216 7936 12222 7948
rect 12360 7945 12388 7976
rect 14369 7973 14381 8007
rect 14415 8004 14427 8007
rect 14642 8004 14648 8016
rect 14415 7976 14648 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 14642 7964 14648 7976
rect 14700 7964 14706 8016
rect 15651 8007 15709 8013
rect 15651 7973 15663 8007
rect 15697 8004 15709 8007
rect 15746 8004 15752 8016
rect 15697 7976 15752 8004
rect 15697 7973 15709 7976
rect 15651 7967 15709 7973
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 17586 8004 17592 8016
rect 16224 7976 17592 8004
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 12216 7908 12357 7936
rect 12216 7896 12222 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 3559 7840 4169 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 4157 7837 4169 7840
rect 4203 7868 4215 7871
rect 4246 7868 4252 7880
rect 4203 7840 4252 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 6914 7868 6920 7880
rect 6871 7840 6920 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 9950 7828 9956 7880
rect 10008 7868 10014 7880
rect 10980 7868 11008 7896
rect 10008 7840 11008 7868
rect 10008 7828 10014 7840
rect 12636 7812 12664 7899
rect 12710 7896 12716 7948
rect 12768 7936 12774 7948
rect 13814 7936 13820 7948
rect 12768 7908 13820 7936
rect 12768 7896 12774 7908
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 13998 7896 14004 7948
rect 14056 7936 14062 7948
rect 16224 7945 16252 7976
rect 17586 7964 17592 7976
rect 17644 8004 17650 8016
rect 17681 8007 17739 8013
rect 17681 8004 17693 8007
rect 17644 7976 17693 8004
rect 17644 7964 17650 7976
rect 17681 7973 17693 7976
rect 17727 8004 17739 8007
rect 17727 7976 18736 8004
rect 17727 7973 17739 7976
rect 17681 7967 17739 7973
rect 18708 7948 18736 7976
rect 19150 7964 19156 8016
rect 19208 8004 19214 8016
rect 19254 8007 19312 8013
rect 19254 8004 19266 8007
rect 19208 7976 19266 8004
rect 19208 7964 19214 7976
rect 19254 7973 19266 7976
rect 19300 7973 19312 8007
rect 19254 7967 19312 7973
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 8004 21695 8007
rect 22002 8004 22008 8016
rect 21683 7976 22008 8004
rect 21683 7973 21695 7976
rect 21637 7967 21695 7973
rect 22002 7964 22008 7976
rect 22060 7964 22066 8016
rect 24670 7964 24676 8016
rect 24728 8004 24734 8016
rect 26878 8013 26884 8016
rect 24810 8007 24868 8013
rect 24810 8004 24822 8007
rect 24728 7976 24822 8004
rect 24728 7964 24734 7976
rect 24810 7973 24822 7976
rect 24856 7973 24868 8007
rect 26875 8004 26884 8013
rect 26839 7976 26884 8004
rect 24810 7967 24868 7973
rect 26875 7967 26884 7976
rect 26878 7964 26884 7967
rect 26936 7964 26942 8016
rect 29178 7964 29184 8016
rect 29236 8013 29242 8016
rect 29236 8007 29284 8013
rect 29236 7973 29238 8007
rect 29272 7973 29284 8007
rect 29236 7967 29284 7973
rect 33867 8007 33925 8013
rect 33867 7973 33879 8007
rect 33913 8004 33925 8007
rect 34146 8004 34152 8016
rect 33913 7976 34152 8004
rect 33913 7973 33925 7976
rect 33867 7967 33925 7973
rect 29236 7964 29242 7967
rect 34146 7964 34152 7976
rect 34204 7964 34210 8016
rect 35434 8004 35440 8016
rect 35347 7976 35440 8004
rect 35434 7964 35440 7976
rect 35492 7964 35498 8016
rect 35986 8004 35992 8016
rect 35947 7976 35992 8004
rect 35986 7964 35992 7976
rect 36044 7964 36050 8016
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 14056 7908 14105 7936
rect 14056 7896 14062 7908
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 16209 7939 16267 7945
rect 16209 7905 16221 7939
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 18877 7939 18935 7945
rect 18877 7936 18889 7939
rect 18748 7908 18889 7936
rect 18748 7896 18754 7908
rect 18877 7905 18889 7908
rect 18923 7905 18935 7939
rect 18877 7899 18935 7905
rect 22646 7896 22652 7948
rect 22704 7936 22710 7948
rect 23017 7939 23075 7945
rect 23017 7936 23029 7939
rect 22704 7908 23029 7936
rect 22704 7896 22710 7908
rect 23017 7905 23029 7908
rect 23063 7905 23075 7939
rect 23017 7899 23075 7905
rect 23201 7939 23259 7945
rect 23201 7905 23213 7939
rect 23247 7936 23259 7939
rect 23382 7936 23388 7948
rect 23247 7908 23388 7936
rect 23247 7905 23259 7908
rect 23201 7899 23259 7905
rect 23382 7896 23388 7908
rect 23440 7896 23446 7948
rect 28994 7896 29000 7948
rect 29052 7936 29058 7948
rect 30098 7936 30104 7948
rect 29052 7908 30104 7936
rect 29052 7896 29058 7908
rect 30098 7896 30104 7908
rect 30156 7896 30162 7948
rect 30558 7896 30564 7948
rect 30616 7936 30622 7948
rect 32560 7939 32618 7945
rect 32560 7936 32572 7939
rect 30616 7908 32572 7936
rect 30616 7896 30622 7908
rect 32560 7905 32572 7908
rect 32606 7936 32618 7939
rect 32766 7936 32772 7948
rect 32606 7908 32772 7936
rect 32606 7905 32618 7908
rect 32560 7899 32618 7905
rect 32766 7896 32772 7908
rect 32824 7936 32830 7948
rect 35158 7936 35164 7948
rect 32824 7908 35164 7936
rect 32824 7896 32830 7908
rect 35158 7896 35164 7908
rect 35216 7896 35222 7948
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 14550 7868 14556 7880
rect 12851 7840 14556 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 14550 7828 14556 7840
rect 14608 7868 14614 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 14608 7840 15301 7868
rect 14608 7828 14614 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 17589 7871 17647 7877
rect 17589 7837 17601 7871
rect 17635 7868 17647 7871
rect 17954 7868 17960 7880
rect 17635 7840 17960 7868
rect 17635 7837 17647 7840
rect 17589 7831 17647 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18233 7871 18291 7877
rect 18233 7837 18245 7871
rect 18279 7868 18291 7871
rect 18598 7868 18604 7880
rect 18279 7840 18604 7868
rect 18279 7837 18291 7840
rect 18233 7831 18291 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19153 7871 19211 7877
rect 19153 7868 19165 7871
rect 19024 7840 19165 7868
rect 19024 7828 19030 7840
rect 19153 7837 19165 7840
rect 19199 7837 19211 7871
rect 19518 7868 19524 7880
rect 19479 7840 19524 7868
rect 19153 7831 19211 7837
rect 19518 7828 19524 7840
rect 19576 7868 19582 7880
rect 21269 7871 21327 7877
rect 21269 7868 21281 7871
rect 19576 7840 21281 7868
rect 19576 7828 19582 7840
rect 21269 7837 21281 7840
rect 21315 7868 21327 7871
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 21315 7840 21557 7868
rect 21315 7837 21327 7840
rect 21269 7831 21327 7837
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7868 24547 7871
rect 25038 7868 25044 7880
rect 24535 7840 25044 7868
rect 24535 7837 24547 7840
rect 24489 7831 24547 7837
rect 12618 7800 12624 7812
rect 12531 7772 12624 7800
rect 12618 7760 12624 7772
rect 12676 7800 12682 7812
rect 12676 7772 14044 7800
rect 12676 7760 12682 7772
rect 14016 7744 14044 7772
rect 19058 7760 19064 7812
rect 19116 7760 19122 7812
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 23584 7800 23612 7831
rect 25038 7828 25044 7840
rect 25096 7828 25102 7880
rect 26510 7868 26516 7880
rect 26471 7840 26516 7868
rect 26510 7828 26516 7840
rect 26568 7828 26574 7880
rect 28718 7828 28724 7880
rect 28776 7868 28782 7880
rect 28905 7871 28963 7877
rect 28905 7868 28917 7871
rect 28776 7840 28917 7868
rect 28776 7828 28782 7840
rect 28905 7837 28917 7840
rect 28951 7837 28963 7871
rect 33502 7868 33508 7880
rect 33463 7840 33508 7868
rect 28905 7831 28963 7837
rect 33502 7828 33508 7840
rect 33560 7828 33566 7880
rect 35342 7868 35348 7880
rect 35303 7840 35348 7868
rect 35342 7828 35348 7840
rect 35400 7828 35406 7880
rect 24854 7800 24860 7812
rect 22152 7772 22197 7800
rect 23584 7772 24860 7800
rect 22152 7760 22158 7772
rect 24854 7760 24860 7772
rect 24912 7760 24918 7812
rect 31018 7760 31024 7812
rect 31076 7800 31082 7812
rect 33321 7803 33379 7809
rect 33321 7800 33333 7803
rect 31076 7772 33333 7800
rect 31076 7760 31082 7772
rect 33321 7769 33333 7772
rect 33367 7800 33379 7803
rect 33594 7800 33600 7812
rect 33367 7772 33600 7800
rect 33367 7769 33379 7772
rect 33321 7763 33379 7769
rect 33594 7760 33600 7772
rect 33652 7760 33658 7812
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 3510 7732 3516 7744
rect 3099 7704 3516 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 9824 7704 10057 7732
rect 9824 7692 9830 7704
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13630 7732 13636 7744
rect 13587 7704 13636 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 14056 7704 16589 7732
rect 14056 7692 14062 7704
rect 16577 7701 16589 7704
rect 16623 7732 16635 7735
rect 16942 7732 16948 7744
rect 16623 7704 16948 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 18414 7692 18420 7744
rect 18472 7732 18478 7744
rect 19076 7732 19104 7760
rect 19242 7732 19248 7744
rect 18472 7704 19248 7732
rect 18472 7692 18478 7704
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 22554 7732 22560 7744
rect 20864 7704 22560 7732
rect 20864 7692 20870 7704
rect 22554 7692 22560 7704
rect 22612 7732 22618 7744
rect 23290 7732 23296 7744
rect 22612 7704 23296 7732
rect 22612 7692 22618 7704
rect 23290 7692 23296 7704
rect 23348 7692 23354 7744
rect 24210 7732 24216 7744
rect 24171 7704 24216 7732
rect 24210 7692 24216 7704
rect 24268 7692 24274 7744
rect 27430 7732 27436 7744
rect 27391 7704 27436 7732
rect 27430 7692 27436 7704
rect 27488 7692 27494 7744
rect 27706 7732 27712 7744
rect 27667 7704 27712 7732
rect 27706 7692 27712 7704
rect 27764 7692 27770 7744
rect 32631 7735 32689 7741
rect 32631 7701 32643 7735
rect 32677 7732 32689 7735
rect 33134 7732 33140 7744
rect 32677 7704 33140 7732
rect 32677 7701 32689 7704
rect 32631 7695 32689 7701
rect 33134 7692 33140 7704
rect 33192 7692 33198 7744
rect 34882 7732 34888 7744
rect 34843 7704 34888 7732
rect 34882 7692 34888 7704
rect 34940 7692 34946 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 5718 7528 5724 7540
rect 5679 7500 5724 7528
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 8754 7528 8760 7540
rect 8715 7500 8760 7528
rect 8754 7488 8760 7500
rect 8812 7488 8818 7540
rect 9674 7528 9680 7540
rect 9635 7500 9680 7528
rect 9674 7488 9680 7500
rect 9732 7528 9738 7540
rect 10226 7528 10232 7540
rect 9732 7500 10232 7528
rect 9732 7488 9738 7500
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10778 7488 10784 7540
rect 10836 7528 10842 7540
rect 11149 7531 11207 7537
rect 11149 7528 11161 7531
rect 10836 7500 11161 7528
rect 10836 7488 10842 7500
rect 11149 7497 11161 7500
rect 11195 7497 11207 7531
rect 11149 7491 11207 7497
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 12618 7528 12624 7540
rect 11839 7500 12624 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13722 7528 13728 7540
rect 13495 7500 13728 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14550 7528 14556 7540
rect 14511 7500 14556 7528
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 15286 7528 15292 7540
rect 15247 7500 15292 7528
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 17586 7528 17592 7540
rect 17547 7500 17592 7528
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 19076 7500 20085 7528
rect 9950 7460 9956 7472
rect 9911 7432 9956 7460
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 12158 7460 12164 7472
rect 12119 7432 12164 7460
rect 12158 7420 12164 7432
rect 12216 7420 12222 7472
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 18782 7460 18788 7472
rect 13596 7432 18788 7460
rect 13596 7420 13602 7432
rect 18782 7420 18788 7432
rect 18840 7420 18846 7472
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 9088 7364 10517 7392
rect 9088 7352 9094 7364
rect 10505 7361 10517 7364
rect 10551 7392 10563 7395
rect 10962 7392 10968 7404
rect 10551 7364 10968 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 13909 7395 13967 7401
rect 13909 7392 13921 7395
rect 13872 7364 13921 7392
rect 13872 7352 13878 7364
rect 13909 7361 13921 7364
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 17034 7392 17040 7404
rect 16255 7364 17040 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 18693 7395 18751 7401
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 19076 7392 19104 7500
rect 20073 7497 20085 7500
rect 20119 7528 20131 7531
rect 20622 7528 20628 7540
rect 20119 7500 20628 7528
rect 20119 7497 20131 7500
rect 20073 7491 20131 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 22002 7488 22008 7540
rect 22060 7528 22066 7540
rect 22373 7531 22431 7537
rect 22373 7528 22385 7531
rect 22060 7500 22385 7528
rect 22060 7488 22066 7500
rect 22373 7497 22385 7500
rect 22419 7497 22431 7531
rect 22373 7491 22431 7497
rect 26878 7488 26884 7540
rect 26936 7528 26942 7540
rect 29089 7531 29147 7537
rect 29089 7528 29101 7531
rect 26936 7500 29101 7528
rect 26936 7488 26942 7500
rect 29089 7497 29101 7500
rect 29135 7497 29147 7531
rect 31018 7528 31024 7540
rect 30979 7500 31024 7528
rect 29089 7491 29147 7497
rect 31018 7488 31024 7500
rect 31076 7488 31082 7540
rect 32766 7528 32772 7540
rect 32727 7500 32772 7528
rect 32766 7488 32772 7500
rect 32824 7488 32830 7540
rect 34146 7488 34152 7540
rect 34204 7528 34210 7540
rect 34241 7531 34299 7537
rect 34241 7528 34253 7531
rect 34204 7500 34253 7528
rect 34204 7488 34210 7500
rect 34241 7497 34253 7500
rect 34287 7497 34299 7531
rect 34241 7491 34299 7497
rect 35434 7488 35440 7540
rect 35492 7528 35498 7540
rect 35897 7531 35955 7537
rect 35897 7528 35909 7531
rect 35492 7500 35909 7528
rect 35492 7488 35498 7500
rect 35897 7497 35909 7500
rect 35943 7497 35955 7531
rect 36630 7528 36636 7540
rect 36591 7500 36636 7528
rect 35897 7491 35955 7497
rect 36630 7488 36636 7500
rect 36688 7488 36694 7540
rect 19245 7463 19303 7469
rect 19245 7429 19257 7463
rect 19291 7460 19303 7463
rect 19518 7460 19524 7472
rect 19291 7432 19524 7460
rect 19291 7429 19303 7432
rect 19245 7423 19303 7429
rect 19518 7420 19524 7432
rect 19576 7420 19582 7472
rect 32355 7463 32413 7469
rect 32355 7429 32367 7463
rect 32401 7460 32413 7463
rect 34882 7460 34888 7472
rect 32401 7432 34888 7460
rect 32401 7429 32413 7432
rect 32355 7423 32413 7429
rect 34882 7420 34888 7432
rect 34940 7460 34946 7472
rect 34940 7432 35020 7460
rect 34940 7420 34946 7432
rect 18739 7364 19104 7392
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 20303 7395 20361 7401
rect 20303 7392 20315 7395
rect 19208 7364 20315 7392
rect 19208 7352 19214 7364
rect 20303 7361 20315 7364
rect 20349 7361 20361 7395
rect 20303 7355 20361 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 21542 7392 21548 7404
rect 21499 7364 21548 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 24210 7392 24216 7404
rect 24171 7364 24216 7392
rect 24210 7352 24216 7364
rect 24268 7352 24274 7404
rect 25869 7395 25927 7401
rect 25869 7361 25881 7395
rect 25915 7392 25927 7395
rect 26142 7392 26148 7404
rect 25915 7364 26148 7392
rect 25915 7361 25927 7364
rect 25869 7355 25927 7361
rect 26142 7352 26148 7364
rect 26200 7352 26206 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7392 27770 7404
rect 27982 7392 27988 7404
rect 27764 7364 27988 7392
rect 27764 7352 27770 7364
rect 27982 7352 27988 7364
rect 28040 7352 28046 7404
rect 28074 7352 28080 7404
rect 28132 7392 28138 7404
rect 30098 7392 30104 7404
rect 28132 7364 28177 7392
rect 30059 7364 30104 7392
rect 28132 7352 28138 7364
rect 30098 7352 30104 7364
rect 30156 7352 30162 7404
rect 32674 7392 32680 7404
rect 31623 7364 32680 7392
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7324 2283 7327
rect 3510 7324 3516 7336
rect 2271 7296 3516 7324
rect 2271 7293 2283 7296
rect 2225 7287 2283 7293
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6730 7324 6736 7336
rect 6687 7296 6736 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6730 7284 6736 7296
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8018 7324 8024 7336
rect 7883 7296 8024 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 12618 7333 12624 7336
rect 12596 7327 12624 7333
rect 12596 7293 12608 7327
rect 12676 7324 12682 7336
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 12676 7296 13124 7324
rect 12596 7287 12624 7293
rect 12618 7284 12624 7287
rect 12676 7284 12682 7296
rect 2546 7259 2604 7265
rect 2546 7256 2558 7259
rect 2332 7228 2558 7256
rect 2332 7200 2360 7228
rect 2546 7225 2558 7228
rect 2592 7225 2604 7259
rect 4478 7259 4536 7265
rect 4478 7256 4490 7259
rect 2546 7219 2604 7225
rect 3988 7228 4490 7256
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2314 7188 2320 7200
rect 1903 7160 2320 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2314 7148 2320 7160
rect 2372 7148 2378 7200
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 3602 7188 3608 7200
rect 3559 7160 3608 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 3602 7148 3608 7160
rect 3660 7188 3666 7200
rect 3988 7197 4016 7228
rect 4478 7225 4490 7228
rect 4524 7256 4536 7259
rect 5534 7256 5540 7268
rect 4524 7228 5540 7256
rect 4524 7225 4536 7228
rect 4478 7219 4536 7225
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 8158 7259 8216 7265
rect 8158 7256 8170 7259
rect 7668 7228 8170 7256
rect 3973 7191 4031 7197
rect 3973 7188 3985 7191
rect 3660 7160 3985 7188
rect 3660 7148 3666 7160
rect 3973 7157 3985 7160
rect 4019 7157 4031 7191
rect 5074 7188 5080 7200
rect 5035 7160 5080 7188
rect 3973 7151 4031 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6914 7188 6920 7200
rect 6319 7160 6920 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7098 7188 7104 7200
rect 7055 7160 7104 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 7668 7197 7696 7228
rect 8158 7225 8170 7228
rect 8204 7225 8216 7259
rect 10226 7256 10232 7268
rect 10187 7228 10232 7256
rect 8158 7219 8216 7225
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10321 7259 10379 7265
rect 10321 7225 10333 7259
rect 10367 7225 10379 7259
rect 10321 7219 10379 7225
rect 7285 7191 7343 7197
rect 7285 7188 7297 7191
rect 7248 7160 7297 7188
rect 7248 7148 7254 7160
rect 7285 7157 7297 7160
rect 7331 7188 7343 7191
rect 7653 7191 7711 7197
rect 7653 7188 7665 7191
rect 7331 7160 7665 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7653 7157 7665 7160
rect 7699 7157 7711 7191
rect 7653 7151 7711 7157
rect 9309 7191 9367 7197
rect 9309 7157 9321 7191
rect 9355 7188 9367 7191
rect 10336 7188 10364 7219
rect 13096 7200 13124 7296
rect 14936 7296 15117 7324
rect 13630 7256 13636 7268
rect 13591 7228 13636 7256
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 13780 7228 13825 7256
rect 13780 7216 13786 7228
rect 14936 7200 14964 7296
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15105 7287 15163 7293
rect 17129 7327 17187 7333
rect 17129 7293 17141 7327
rect 17175 7324 17187 7327
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 17175 7296 18429 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 15657 7259 15715 7265
rect 15657 7225 15669 7259
rect 15703 7256 15715 7259
rect 15746 7256 15752 7268
rect 15703 7228 15752 7256
rect 15703 7225 15715 7228
rect 15657 7219 15715 7225
rect 15746 7216 15752 7228
rect 15804 7256 15810 7268
rect 16574 7265 16580 7268
rect 16117 7259 16175 7265
rect 16117 7256 16129 7259
rect 15804 7228 16129 7256
rect 15804 7216 15810 7228
rect 16117 7225 16129 7228
rect 16163 7256 16175 7259
rect 16571 7256 16580 7265
rect 16163 7228 16580 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 16571 7219 16580 7228
rect 16574 7216 16580 7219
rect 16632 7216 16638 7268
rect 10594 7188 10600 7200
rect 9355 7160 10600 7188
rect 9355 7157 9367 7160
rect 9309 7151 9367 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 12667 7191 12725 7197
rect 12667 7157 12679 7191
rect 12713 7188 12725 7191
rect 12802 7188 12808 7200
rect 12713 7160 12808 7188
rect 12713 7157 12725 7160
rect 12667 7151 12725 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13078 7188 13084 7200
rect 13039 7160 13084 7188
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 14918 7188 14924 7200
rect 14879 7160 14924 7188
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 18432 7188 18460 7287
rect 20162 7284 20168 7336
rect 20220 7333 20226 7336
rect 20220 7327 20258 7333
rect 20246 7324 20258 7327
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 20246 7296 20637 7324
rect 20246 7293 20258 7296
rect 20220 7287 20258 7293
rect 20625 7293 20637 7296
rect 20671 7324 20683 7327
rect 22186 7324 22192 7336
rect 20671 7296 22192 7324
rect 20671 7293 20683 7296
rect 20625 7287 20683 7293
rect 20220 7284 20226 7287
rect 22186 7284 22192 7296
rect 22244 7284 22250 7336
rect 23109 7327 23167 7333
rect 23109 7293 23121 7327
rect 23155 7324 23167 7327
rect 23382 7324 23388 7336
rect 23155 7296 23388 7324
rect 23155 7293 23167 7296
rect 23109 7287 23167 7293
rect 23382 7284 23388 7296
rect 23440 7284 23446 7336
rect 23477 7327 23535 7333
rect 23477 7293 23489 7327
rect 23523 7324 23535 7327
rect 23934 7324 23940 7336
rect 23523 7296 23940 7324
rect 23523 7293 23535 7296
rect 23477 7287 23535 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 24118 7324 24124 7336
rect 24079 7296 24124 7324
rect 24118 7284 24124 7296
rect 24176 7284 24182 7336
rect 26789 7327 26847 7333
rect 26789 7293 26801 7327
rect 26835 7324 26847 7327
rect 27433 7327 27491 7333
rect 27433 7324 27445 7327
rect 26835 7296 27445 7324
rect 26835 7293 26847 7296
rect 26789 7287 26847 7293
rect 27433 7293 27445 7296
rect 27479 7293 27491 7327
rect 27433 7287 27491 7293
rect 18785 7259 18843 7265
rect 18785 7225 18797 7259
rect 18831 7225 18843 7259
rect 21358 7256 21364 7268
rect 21271 7228 21364 7256
rect 18785 7219 18843 7225
rect 18598 7188 18604 7200
rect 18432 7160 18604 7188
rect 18598 7148 18604 7160
rect 18656 7188 18662 7200
rect 18800 7188 18828 7219
rect 21358 7216 21364 7228
rect 21416 7256 21422 7268
rect 21815 7259 21873 7265
rect 21815 7256 21827 7259
rect 21416 7228 21827 7256
rect 21416 7216 21422 7228
rect 21815 7225 21827 7228
rect 21861 7256 21873 7259
rect 25685 7259 25743 7265
rect 25685 7256 25697 7259
rect 21861 7228 25697 7256
rect 21861 7225 21873 7228
rect 21815 7219 21873 7225
rect 24688 7200 24716 7228
rect 25685 7225 25697 7228
rect 25731 7256 25743 7259
rect 26190 7259 26248 7265
rect 26190 7256 26202 7259
rect 25731 7228 26202 7256
rect 25731 7225 25743 7228
rect 25685 7219 25743 7225
rect 26190 7225 26202 7228
rect 26236 7256 26248 7259
rect 26878 7256 26884 7268
rect 26236 7228 26884 7256
rect 26236 7225 26248 7228
rect 26190 7219 26248 7225
rect 26878 7216 26884 7228
rect 26936 7256 26942 7268
rect 27065 7259 27123 7265
rect 27065 7256 27077 7259
rect 26936 7228 27077 7256
rect 26936 7216 26942 7228
rect 27065 7225 27077 7228
rect 27111 7225 27123 7259
rect 27065 7219 27123 7225
rect 18656 7160 18828 7188
rect 18656 7148 18662 7160
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19300 7160 19625 7188
rect 19300 7148 19306 7160
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 22646 7188 22652 7200
rect 22607 7160 22652 7188
rect 19613 7151 19671 7157
rect 22646 7148 22652 7160
rect 22704 7148 22710 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 25038 7188 25044 7200
rect 24999 7160 25044 7188
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 27448 7188 27476 7287
rect 27801 7259 27859 7265
rect 27801 7225 27813 7259
rect 27847 7225 27859 7259
rect 27801 7219 27859 7225
rect 27816 7188 27844 7219
rect 28718 7216 28724 7268
rect 28776 7256 28782 7268
rect 29457 7259 29515 7265
rect 29457 7256 29469 7259
rect 28776 7228 29469 7256
rect 28776 7216 28782 7228
rect 29457 7225 29469 7228
rect 29503 7225 29515 7259
rect 29457 7219 29515 7225
rect 30009 7259 30067 7265
rect 30009 7225 30021 7259
rect 30055 7256 30067 7259
rect 30463 7259 30521 7265
rect 30463 7256 30475 7259
rect 30055 7228 30475 7256
rect 30055 7225 30067 7228
rect 30009 7219 30067 7225
rect 30463 7225 30475 7228
rect 30509 7256 30521 7259
rect 31623 7256 31651 7364
rect 32674 7352 32680 7364
rect 32732 7352 32738 7404
rect 33134 7352 33140 7404
rect 33192 7392 33198 7404
rect 34992 7401 35020 7432
rect 33321 7395 33379 7401
rect 33321 7392 33333 7395
rect 33192 7364 33333 7392
rect 33192 7352 33198 7364
rect 33321 7361 33333 7364
rect 33367 7361 33379 7395
rect 33321 7355 33379 7361
rect 34977 7395 35035 7401
rect 34977 7361 34989 7395
rect 35023 7361 35035 7395
rect 35342 7392 35348 7404
rect 35303 7364 35348 7392
rect 34977 7355 35035 7361
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 32030 7284 32036 7336
rect 32088 7324 32094 7336
rect 32284 7327 32342 7333
rect 32284 7324 32296 7327
rect 32088 7296 32296 7324
rect 32088 7284 32094 7296
rect 32284 7293 32296 7296
rect 32330 7324 32342 7327
rect 32493 7327 32551 7333
rect 32493 7324 32505 7327
rect 32330 7296 32505 7324
rect 32330 7293 32342 7296
rect 32284 7287 32342 7293
rect 32493 7293 32505 7296
rect 32539 7293 32551 7327
rect 32493 7287 32551 7293
rect 33965 7327 34023 7333
rect 33965 7293 33977 7327
rect 34011 7324 34023 7327
rect 34422 7324 34428 7336
rect 34011 7296 34428 7324
rect 34011 7293 34023 7296
rect 33965 7287 34023 7293
rect 34422 7284 34428 7296
rect 34480 7284 34486 7336
rect 36446 7324 36452 7336
rect 36359 7296 36452 7324
rect 36446 7284 36452 7296
rect 36504 7324 36510 7336
rect 37001 7327 37059 7333
rect 37001 7324 37013 7327
rect 36504 7296 37013 7324
rect 36504 7284 36510 7296
rect 37001 7293 37013 7296
rect 37047 7293 37059 7327
rect 37001 7287 37059 7293
rect 30509 7228 31651 7256
rect 33422 7259 33480 7265
rect 30509 7225 30521 7228
rect 30463 7219 30521 7225
rect 33422 7225 33434 7259
rect 33468 7256 33480 7259
rect 33594 7256 33600 7268
rect 33468 7228 33600 7256
rect 33468 7225 33480 7228
rect 33422 7219 33480 7225
rect 27448 7160 27844 7188
rect 28997 7191 29055 7197
rect 28997 7157 29009 7191
rect 29043 7188 29055 7191
rect 29089 7191 29147 7197
rect 29089 7188 29101 7191
rect 29043 7160 29101 7188
rect 29043 7157 29055 7160
rect 28997 7151 29055 7157
rect 29089 7157 29101 7160
rect 29135 7188 29147 7191
rect 30024 7188 30052 7219
rect 33594 7216 33600 7228
rect 33652 7256 33658 7268
rect 34609 7259 34667 7265
rect 34609 7256 34621 7259
rect 33652 7228 34621 7256
rect 33652 7216 33658 7228
rect 34609 7225 34621 7228
rect 34655 7256 34667 7259
rect 35069 7259 35127 7265
rect 35069 7256 35081 7259
rect 34655 7228 35081 7256
rect 34655 7225 34667 7228
rect 34609 7219 34667 7225
rect 35069 7225 35081 7228
rect 35115 7225 35127 7259
rect 35069 7219 35127 7225
rect 29135 7160 30052 7188
rect 32493 7191 32551 7197
rect 29135 7157 29147 7160
rect 29089 7151 29147 7157
rect 32493 7157 32505 7191
rect 32539 7188 32551 7191
rect 33137 7191 33195 7197
rect 33137 7188 33149 7191
rect 32539 7160 33149 7188
rect 32539 7157 32551 7160
rect 32493 7151 32551 7157
rect 33137 7157 33149 7160
rect 33183 7188 33195 7191
rect 33226 7188 33232 7200
rect 33183 7160 33232 7188
rect 33183 7157 33195 7160
rect 33137 7151 33195 7157
rect 33226 7148 33232 7160
rect 33284 7148 33290 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 1762 6984 1768 6996
rect 1723 6956 1768 6984
rect 1762 6944 1768 6956
rect 1820 6944 1826 6996
rect 10594 6984 10600 6996
rect 10555 6956 10600 6984
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 13998 6984 14004 6996
rect 13771 6956 14004 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 17497 6987 17555 6993
rect 17497 6953 17509 6987
rect 17543 6984 17555 6987
rect 17954 6984 17960 6996
rect 17543 6956 17960 6984
rect 17543 6953 17555 6956
rect 17497 6947 17555 6953
rect 17954 6944 17960 6956
rect 18012 6944 18018 6996
rect 22002 6984 22008 6996
rect 21963 6956 22008 6984
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 25961 6987 26019 6993
rect 25961 6953 25973 6987
rect 26007 6984 26019 6987
rect 26142 6984 26148 6996
rect 26007 6956 26148 6984
rect 26007 6953 26019 6956
rect 25961 6947 26019 6953
rect 26142 6944 26148 6956
rect 26200 6944 26206 6996
rect 33134 6944 33140 6996
rect 33192 6984 33198 6996
rect 33873 6987 33931 6993
rect 33873 6984 33885 6987
rect 33192 6956 33885 6984
rect 33192 6944 33198 6956
rect 33873 6953 33885 6956
rect 33919 6953 33931 6987
rect 35342 6984 35348 6996
rect 33873 6947 33931 6953
rect 35176 6956 35348 6984
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 2546 6919 2604 6925
rect 2546 6916 2558 6919
rect 2372 6888 2558 6916
rect 2372 6876 2378 6888
rect 2546 6885 2558 6888
rect 2592 6916 2604 6919
rect 3602 6916 3608 6928
rect 2592 6888 3608 6916
rect 2592 6885 2604 6888
rect 2546 6879 2604 6885
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 4430 6916 4436 6928
rect 4264 6888 4436 6916
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4154 6848 4160 6860
rect 3927 6820 4160 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 4154 6808 4160 6820
rect 4212 6848 4218 6860
rect 4264 6848 4292 6888
rect 4430 6876 4436 6888
rect 4488 6916 4494 6928
rect 4525 6919 4583 6925
rect 4525 6916 4537 6919
rect 4488 6888 4537 6916
rect 4488 6876 4494 6888
rect 4525 6885 4537 6888
rect 4571 6916 4583 6919
rect 5074 6916 5080 6928
rect 4571 6888 5080 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 6911 6919 6969 6925
rect 6911 6885 6923 6919
rect 6957 6916 6969 6919
rect 7190 6916 7196 6928
rect 6957 6888 7196 6916
rect 6957 6885 6969 6888
rect 6911 6879 6969 6885
rect 4212 6820 4292 6848
rect 4212 6808 4218 6820
rect 6638 6808 6644 6860
rect 6696 6848 6702 6860
rect 6932 6848 6960 6879
rect 7190 6876 7196 6888
rect 7248 6876 7254 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 9998 6919 10056 6925
rect 9998 6916 10010 6919
rect 9824 6888 10010 6916
rect 9824 6876 9830 6888
rect 9998 6885 10010 6888
rect 10044 6885 10056 6919
rect 9998 6879 10056 6885
rect 12339 6919 12397 6925
rect 12339 6885 12351 6919
rect 12385 6885 12397 6919
rect 12339 6879 12397 6885
rect 15841 6919 15899 6925
rect 15841 6885 15853 6919
rect 15887 6916 15899 6919
rect 16117 6919 16175 6925
rect 16117 6916 16129 6919
rect 15887 6888 16129 6916
rect 15887 6885 15899 6888
rect 15841 6879 15899 6885
rect 16117 6885 16129 6888
rect 16163 6916 16175 6919
rect 16298 6916 16304 6928
rect 16163 6888 16304 6916
rect 16163 6885 16175 6888
rect 16117 6879 16175 6885
rect 6696 6820 6960 6848
rect 8573 6851 8631 6857
rect 6696 6808 6702 6820
rect 8573 6817 8585 6851
rect 8619 6848 8631 6851
rect 8662 6848 8668 6860
rect 8619 6820 8668 6848
rect 8619 6817 8631 6820
rect 8573 6811 8631 6817
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12360 6848 12388 6879
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 19331 6919 19389 6925
rect 19331 6885 19343 6919
rect 19377 6916 19389 6919
rect 21085 6919 21143 6925
rect 21085 6916 21097 6919
rect 19377 6888 19411 6916
rect 20824 6888 21097 6916
rect 19377 6885 19389 6888
rect 19331 6879 19389 6885
rect 12124 6820 12388 6848
rect 14185 6851 14243 6857
rect 12124 6808 12130 6820
rect 14185 6817 14197 6851
rect 14231 6848 14243 6851
rect 15010 6848 15016 6860
rect 14231 6820 15016 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 17589 6851 17647 6857
rect 16724 6820 16769 6848
rect 16724 6808 16730 6820
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 17770 6848 17776 6860
rect 17731 6820 17776 6848
rect 17589 6811 17647 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2590 6780 2596 6792
rect 2271 6752 2596 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4433 6783 4491 6789
rect 4433 6780 4445 6783
rect 4120 6752 4445 6780
rect 4120 6740 4126 6752
rect 4433 6749 4445 6752
rect 4479 6780 4491 6783
rect 5258 6780 5264 6792
rect 4479 6752 5264 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6822 6780 6828 6792
rect 6595 6752 6828 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 9677 6783 9735 6789
rect 9677 6749 9689 6783
rect 9723 6780 9735 6783
rect 10226 6780 10232 6792
rect 9723 6752 10232 6780
rect 9723 6749 9735 6752
rect 9677 6743 9735 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 14826 6740 14832 6792
rect 14884 6780 14890 6792
rect 16025 6783 16083 6789
rect 16025 6780 16037 6783
rect 14884 6752 16037 6780
rect 14884 6740 14890 6752
rect 16025 6749 16037 6752
rect 16071 6780 16083 6783
rect 16850 6780 16856 6792
rect 16071 6752 16856 6780
rect 16071 6749 16083 6752
rect 16025 6743 16083 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4985 6715 5043 6721
rect 4985 6712 4997 6715
rect 3384 6684 4997 6712
rect 3384 6672 3390 6684
rect 4985 6681 4997 6684
rect 5031 6681 5043 6715
rect 8754 6712 8760 6724
rect 8715 6684 8760 6712
rect 4985 6675 5043 6681
rect 8754 6672 8760 6684
rect 8812 6672 8818 6724
rect 14182 6672 14188 6724
rect 14240 6712 14246 6724
rect 14369 6715 14427 6721
rect 14369 6712 14381 6715
rect 14240 6684 14381 6712
rect 14240 6672 14246 6684
rect 14369 6681 14381 6684
rect 14415 6681 14427 6715
rect 17604 6712 17632 6811
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 18506 6848 18512 6860
rect 18419 6820 18512 6848
rect 18506 6808 18512 6820
rect 18564 6848 18570 6860
rect 19150 6848 19156 6860
rect 18564 6820 19156 6848
rect 18564 6808 18570 6820
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19242 6808 19248 6860
rect 19300 6848 19306 6860
rect 19346 6848 19374 6879
rect 20824 6860 20852 6888
rect 21085 6885 21097 6888
rect 21131 6885 21143 6919
rect 23934 6916 23940 6928
rect 21085 6879 21143 6885
rect 23400 6888 23940 6916
rect 19610 6848 19616 6860
rect 19300 6820 19616 6848
rect 19300 6808 19306 6820
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 19889 6851 19947 6857
rect 19889 6817 19901 6851
rect 19935 6848 19947 6851
rect 20806 6848 20812 6860
rect 19935 6820 20812 6848
rect 19935 6817 19947 6820
rect 19889 6811 19947 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 22500 6851 22558 6857
rect 22500 6848 22512 6851
rect 22388 6820 22512 6848
rect 18138 6780 18144 6792
rect 18099 6752 18144 6780
rect 18138 6740 18144 6752
rect 18196 6740 18202 6792
rect 18969 6783 19027 6789
rect 18969 6749 18981 6783
rect 19015 6749 19027 6783
rect 20714 6780 20720 6792
rect 20675 6752 20720 6780
rect 18969 6743 19027 6749
rect 18414 6712 18420 6724
rect 17604 6684 18420 6712
rect 14369 6675 14427 6681
rect 18414 6672 18420 6684
rect 18472 6672 18478 6724
rect 18984 6656 19012 6743
rect 20714 6740 20720 6752
rect 20772 6780 20778 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20772 6752 21005 6780
rect 20772 6740 20778 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 21634 6780 21640 6792
rect 21595 6752 21640 6780
rect 20993 6743 21051 6749
rect 21634 6740 21640 6752
rect 21692 6780 21698 6792
rect 22094 6780 22100 6792
rect 21692 6752 22100 6780
rect 21692 6740 21698 6752
rect 22094 6740 22100 6752
rect 22152 6780 22158 6792
rect 22388 6780 22416 6820
rect 22500 6817 22512 6820
rect 22546 6817 22558 6851
rect 22500 6811 22558 6817
rect 22152 6752 22416 6780
rect 22152 6740 22158 6752
rect 21266 6672 21272 6724
rect 21324 6712 21330 6724
rect 21818 6712 21824 6724
rect 21324 6684 21824 6712
rect 21324 6672 21330 6684
rect 21818 6672 21824 6684
rect 21876 6712 21882 6724
rect 23400 6712 23428 6888
rect 23934 6876 23940 6888
rect 23992 6876 23998 6928
rect 24489 6919 24547 6925
rect 24489 6885 24501 6919
rect 24535 6916 24547 6919
rect 25038 6916 25044 6928
rect 24535 6888 25044 6916
rect 24535 6885 24547 6888
rect 24489 6879 24547 6885
rect 25038 6876 25044 6888
rect 25096 6876 25102 6928
rect 27249 6919 27307 6925
rect 27249 6885 27261 6919
rect 27295 6916 27307 6919
rect 27430 6916 27436 6928
rect 27295 6888 27436 6916
rect 27295 6885 27307 6888
rect 27249 6879 27307 6885
rect 27430 6876 27436 6888
rect 27488 6876 27494 6928
rect 27801 6919 27859 6925
rect 27801 6885 27813 6919
rect 27847 6916 27859 6919
rect 28074 6916 28080 6928
rect 27847 6888 28080 6916
rect 27847 6885 27859 6888
rect 27801 6879 27859 6885
rect 28074 6876 28080 6888
rect 28132 6876 28138 6928
rect 28810 6916 28816 6928
rect 28771 6888 28816 6916
rect 28810 6876 28816 6888
rect 28868 6876 28874 6928
rect 32487 6919 32545 6925
rect 30852 6888 31064 6916
rect 24026 6848 24032 6860
rect 23987 6820 24032 6848
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 24305 6851 24363 6857
rect 24305 6817 24317 6851
rect 24351 6817 24363 6851
rect 24305 6811 24363 6817
rect 24320 6780 24348 6811
rect 24854 6808 24860 6860
rect 24912 6848 24918 6860
rect 25314 6848 25320 6860
rect 24912 6820 25320 6848
rect 24912 6808 24918 6820
rect 25314 6808 25320 6820
rect 25372 6808 25378 6860
rect 30374 6848 30380 6860
rect 30335 6820 30380 6848
rect 30374 6808 30380 6820
rect 30432 6808 30438 6860
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 30745 6851 30803 6857
rect 30745 6848 30757 6851
rect 30616 6820 30757 6848
rect 30616 6808 30622 6820
rect 30745 6817 30757 6820
rect 30791 6848 30803 6851
rect 30852 6848 30880 6888
rect 30791 6820 30880 6848
rect 30929 6851 30987 6857
rect 30791 6817 30803 6820
rect 30745 6811 30803 6817
rect 30929 6817 30941 6851
rect 30975 6817 30987 6851
rect 31036 6848 31064 6888
rect 32487 6885 32499 6919
rect 32533 6916 32545 6919
rect 32674 6916 32680 6928
rect 32533 6888 32680 6916
rect 32533 6885 32545 6888
rect 32487 6879 32545 6885
rect 32674 6876 32680 6888
rect 32732 6876 32738 6928
rect 34606 6916 34612 6928
rect 34567 6888 34612 6916
rect 34606 6876 34612 6888
rect 34664 6876 34670 6928
rect 35176 6925 35204 6956
rect 35342 6944 35348 6956
rect 35400 6984 35406 6996
rect 35437 6987 35495 6993
rect 35437 6984 35449 6987
rect 35400 6956 35449 6984
rect 35400 6944 35406 6956
rect 35437 6953 35449 6956
rect 35483 6953 35495 6987
rect 35437 6947 35495 6953
rect 35161 6919 35219 6925
rect 35161 6885 35173 6919
rect 35207 6885 35219 6919
rect 36170 6916 36176 6928
rect 36131 6888 36176 6916
rect 35161 6879 35219 6885
rect 36170 6876 36176 6888
rect 36228 6876 36234 6928
rect 31570 6848 31576 6860
rect 31036 6820 31576 6848
rect 30929 6811 30987 6817
rect 24320 6752 24992 6780
rect 24964 6724 24992 6752
rect 26326 6740 26332 6792
rect 26384 6780 26390 6792
rect 27157 6783 27215 6789
rect 27157 6780 27169 6783
rect 26384 6752 27169 6780
rect 26384 6740 26390 6752
rect 27157 6749 27169 6752
rect 27203 6749 27215 6783
rect 27157 6743 27215 6749
rect 28537 6783 28595 6789
rect 28537 6749 28549 6783
rect 28583 6780 28595 6783
rect 28721 6783 28779 6789
rect 28721 6780 28733 6783
rect 28583 6752 28733 6780
rect 28583 6749 28595 6752
rect 28537 6743 28595 6749
rect 28721 6749 28733 6752
rect 28767 6780 28779 6783
rect 28902 6780 28908 6792
rect 28767 6752 28908 6780
rect 28767 6749 28779 6752
rect 28721 6743 28779 6749
rect 28902 6740 28908 6752
rect 28960 6740 28966 6792
rect 29086 6780 29092 6792
rect 29047 6752 29092 6780
rect 29086 6740 29092 6752
rect 29144 6740 29150 6792
rect 30392 6780 30420 6808
rect 30944 6780 30972 6811
rect 31570 6808 31576 6820
rect 31628 6808 31634 6860
rect 31110 6780 31116 6792
rect 30392 6752 31116 6780
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 31205 6783 31263 6789
rect 31205 6749 31217 6783
rect 31251 6780 31263 6783
rect 32125 6783 32183 6789
rect 32125 6780 32137 6783
rect 31251 6752 32137 6780
rect 31251 6749 31263 6752
rect 31205 6743 31263 6749
rect 32125 6749 32137 6752
rect 32171 6780 32183 6783
rect 33870 6780 33876 6792
rect 32171 6752 33876 6780
rect 32171 6749 32183 6752
rect 32125 6743 32183 6749
rect 33870 6740 33876 6752
rect 33928 6740 33934 6792
rect 34146 6740 34152 6792
rect 34204 6780 34210 6792
rect 34517 6783 34575 6789
rect 34517 6780 34529 6783
rect 34204 6752 34529 6780
rect 34204 6740 34210 6752
rect 34517 6749 34529 6752
rect 34563 6749 34575 6783
rect 36078 6780 36084 6792
rect 36039 6752 36084 6780
rect 34517 6743 34575 6749
rect 36078 6740 36084 6752
rect 36136 6740 36142 6792
rect 36354 6780 36360 6792
rect 36315 6752 36360 6780
rect 36354 6740 36360 6752
rect 36412 6740 36418 6792
rect 21876 6684 23428 6712
rect 21876 6672 21882 6684
rect 24946 6672 24952 6724
rect 25004 6712 25010 6724
rect 25501 6715 25559 6721
rect 25501 6712 25513 6715
rect 25004 6684 25513 6712
rect 25004 6672 25010 6684
rect 25501 6681 25513 6684
rect 25547 6712 25559 6715
rect 26050 6712 26056 6724
rect 25547 6684 26056 6712
rect 25547 6681 25559 6684
rect 25501 6675 25559 6681
rect 26050 6672 26056 6684
rect 26108 6672 26114 6724
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3145 6647 3203 6653
rect 3145 6644 3157 6647
rect 2832 6616 3157 6644
rect 2832 6604 2838 6616
rect 3145 6613 3157 6616
rect 3191 6613 3203 6647
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3145 6607 3203 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 7064 6616 7481 6644
rect 7064 6604 7070 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8018 6644 8024 6656
rect 7975 6616 8024 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8018 6604 8024 6616
rect 8076 6644 8082 6656
rect 8478 6644 8484 6656
rect 8076 6616 8484 6644
rect 8076 6604 8082 6616
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 9030 6644 9036 6656
rect 8991 6616 9036 6644
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 12894 6644 12900 6656
rect 12855 6616 12900 6644
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13998 6644 14004 6656
rect 13959 6616 14004 6644
rect 13998 6604 14004 6616
rect 14056 6604 14062 6656
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 18966 6644 18972 6656
rect 18923 6616 18972 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 21542 6604 21548 6656
rect 21600 6644 21606 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 21600 6616 22293 6644
rect 21600 6604 21606 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 22603 6647 22661 6653
rect 22603 6613 22615 6647
rect 22649 6644 22661 6647
rect 23382 6644 23388 6656
rect 22649 6616 23388 6644
rect 22649 6613 22661 6616
rect 22603 6607 22661 6613
rect 23382 6604 23388 6616
rect 23440 6604 23446 6656
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 26510 6644 26516 6656
rect 26292 6616 26516 6644
rect 26292 6604 26298 6616
rect 26510 6604 26516 6616
rect 26568 6644 26574 6656
rect 26697 6647 26755 6653
rect 26697 6644 26709 6647
rect 26568 6616 26709 6644
rect 26568 6604 26574 6616
rect 26697 6613 26709 6616
rect 26743 6613 26755 6647
rect 33042 6644 33048 6656
rect 33003 6616 33048 6644
rect 26697 6607 26755 6613
rect 33042 6604 33048 6616
rect 33100 6604 33106 6656
rect 33502 6644 33508 6656
rect 33463 6616 33508 6644
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2222 6440 2228 6452
rect 2087 6412 2228 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6403
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 4154 6440 4160 6452
rect 4115 6412 4160 6440
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 5258 6440 5264 6452
rect 5219 6412 5264 6440
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 5592 6412 6561 6440
rect 5592 6400 5598 6412
rect 6549 6409 6561 6412
rect 6595 6440 6607 6443
rect 6638 6440 6644 6452
rect 6595 6412 6644 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 12066 6440 12072 6452
rect 12027 6412 12072 6440
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13722 6440 13728 6452
rect 13403 6412 13728 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13722 6400 13728 6412
rect 13780 6440 13786 6452
rect 13998 6440 14004 6452
rect 13780 6412 14004 6440
rect 13780 6400 13786 6412
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 16574 6440 16580 6452
rect 16535 6412 16580 6440
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16908 6412 16957 6440
rect 16908 6400 16914 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 16945 6403 17003 6409
rect 17681 6443 17739 6449
rect 17681 6409 17693 6443
rect 17727 6440 17739 6443
rect 17770 6440 17776 6452
rect 17727 6412 17776 6440
rect 17727 6409 17739 6412
rect 17681 6403 17739 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21177 6443 21235 6449
rect 21177 6440 21189 6443
rect 20864 6412 21189 6440
rect 20864 6400 20870 6412
rect 21177 6409 21189 6412
rect 21223 6409 21235 6443
rect 21818 6440 21824 6452
rect 21779 6412 21824 6440
rect 21177 6403 21235 6409
rect 21818 6400 21824 6412
rect 21876 6400 21882 6452
rect 23106 6440 23112 6452
rect 23019 6412 23112 6440
rect 23106 6400 23112 6412
rect 23164 6440 23170 6452
rect 24026 6440 24032 6452
rect 23164 6412 24032 6440
rect 23164 6400 23170 6412
rect 24026 6400 24032 6412
rect 24084 6400 24090 6452
rect 24946 6440 24952 6452
rect 24907 6412 24952 6440
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 25314 6440 25320 6452
rect 25275 6412 25320 6440
rect 25314 6400 25320 6412
rect 25372 6400 25378 6452
rect 27157 6443 27215 6449
rect 27157 6409 27169 6443
rect 27203 6440 27215 6443
rect 27430 6440 27436 6452
rect 27203 6412 27436 6440
rect 27203 6409 27215 6412
rect 27157 6403 27215 6409
rect 27430 6400 27436 6412
rect 27488 6400 27494 6452
rect 28721 6443 28779 6449
rect 28721 6409 28733 6443
rect 28767 6440 28779 6443
rect 28810 6440 28816 6452
rect 28767 6412 28816 6440
rect 28767 6409 28779 6412
rect 28721 6403 28779 6409
rect 28810 6400 28816 6412
rect 28868 6400 28874 6452
rect 30558 6440 30564 6452
rect 30519 6412 30564 6440
rect 30558 6400 30564 6412
rect 30616 6400 30622 6452
rect 32217 6443 32275 6449
rect 32217 6409 32229 6443
rect 32263 6440 32275 6443
rect 32493 6443 32551 6449
rect 32493 6440 32505 6443
rect 32263 6412 32505 6440
rect 32263 6409 32275 6412
rect 32217 6403 32275 6409
rect 32493 6409 32505 6412
rect 32539 6440 32551 6443
rect 32674 6440 32680 6452
rect 32539 6412 32680 6440
rect 32539 6409 32551 6412
rect 32493 6403 32551 6409
rect 32674 6400 32680 6412
rect 32732 6400 32738 6452
rect 33870 6440 33876 6452
rect 33831 6412 33876 6440
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 36078 6400 36084 6452
rect 36136 6440 36142 6452
rect 36446 6440 36452 6452
rect 36136 6412 36452 6440
rect 36136 6400 36142 6412
rect 36446 6400 36452 6412
rect 36504 6440 36510 6452
rect 36587 6443 36645 6449
rect 36587 6440 36599 6443
rect 36504 6412 36599 6440
rect 36504 6400 36510 6412
rect 36587 6409 36599 6412
rect 36633 6409 36645 6443
rect 36587 6403 36645 6409
rect 3326 6372 3332 6384
rect 3287 6344 3332 6372
rect 3326 6332 3332 6344
rect 3384 6332 3390 6384
rect 24578 6372 24584 6384
rect 24539 6344 24584 6372
rect 24578 6332 24584 6344
rect 24636 6332 24642 6384
rect 28074 6372 28080 6384
rect 27724 6344 28080 6372
rect 2498 6264 2504 6316
rect 2556 6304 2562 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2556 6276 2789 6304
rect 2556 6264 2562 6276
rect 2777 6273 2789 6276
rect 2823 6304 2835 6307
rect 3418 6304 3424 6316
rect 2823 6276 3424 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4614 6304 4620 6316
rect 4575 6276 4620 6304
rect 4614 6264 4620 6276
rect 4672 6264 4678 6316
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7006 6304 7012 6316
rect 6319 6276 7012 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 9030 6304 9036 6316
rect 7607 6276 9036 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 11054 6304 11060 6316
rect 11015 6276 11060 6304
rect 11054 6264 11060 6276
rect 11112 6264 11118 6316
rect 18506 6304 18512 6316
rect 18467 6276 18512 6304
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 18690 6264 18696 6316
rect 18748 6304 18754 6316
rect 27724 6313 27752 6344
rect 28074 6332 28080 6344
rect 28132 6332 28138 6384
rect 18785 6307 18843 6313
rect 18785 6304 18797 6307
rect 18748 6276 18797 6304
rect 18748 6264 18754 6276
rect 18785 6273 18797 6276
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 27709 6307 27767 6313
rect 27709 6273 27721 6307
rect 27755 6273 27767 6307
rect 27982 6304 27988 6316
rect 27943 6276 27988 6304
rect 27709 6267 27767 6273
rect 27982 6264 27988 6276
rect 28040 6264 28046 6316
rect 29086 6264 29092 6316
rect 29144 6304 29150 6316
rect 29641 6307 29699 6313
rect 29641 6304 29653 6307
rect 29144 6276 29653 6304
rect 29144 6264 29150 6276
rect 29641 6273 29653 6276
rect 29687 6273 29699 6307
rect 29641 6267 29699 6273
rect 31110 6264 31116 6316
rect 31168 6304 31174 6316
rect 32692 6304 32720 6400
rect 33042 6332 33048 6384
rect 33100 6372 33106 6384
rect 34241 6375 34299 6381
rect 34241 6372 34253 6375
rect 33100 6344 34253 6372
rect 33100 6332 33106 6344
rect 34241 6341 34253 6344
rect 34287 6372 34299 6375
rect 34606 6372 34612 6384
rect 34287 6344 34612 6372
rect 34287 6341 34299 6344
rect 34241 6335 34299 6341
rect 34606 6332 34612 6344
rect 34664 6372 34670 6384
rect 35989 6375 36047 6381
rect 35989 6372 36001 6375
rect 34664 6344 36001 6372
rect 34664 6332 34670 6344
rect 35989 6341 36001 6344
rect 36035 6372 36047 6375
rect 36170 6372 36176 6384
rect 36035 6344 36176 6372
rect 36035 6341 36047 6344
rect 35989 6335 36047 6341
rect 36170 6332 36176 6344
rect 36228 6332 36234 6384
rect 35342 6304 35348 6316
rect 31168 6276 31616 6304
rect 32692 6276 32812 6304
rect 35303 6276 35348 6304
rect 31168 6264 31174 6276
rect 8662 6236 8668 6248
rect 1443 6208 2084 6236
rect 8623 6208 8668 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 8849 6239 8907 6245
rect 8849 6205 8861 6239
rect 8895 6205 8907 6239
rect 8849 6199 8907 6205
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6236 12495 6239
rect 12986 6236 12992 6248
rect 12483 6208 12992 6236
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 2314 6168 2320 6180
rect 1728 6140 2320 6168
rect 1728 6128 1734 6140
rect 2314 6128 2320 6140
rect 2372 6128 2378 6180
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3142 6168 3148 6180
rect 2915 6140 3148 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6137 4491 6171
rect 4433 6131 4491 6137
rect 2774 6060 2780 6112
rect 2832 6100 2838 6112
rect 3697 6103 3755 6109
rect 3697 6100 3709 6103
rect 2832 6072 3709 6100
rect 2832 6060 2838 6072
rect 3697 6069 3709 6072
rect 3743 6100 3755 6103
rect 4448 6100 4476 6131
rect 4614 6128 4620 6180
rect 4672 6168 4678 6180
rect 6917 6171 6975 6177
rect 6917 6168 6929 6171
rect 4672 6140 6929 6168
rect 4672 6128 4678 6140
rect 6917 6137 6929 6140
rect 6963 6137 6975 6171
rect 6917 6131 6975 6137
rect 3743 6072 4476 6100
rect 6932 6100 6960 6131
rect 7006 6128 7012 6180
rect 7064 6168 7070 6180
rect 7064 6140 7109 6168
rect 7064 6128 7070 6140
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 8864 6168 8892 6199
rect 12986 6196 12992 6208
rect 13044 6236 13050 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13044 6208 13645 6236
rect 13044 6196 13050 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13633 6199 13691 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14182 6236 14188 6248
rect 14139 6208 14188 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14182 6196 14188 6208
rect 14240 6196 14246 6248
rect 15378 6236 15384 6248
rect 15339 6208 15384 6236
rect 15378 6196 15384 6208
rect 15436 6196 15442 6248
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6236 20039 6239
rect 20162 6236 20168 6248
rect 20027 6208 20168 6236
rect 20027 6205 20039 6208
rect 19981 6199 20039 6205
rect 20162 6196 20168 6208
rect 20220 6196 20226 6248
rect 21818 6196 21824 6248
rect 21876 6236 21882 6248
rect 22005 6239 22063 6245
rect 22005 6236 22017 6239
rect 21876 6208 22017 6236
rect 21876 6196 21882 6208
rect 22005 6205 22017 6208
rect 22051 6205 22063 6239
rect 22554 6236 22560 6248
rect 22515 6208 22560 6236
rect 22005 6199 22063 6205
rect 22554 6196 22560 6208
rect 22612 6196 22618 6248
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6196 23722 6248
rect 25866 6236 25872 6248
rect 25827 6208 25872 6236
rect 25866 6196 25872 6208
rect 25924 6196 25930 6248
rect 31021 6239 31079 6245
rect 31021 6205 31033 6239
rect 31067 6236 31079 6239
rect 31386 6236 31392 6248
rect 31067 6208 31392 6236
rect 31067 6205 31079 6208
rect 31021 6199 31079 6205
rect 31386 6196 31392 6208
rect 31444 6196 31450 6248
rect 31588 6245 31616 6276
rect 31573 6239 31631 6245
rect 31573 6205 31585 6239
rect 31619 6205 31631 6239
rect 31573 6199 31631 6205
rect 31849 6239 31907 6245
rect 31849 6205 31861 6239
rect 31895 6236 31907 6239
rect 32674 6236 32680 6248
rect 31895 6208 32680 6236
rect 31895 6205 31907 6208
rect 31849 6199 31907 6205
rect 32674 6196 32680 6208
rect 32732 6196 32738 6248
rect 10778 6168 10784 6180
rect 8352 6140 8892 6168
rect 10739 6140 10784 6168
rect 8352 6128 8358 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 10928 6140 10973 6168
rect 10928 6128 10934 6140
rect 12066 6128 12072 6180
rect 12124 6168 12130 6180
rect 12799 6171 12857 6177
rect 12799 6168 12811 6171
rect 12124 6140 12811 6168
rect 12124 6128 12130 6140
rect 12799 6137 12811 6140
rect 12845 6168 12857 6171
rect 13170 6168 13176 6180
rect 12845 6140 13176 6168
rect 12845 6137 12857 6140
rect 12799 6131 12857 6137
rect 13170 6128 13176 6140
rect 13228 6168 13234 6180
rect 15746 6177 15752 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 13228 6140 15301 6168
rect 13228 6128 13234 6140
rect 15289 6137 15301 6140
rect 15335 6168 15347 6171
rect 15743 6168 15752 6177
rect 15335 6140 15752 6168
rect 15335 6137 15347 6140
rect 15289 6131 15347 6137
rect 15743 6131 15752 6140
rect 15746 6128 15752 6131
rect 15804 6128 15810 6180
rect 18598 6168 18604 6180
rect 18559 6140 18604 6168
rect 18598 6128 18604 6140
rect 18656 6128 18662 6180
rect 19521 6171 19579 6177
rect 19521 6137 19533 6171
rect 19567 6168 19579 6171
rect 19610 6168 19616 6180
rect 19567 6140 19616 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 19610 6128 19616 6140
rect 19668 6168 19674 6180
rect 19889 6171 19947 6177
rect 19889 6168 19901 6171
rect 19668 6140 19901 6168
rect 19668 6128 19674 6140
rect 19889 6137 19901 6140
rect 19935 6168 19947 6171
rect 20343 6171 20401 6177
rect 20343 6168 20355 6171
rect 19935 6140 20355 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20343 6137 20355 6140
rect 20389 6168 20401 6171
rect 21358 6168 21364 6180
rect 20389 6140 21364 6168
rect 20389 6137 20401 6140
rect 20343 6131 20401 6137
rect 21358 6128 21364 6140
rect 21416 6128 21422 6180
rect 23982 6171 24040 6177
rect 23982 6137 23994 6171
rect 24028 6168 24040 6171
rect 26190 6171 26248 6177
rect 26190 6168 26202 6171
rect 24028 6140 24062 6168
rect 25700 6140 26202 6168
rect 24028 6137 24040 6140
rect 23982 6131 24040 6137
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 6932 6072 7849 6100
rect 3743 6069 3755 6072
rect 3697 6063 3755 6069
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 8478 6100 8484 6112
rect 8439 6072 8484 6100
rect 7837 6063 7895 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9766 6100 9772 6112
rect 9727 6072 9772 6100
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10226 6100 10232 6112
rect 10183 6072 10232 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10597 6103 10655 6109
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 10888 6100 10916 6128
rect 10643 6072 10916 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 14182 6060 14188 6112
rect 14240 6100 14246 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 14240 6072 14381 6100
rect 14240 6060 14246 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14369 6063 14427 6069
rect 14737 6103 14795 6109
rect 14737 6069 14749 6103
rect 14783 6100 14795 6103
rect 15010 6100 15016 6112
rect 14783 6072 15016 6100
rect 14783 6069 14795 6072
rect 14737 6063 14795 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 18325 6103 18383 6109
rect 18325 6069 18337 6103
rect 18371 6100 18383 6103
rect 18414 6100 18420 6112
rect 18371 6072 18420 6100
rect 18371 6069 18383 6072
rect 18325 6063 18383 6069
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20772 6072 20913 6100
rect 20772 6060 20778 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 22278 6100 22284 6112
rect 22239 6072 22284 6100
rect 20901 6063 20959 6069
rect 22278 6060 22284 6072
rect 22336 6060 22342 6112
rect 23382 6100 23388 6112
rect 23343 6072 23388 6100
rect 23382 6060 23388 6072
rect 23440 6100 23446 6112
rect 23997 6100 24025 6131
rect 24670 6100 24676 6112
rect 23440 6072 24676 6100
rect 23440 6060 23446 6072
rect 24670 6060 24676 6072
rect 24728 6100 24734 6112
rect 25700 6109 25728 6140
rect 26190 6137 26202 6140
rect 26236 6137 26248 6171
rect 26190 6131 26248 6137
rect 27801 6171 27859 6177
rect 27801 6137 27813 6171
rect 27847 6168 27859 6171
rect 28810 6168 28816 6180
rect 27847 6140 28816 6168
rect 27847 6137 27859 6140
rect 27801 6131 27859 6137
rect 25685 6103 25743 6109
rect 25685 6100 25697 6103
rect 24728 6072 25697 6100
rect 24728 6060 24734 6072
rect 25685 6069 25697 6072
rect 25731 6069 25743 6103
rect 25685 6063 25743 6069
rect 26789 6103 26847 6109
rect 26789 6069 26801 6103
rect 26835 6100 26847 6103
rect 27525 6103 27583 6109
rect 27525 6100 27537 6103
rect 26835 6072 27537 6100
rect 26835 6069 26847 6072
rect 26789 6063 26847 6069
rect 27525 6069 27537 6072
rect 27571 6100 27583 6103
rect 27816 6100 27844 6131
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 29362 6168 29368 6180
rect 29323 6140 29368 6168
rect 29362 6128 29368 6140
rect 29420 6128 29426 6180
rect 29457 6171 29515 6177
rect 29457 6137 29469 6171
rect 29503 6137 29515 6171
rect 32784 6168 32812 6276
rect 35342 6264 35348 6276
rect 35400 6264 35406 6316
rect 33597 6239 33655 6245
rect 33597 6205 33609 6239
rect 33643 6236 33655 6239
rect 34606 6236 34612 6248
rect 33643 6208 34612 6236
rect 33643 6205 33655 6208
rect 33597 6199 33655 6205
rect 34606 6196 34612 6208
rect 34664 6196 34670 6248
rect 35894 6196 35900 6248
rect 35952 6236 35958 6248
rect 36484 6239 36542 6245
rect 36484 6236 36496 6239
rect 35952 6208 36496 6236
rect 35952 6196 35958 6208
rect 36484 6205 36496 6208
rect 36530 6236 36542 6239
rect 36909 6239 36967 6245
rect 36909 6236 36921 6239
rect 36530 6208 36921 6236
rect 36530 6205 36542 6208
rect 36484 6199 36542 6205
rect 36909 6205 36921 6208
rect 36955 6205 36967 6239
rect 36909 6199 36967 6205
rect 32998 6171 33056 6177
rect 32998 6168 33010 6171
rect 32784 6140 33010 6168
rect 29457 6131 29515 6137
rect 32998 6137 33010 6140
rect 33044 6137 33056 6171
rect 34974 6168 34980 6180
rect 34935 6140 34980 6168
rect 32998 6131 33056 6137
rect 27571 6072 27844 6100
rect 29089 6103 29147 6109
rect 27571 6069 27583 6072
rect 27525 6063 27583 6069
rect 29089 6069 29101 6103
rect 29135 6100 29147 6103
rect 29178 6100 29184 6112
rect 29135 6072 29184 6100
rect 29135 6069 29147 6072
rect 29089 6063 29147 6069
rect 29178 6060 29184 6072
rect 29236 6100 29242 6112
rect 29472 6100 29500 6131
rect 34974 6128 34980 6140
rect 35032 6128 35038 6180
rect 35069 6171 35127 6177
rect 35069 6137 35081 6171
rect 35115 6137 35127 6171
rect 35069 6131 35127 6137
rect 29236 6072 29500 6100
rect 29236 6060 29242 6072
rect 34606 6060 34612 6112
rect 34664 6100 34670 6112
rect 35084 6100 35112 6131
rect 34664 6072 35112 6100
rect 34664 6060 34670 6072
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 2961 5899 3019 5905
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3142 5896 3148 5908
rect 3007 5868 3148 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4396 5868 5089 5896
rect 4396 5856 4402 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 5077 5859 5135 5865
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 6822 5896 6828 5908
rect 6779 5868 6828 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 6972 5868 7297 5896
rect 6972 5856 6978 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 8662 5896 8668 5908
rect 8527 5868 8668 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 8662 5856 8668 5868
rect 8720 5856 8726 5908
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 9582 5896 9588 5908
rect 9180 5868 9588 5896
rect 9180 5856 9186 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5865 10655 5899
rect 11974 5896 11980 5908
rect 11935 5868 11980 5896
rect 10597 5859 10655 5865
rect 2038 5828 2044 5840
rect 1999 5800 2044 5828
rect 2038 5788 2044 5800
rect 2096 5788 2102 5840
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 5810 5828 5816 5840
rect 4295 5800 5816 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 7098 5828 7104 5840
rect 7011 5800 7104 5828
rect 7098 5788 7104 5800
rect 7156 5828 7162 5840
rect 9490 5828 9496 5840
rect 7156 5800 9496 5828
rect 7156 5788 7162 5800
rect 7484 5769 7512 5800
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9998 5831 10056 5837
rect 9998 5828 10010 5831
rect 9824 5800 10010 5828
rect 9824 5788 9830 5800
rect 9998 5797 10010 5800
rect 10044 5797 10056 5831
rect 10612 5828 10640 5859
rect 11974 5856 11980 5868
rect 12032 5896 12038 5908
rect 12342 5896 12348 5908
rect 12032 5868 12348 5896
rect 12032 5856 12038 5868
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 13170 5896 13176 5908
rect 13131 5868 13176 5896
rect 13170 5856 13176 5868
rect 13228 5856 13234 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13906 5896 13912 5908
rect 13587 5868 13912 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13906 5856 13912 5868
rect 13964 5856 13970 5908
rect 16485 5899 16543 5905
rect 16485 5865 16497 5899
rect 16531 5896 16543 5899
rect 16666 5896 16672 5908
rect 16531 5868 16672 5896
rect 16531 5865 16543 5868
rect 16485 5859 16543 5865
rect 16666 5856 16672 5868
rect 16724 5896 16730 5908
rect 17770 5896 17776 5908
rect 16724 5868 17776 5896
rect 16724 5856 16730 5868
rect 17770 5856 17776 5868
rect 17828 5856 17834 5908
rect 18509 5899 18567 5905
rect 18509 5865 18521 5899
rect 18555 5896 18567 5899
rect 18598 5896 18604 5908
rect 18555 5868 18604 5896
rect 18555 5865 18567 5868
rect 18509 5859 18567 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 19886 5896 19892 5908
rect 19847 5868 19892 5896
rect 19886 5856 19892 5868
rect 19944 5856 19950 5908
rect 22097 5899 22155 5905
rect 22097 5865 22109 5899
rect 22143 5896 22155 5899
rect 22554 5896 22560 5908
rect 22143 5868 22560 5896
rect 22143 5865 22155 5868
rect 22097 5859 22155 5865
rect 22554 5856 22560 5868
rect 22612 5856 22618 5908
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23716 5868 24409 5896
rect 23716 5856 23722 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 26326 5896 26332 5908
rect 26287 5868 26332 5896
rect 24397 5859 24455 5865
rect 26326 5856 26332 5868
rect 26384 5856 26390 5908
rect 31110 5896 31116 5908
rect 31071 5868 31116 5896
rect 31110 5856 31116 5868
rect 31168 5856 31174 5908
rect 32674 5896 32680 5908
rect 32635 5868 32680 5896
rect 32674 5856 32680 5868
rect 32732 5856 32738 5908
rect 33551 5899 33609 5905
rect 33551 5865 33563 5899
rect 33597 5896 33609 5899
rect 34146 5896 34152 5908
rect 33597 5868 34152 5896
rect 33597 5865 33609 5868
rect 33551 5859 33609 5865
rect 34146 5856 34152 5868
rect 34204 5896 34210 5908
rect 34241 5899 34299 5905
rect 34241 5896 34253 5899
rect 34204 5868 34253 5896
rect 34204 5856 34210 5868
rect 34241 5865 34253 5868
rect 34287 5865 34299 5899
rect 34241 5859 34299 5865
rect 34974 5856 34980 5908
rect 35032 5896 35038 5908
rect 35437 5899 35495 5905
rect 35437 5896 35449 5899
rect 35032 5868 35449 5896
rect 35032 5856 35038 5868
rect 35437 5865 35449 5868
rect 35483 5865 35495 5899
rect 36446 5896 36452 5908
rect 36407 5868 36452 5896
rect 35437 5859 35495 5865
rect 36446 5856 36452 5868
rect 36504 5856 36510 5908
rect 12158 5828 12164 5840
rect 10612 5800 12164 5828
rect 9998 5791 10056 5797
rect 12158 5788 12164 5800
rect 12216 5828 12222 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 12216 5800 12265 5828
rect 12216 5788 12222 5800
rect 12253 5797 12265 5800
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 13446 5828 13452 5840
rect 12860 5800 13452 5828
rect 12860 5788 12866 5800
rect 13446 5788 13452 5800
rect 13504 5828 13510 5840
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13504 5800 13737 5828
rect 13504 5788 13510 5800
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 13725 5791 13783 5797
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 14090 5828 14096 5840
rect 13863 5800 14096 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 14090 5788 14096 5800
rect 14148 5828 14154 5840
rect 15473 5831 15531 5837
rect 15473 5828 15485 5831
rect 14148 5800 15485 5828
rect 14148 5788 14154 5800
rect 15473 5797 15485 5800
rect 15519 5797 15531 5831
rect 15473 5791 15531 5797
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 16942 5828 16948 5840
rect 16448 5800 16948 5828
rect 16448 5788 16454 5800
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 17037 5831 17095 5837
rect 17037 5797 17049 5831
rect 17083 5828 17095 5831
rect 18963 5831 19021 5837
rect 17083 5800 18000 5828
rect 17083 5797 17095 5800
rect 17037 5791 17095 5797
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5729 7527 5763
rect 7469 5723 7527 5729
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 8294 5760 8300 5772
rect 7791 5732 8300 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 1949 5695 2007 5701
rect 1949 5661 1961 5695
rect 1995 5692 2007 5695
rect 3513 5695 3571 5701
rect 3513 5692 3525 5695
rect 1995 5664 3525 5692
rect 1995 5661 2007 5664
rect 1949 5655 2007 5661
rect 3513 5661 3525 5664
rect 3559 5661 3571 5695
rect 4154 5692 4160 5704
rect 4115 5664 4160 5692
rect 3513 5655 3571 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4614 5692 4620 5704
rect 4479 5664 4620 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 2501 5627 2559 5633
rect 2501 5593 2513 5627
rect 2547 5624 2559 5627
rect 4448 5624 4476 5655
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5592 5664 5733 5692
rect 5592 5652 5598 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5721 5655 5779 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6822 5652 6828 5704
rect 6880 5692 6886 5704
rect 7760 5692 7788 5723
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 9674 5692 9680 5704
rect 6880 5664 7788 5692
rect 9635 5664 9680 5692
rect 6880 5652 6886 5664
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11940 5664 12173 5692
rect 11940 5652 11946 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 14369 5695 14427 5701
rect 14369 5661 14381 5695
rect 14415 5692 14427 5695
rect 14918 5692 14924 5704
rect 14415 5664 14924 5692
rect 14415 5661 14427 5664
rect 14369 5655 14427 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15381 5695 15439 5701
rect 15381 5692 15393 5695
rect 15252 5664 15393 5692
rect 15252 5652 15258 5664
rect 15381 5661 15393 5664
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 10870 5624 10876 5636
rect 2547 5596 4476 5624
rect 10831 5596 10876 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 12713 5627 12771 5633
rect 12713 5593 12725 5627
rect 12759 5624 12771 5627
rect 13722 5624 13728 5636
rect 12759 5596 13728 5624
rect 12759 5593 12771 5596
rect 12713 5587 12771 5593
rect 13722 5584 13728 5596
rect 13780 5624 13786 5636
rect 15672 5624 15700 5655
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 16816 5664 17233 5692
rect 16816 5652 16822 5664
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17972 5633 18000 5800
rect 18963 5797 18975 5831
rect 19009 5828 19021 5831
rect 19610 5828 19616 5840
rect 19009 5800 19616 5828
rect 19009 5797 19021 5800
rect 18963 5791 19021 5797
rect 19610 5788 19616 5800
rect 19668 5788 19674 5840
rect 20714 5788 20720 5840
rect 20772 5828 20778 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 20772 5800 21097 5828
rect 20772 5788 20778 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21634 5828 21640 5840
rect 21547 5800 21640 5828
rect 21085 5791 21143 5797
rect 21634 5788 21640 5800
rect 21692 5828 21698 5840
rect 22465 5831 22523 5837
rect 22465 5828 22477 5831
rect 21692 5800 22477 5828
rect 21692 5788 21698 5800
rect 22465 5797 22477 5800
rect 22511 5797 22523 5831
rect 22465 5791 22523 5797
rect 23382 5788 23388 5840
rect 23440 5828 23446 5840
rect 23522 5831 23580 5837
rect 23522 5828 23534 5831
rect 23440 5800 23534 5828
rect 23440 5788 23446 5800
rect 23522 5797 23534 5800
rect 23568 5797 23580 5831
rect 27154 5828 27160 5840
rect 27115 5800 27160 5828
rect 23522 5791 23580 5797
rect 27154 5788 27160 5800
rect 27212 5788 27218 5840
rect 27709 5831 27767 5837
rect 27709 5797 27721 5831
rect 27755 5828 27767 5831
rect 27982 5828 27988 5840
rect 27755 5800 27988 5828
rect 27755 5797 27767 5800
rect 27709 5791 27767 5797
rect 27982 5788 27988 5800
rect 28040 5788 28046 5840
rect 28626 5788 28632 5840
rect 28684 5828 28690 5840
rect 28721 5831 28779 5837
rect 28721 5828 28733 5831
rect 28684 5800 28733 5828
rect 28684 5788 28690 5800
rect 28721 5797 28733 5800
rect 28767 5797 28779 5831
rect 30834 5828 30840 5840
rect 30795 5800 30840 5828
rect 28721 5791 28779 5797
rect 30834 5788 30840 5800
rect 30892 5788 30898 5840
rect 18322 5720 18328 5772
rect 18380 5760 18386 5772
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18380 5732 18613 5760
rect 18380 5720 18386 5732
rect 18601 5729 18613 5732
rect 18647 5760 18659 5763
rect 19242 5760 19248 5772
rect 18647 5732 19248 5760
rect 18647 5729 18659 5732
rect 18601 5723 18659 5729
rect 19242 5720 19248 5732
rect 19300 5720 19306 5772
rect 24854 5720 24860 5772
rect 24912 5760 24918 5772
rect 24949 5763 25007 5769
rect 24949 5760 24961 5763
rect 24912 5732 24961 5760
rect 24912 5720 24918 5732
rect 24949 5729 24961 5732
rect 24995 5729 25007 5763
rect 25130 5760 25136 5772
rect 25091 5732 25136 5760
rect 24949 5723 25007 5729
rect 25130 5720 25136 5732
rect 25188 5720 25194 5772
rect 29270 5720 29276 5772
rect 29328 5760 29334 5772
rect 30098 5760 30104 5772
rect 29328 5732 30104 5760
rect 29328 5720 29334 5732
rect 30098 5720 30104 5732
rect 30156 5720 30162 5772
rect 30374 5720 30380 5772
rect 30432 5760 30438 5772
rect 30653 5763 30711 5769
rect 30653 5760 30665 5763
rect 30432 5732 30665 5760
rect 30432 5720 30438 5732
rect 30653 5729 30665 5732
rect 30699 5760 30711 5763
rect 31128 5760 31156 5856
rect 34606 5828 34612 5840
rect 34567 5800 34612 5828
rect 34606 5788 34612 5800
rect 34664 5788 34670 5840
rect 34698 5788 34704 5840
rect 34756 5828 34762 5840
rect 35161 5831 35219 5837
rect 35161 5828 35173 5831
rect 34756 5800 35173 5828
rect 34756 5788 34762 5800
rect 35161 5797 35173 5800
rect 35207 5828 35219 5831
rect 36354 5828 36360 5840
rect 35207 5800 36360 5828
rect 35207 5797 35219 5800
rect 35161 5791 35219 5797
rect 36354 5788 36360 5800
rect 36412 5788 36418 5840
rect 32214 5769 32220 5772
rect 30699 5732 31156 5760
rect 32192 5763 32220 5769
rect 30699 5729 30711 5732
rect 30653 5723 30711 5729
rect 32192 5729 32204 5763
rect 32192 5723 32220 5729
rect 32214 5720 32220 5723
rect 32272 5720 32278 5772
rect 33410 5720 33416 5772
rect 33468 5769 33474 5772
rect 33468 5763 33506 5769
rect 33494 5729 33506 5763
rect 33468 5723 33506 5729
rect 33468 5720 33474 5723
rect 35986 5720 35992 5772
rect 36044 5769 36050 5772
rect 36044 5763 36082 5769
rect 36070 5729 36082 5763
rect 36044 5723 36082 5729
rect 36044 5720 36050 5723
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20864 5664 21005 5692
rect 20864 5652 20870 5664
rect 20993 5661 21005 5664
rect 21039 5661 21051 5695
rect 20993 5655 21051 5661
rect 22278 5652 22284 5704
rect 22336 5692 22342 5704
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22336 5664 23213 5692
rect 22336 5652 22342 5664
rect 23201 5661 23213 5664
rect 23247 5661 23259 5695
rect 25498 5692 25504 5704
rect 25459 5664 25504 5692
rect 23201 5655 23259 5661
rect 25498 5652 25504 5664
rect 25556 5652 25562 5704
rect 26881 5695 26939 5701
rect 26881 5661 26893 5695
rect 26927 5692 26939 5695
rect 27062 5692 27068 5704
rect 26927 5664 27068 5692
rect 26927 5661 26939 5664
rect 26881 5655 26939 5661
rect 27062 5652 27068 5664
rect 27120 5652 27126 5704
rect 28629 5695 28687 5701
rect 28629 5661 28641 5695
rect 28675 5692 28687 5695
rect 28902 5692 28908 5704
rect 28675 5664 28908 5692
rect 28675 5661 28687 5664
rect 28629 5655 28687 5661
rect 28902 5652 28908 5664
rect 28960 5652 28966 5704
rect 29086 5692 29092 5704
rect 29047 5664 29092 5692
rect 29086 5652 29092 5664
rect 29144 5652 29150 5704
rect 34146 5652 34152 5704
rect 34204 5692 34210 5704
rect 34517 5695 34575 5701
rect 34517 5692 34529 5695
rect 34204 5664 34529 5692
rect 34204 5652 34210 5664
rect 34517 5661 34529 5664
rect 34563 5692 34575 5695
rect 36127 5695 36185 5701
rect 36127 5692 36139 5695
rect 34563 5664 36139 5692
rect 34563 5661 34575 5664
rect 34517 5655 34575 5661
rect 36127 5661 36139 5664
rect 36173 5661 36185 5695
rect 36127 5655 36185 5661
rect 13780 5596 15700 5624
rect 17957 5627 18015 5633
rect 13780 5584 13786 5596
rect 17957 5593 17969 5627
rect 18003 5624 18015 5627
rect 19521 5627 19579 5633
rect 19521 5624 19533 5627
rect 18003 5596 19533 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 19521 5593 19533 5596
rect 19567 5593 19579 5627
rect 24118 5624 24124 5636
rect 24079 5596 24124 5624
rect 19521 5587 19579 5593
rect 24118 5584 24124 5596
rect 24176 5584 24182 5636
rect 29362 5584 29368 5636
rect 29420 5624 29426 5636
rect 29641 5627 29699 5633
rect 29641 5624 29653 5627
rect 29420 5596 29653 5624
rect 29420 5584 29426 5596
rect 29641 5593 29653 5596
rect 29687 5624 29699 5627
rect 32263 5627 32321 5633
rect 32263 5624 32275 5627
rect 29687 5596 32275 5624
rect 29687 5593 29699 5596
rect 29641 5587 29699 5593
rect 32263 5593 32275 5596
rect 32309 5593 32321 5627
rect 32263 5587 32321 5593
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 3237 5559 3295 5565
rect 3237 5556 3249 5559
rect 2648 5528 3249 5556
rect 2648 5516 2654 5528
rect 3237 5525 3249 5528
rect 3283 5525 3295 5559
rect 3237 5519 3295 5525
rect 3513 5559 3571 5565
rect 3513 5525 3525 5559
rect 3559 5556 3571 5559
rect 3697 5559 3755 5565
rect 3697 5556 3709 5559
rect 3559 5528 3709 5556
rect 3559 5525 3571 5528
rect 3513 5519 3571 5525
rect 3697 5525 3709 5528
rect 3743 5556 3755 5559
rect 4338 5556 4344 5568
rect 3743 5528 4344 5556
rect 3743 5525 3755 5528
rect 3697 5519 3755 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 8754 5556 8760 5568
rect 8715 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5556 15163 5559
rect 15378 5556 15384 5568
rect 15151 5528 15384 5556
rect 15151 5525 15163 5528
rect 15105 5519 15163 5525
rect 15378 5516 15384 5528
rect 15436 5556 15442 5568
rect 16482 5556 16488 5568
rect 15436 5528 16488 5556
rect 15436 5516 15442 5528
rect 16482 5516 16488 5528
rect 16540 5516 16546 5568
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 19334 5556 19340 5568
rect 18196 5528 19340 5556
rect 18196 5516 18202 5528
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 20162 5556 20168 5568
rect 20123 5528 20168 5556
rect 20162 5516 20168 5528
rect 20220 5516 20226 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 21726 5556 21732 5568
rect 20763 5528 21732 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 21726 5516 21732 5528
rect 21784 5516 21790 5568
rect 25866 5556 25872 5568
rect 25827 5528 25872 5556
rect 25866 5516 25872 5528
rect 25924 5516 25930 5568
rect 28074 5556 28080 5568
rect 27987 5528 28080 5556
rect 28074 5516 28080 5528
rect 28132 5556 28138 5568
rect 29086 5556 29092 5568
rect 28132 5528 29092 5556
rect 28132 5516 28138 5528
rect 29086 5516 29092 5528
rect 29144 5516 29150 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2096 5324 2513 5352
rect 2096 5312 2102 5324
rect 2501 5321 2513 5324
rect 2547 5321 2559 5355
rect 2501 5315 2559 5321
rect 4617 5355 4675 5361
rect 4617 5321 4629 5355
rect 4663 5352 4675 5355
rect 4985 5355 5043 5361
rect 4985 5352 4997 5355
rect 4663 5324 4997 5352
rect 4663 5321 4675 5324
rect 4617 5315 4675 5321
rect 4985 5321 4997 5324
rect 5031 5352 5043 5355
rect 5629 5355 5687 5361
rect 5629 5352 5641 5355
rect 5031 5324 5641 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5629 5321 5641 5324
rect 5675 5352 5687 5355
rect 5810 5352 5816 5364
rect 5675 5324 5816 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 6638 5352 6644 5364
rect 5960 5324 6005 5352
rect 6551 5324 6644 5352
rect 5960 5312 5966 5324
rect 6638 5312 6644 5324
rect 6696 5352 6702 5364
rect 6822 5352 6828 5364
rect 6696 5324 6828 5352
rect 6696 5312 6702 5324
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7282 5352 7288 5364
rect 7243 5324 7288 5352
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 9122 5352 9128 5364
rect 9083 5324 9128 5352
rect 9122 5312 9128 5324
rect 9180 5312 9186 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 9824 5324 10425 5352
rect 9824 5312 9830 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 12158 5352 12164 5364
rect 12119 5324 12164 5352
rect 10413 5315 10471 5321
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 8021 5287 8079 5293
rect 8021 5284 8033 5287
rect 7248 5256 8033 5284
rect 7248 5244 7254 5256
rect 8021 5253 8033 5256
rect 8067 5253 8079 5287
rect 8021 5247 8079 5253
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5148 1639 5151
rect 1762 5148 1768 5160
rect 1627 5120 1768 5148
rect 1627 5117 1639 5120
rect 1581 5111 1639 5117
rect 1762 5108 1768 5120
rect 1820 5148 1826 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 1820 5120 2789 5148
rect 1820 5108 1826 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 3694 5148 3700 5160
rect 3655 5120 3700 5148
rect 2777 5111 2835 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 4154 5148 4160 5160
rect 3896 5120 4160 5148
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 1902 5083 1960 5089
rect 1902 5080 1914 5083
rect 1728 5052 1914 5080
rect 1728 5040 1734 5052
rect 1902 5049 1914 5052
rect 1948 5049 1960 5083
rect 3896 5080 3924 5120
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 5721 5151 5779 5157
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5767 5120 6316 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 6288 5089 6316 5120
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 7101 5151 7159 5157
rect 7101 5148 7113 5151
rect 6420 5120 7113 5148
rect 6420 5108 6426 5120
rect 7101 5117 7113 5120
rect 7147 5148 7159 5151
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7147 5120 7573 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 1902 5043 1960 5049
rect 3252 5052 3924 5080
rect 4059 5083 4117 5089
rect 3252 5024 3280 5052
rect 4059 5049 4071 5083
rect 4105 5049 4117 5083
rect 4059 5043 4117 5049
rect 6273 5083 6331 5089
rect 6273 5049 6285 5083
rect 6319 5080 6331 5083
rect 6822 5080 6828 5092
rect 6319 5052 6828 5080
rect 6319 5049 6331 5052
rect 6273 5043 6331 5049
rect 3234 5012 3240 5024
rect 3195 4984 3240 5012
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3602 5012 3608 5024
rect 3515 4984 3608 5012
rect 3602 4972 3608 4984
rect 3660 5012 3666 5024
rect 4080 5012 4108 5043
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 8036 5080 8064 5247
rect 10428 5216 10456 5315
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 14090 5352 14096 5364
rect 14051 5324 14096 5352
rect 14090 5312 14096 5324
rect 14148 5352 14154 5364
rect 14461 5355 14519 5361
rect 14461 5352 14473 5355
rect 14148 5324 14473 5352
rect 14148 5312 14154 5324
rect 14461 5321 14473 5324
rect 14507 5321 14519 5355
rect 14461 5315 14519 5321
rect 17313 5355 17371 5361
rect 17313 5321 17325 5355
rect 17359 5352 17371 5355
rect 17770 5352 17776 5364
rect 17359 5324 17776 5352
rect 17359 5321 17371 5324
rect 17313 5315 17371 5321
rect 17770 5312 17776 5324
rect 17828 5352 17834 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17828 5324 18337 5352
rect 17828 5312 17834 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 19337 5355 19395 5361
rect 19337 5321 19349 5355
rect 19383 5352 19395 5355
rect 19610 5352 19616 5364
rect 19383 5324 19616 5352
rect 19383 5321 19395 5324
rect 19337 5315 19395 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 20530 5352 20536 5364
rect 20491 5324 20536 5352
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 20806 5312 20812 5364
rect 20864 5352 20870 5364
rect 20901 5355 20959 5361
rect 20901 5352 20913 5355
rect 20864 5324 20913 5352
rect 20864 5312 20870 5324
rect 20901 5321 20913 5324
rect 20947 5321 20959 5355
rect 20901 5315 20959 5321
rect 22278 5312 22284 5364
rect 22336 5352 22342 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22336 5324 22477 5352
rect 22336 5312 22342 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 24762 5352 24768 5364
rect 23532 5324 24768 5352
rect 23532 5312 23538 5324
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 25133 5355 25191 5361
rect 25133 5321 25145 5355
rect 25179 5352 25191 5355
rect 25222 5352 25228 5364
rect 25179 5324 25228 5352
rect 25179 5321 25191 5324
rect 25133 5315 25191 5321
rect 25222 5312 25228 5324
rect 25280 5312 25286 5364
rect 26050 5312 26056 5364
rect 26108 5352 26114 5364
rect 26237 5355 26295 5361
rect 26237 5352 26249 5355
rect 26108 5324 26249 5352
rect 26108 5312 26114 5324
rect 26237 5321 26249 5324
rect 26283 5321 26295 5355
rect 26878 5352 26884 5364
rect 26839 5324 26884 5352
rect 26237 5315 26295 5321
rect 26878 5312 26884 5324
rect 26936 5352 26942 5364
rect 27246 5352 27252 5364
rect 26936 5324 27252 5352
rect 26936 5312 26942 5324
rect 27246 5312 27252 5324
rect 27304 5312 27310 5364
rect 28994 5312 29000 5364
rect 29052 5352 29058 5364
rect 29411 5355 29469 5361
rect 29411 5352 29423 5355
rect 29052 5324 29423 5352
rect 29052 5312 29058 5324
rect 29411 5321 29423 5324
rect 29457 5321 29469 5355
rect 29730 5352 29736 5364
rect 29691 5324 29736 5352
rect 29411 5315 29469 5321
rect 29730 5312 29736 5324
rect 29788 5312 29794 5364
rect 30098 5352 30104 5364
rect 30059 5324 30104 5352
rect 30098 5312 30104 5324
rect 30156 5312 30162 5364
rect 30374 5312 30380 5364
rect 30432 5361 30438 5364
rect 30432 5355 30481 5361
rect 30432 5321 30435 5355
rect 30469 5321 30481 5355
rect 32214 5352 32220 5364
rect 32175 5324 32220 5352
rect 30432 5315 30481 5321
rect 30432 5312 30438 5315
rect 32214 5312 32220 5324
rect 32272 5312 32278 5364
rect 33410 5352 33416 5364
rect 33371 5324 33416 5352
rect 33410 5312 33416 5324
rect 33468 5312 33474 5364
rect 34146 5352 34152 5364
rect 34107 5324 34152 5352
rect 34146 5312 34152 5324
rect 34204 5312 34210 5364
rect 34517 5355 34575 5361
rect 34517 5321 34529 5355
rect 34563 5352 34575 5355
rect 34606 5352 34612 5364
rect 34563 5324 34612 5352
rect 34563 5321 34575 5324
rect 34517 5315 34575 5321
rect 34606 5312 34612 5324
rect 34664 5312 34670 5364
rect 34974 5312 34980 5364
rect 35032 5361 35038 5364
rect 35032 5355 35081 5361
rect 35032 5321 35035 5355
rect 35069 5321 35081 5355
rect 35032 5315 35081 5321
rect 35032 5312 35038 5315
rect 13722 5284 13728 5296
rect 13683 5256 13728 5284
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 30561 5287 30619 5293
rect 30561 5253 30573 5287
rect 30607 5284 30619 5287
rect 30837 5287 30895 5293
rect 30837 5284 30849 5287
rect 30607 5256 30849 5284
rect 30607 5253 30619 5256
rect 30561 5247 30619 5253
rect 30837 5253 30849 5256
rect 30883 5284 30895 5287
rect 32766 5284 32772 5296
rect 30883 5256 32772 5284
rect 30883 5253 30895 5256
rect 30837 5247 30895 5253
rect 32766 5244 32772 5256
rect 32824 5244 32830 5296
rect 10428 5188 10732 5216
rect 8202 5148 8208 5160
rect 8163 5120 8208 5148
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10060 5120 10609 5148
rect 8526 5083 8584 5089
rect 8526 5080 8538 5083
rect 8036 5052 8538 5080
rect 8526 5049 8538 5052
rect 8572 5080 8584 5083
rect 9677 5083 9735 5089
rect 9677 5080 9689 5083
rect 8572 5052 9689 5080
rect 8572 5049 8584 5052
rect 8526 5043 8584 5049
rect 9677 5049 9689 5052
rect 9723 5080 9735 5083
rect 9766 5080 9772 5092
rect 9723 5052 9772 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 9766 5040 9772 5052
rect 9824 5040 9830 5092
rect 10060 5024 10088 5120
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 10704 5080 10732 5188
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 14734 5216 14740 5228
rect 13872 5188 14740 5216
rect 13872 5176 13878 5188
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 14976 5188 15393 5216
rect 14976 5176 14982 5188
rect 15381 5185 15393 5188
rect 15427 5216 15439 5219
rect 16390 5216 16396 5228
rect 15427 5188 16396 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16632 5188 16773 5216
rect 16632 5176 16638 5188
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 20162 5216 20168 5228
rect 20123 5188 20168 5216
rect 16761 5179 16819 5185
rect 20162 5176 20168 5188
rect 20220 5176 20226 5228
rect 25866 5216 25872 5228
rect 25827 5188 25872 5216
rect 25866 5176 25872 5188
rect 25924 5176 25930 5228
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5216 27859 5219
rect 27982 5216 27988 5228
rect 27847 5188 27988 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28902 5176 28908 5228
rect 28960 5216 28966 5228
rect 28997 5219 29055 5225
rect 28997 5216 29009 5219
rect 28960 5188 29009 5216
rect 28960 5176 28966 5188
rect 28997 5185 29009 5188
rect 29043 5216 29055 5219
rect 31435 5219 31493 5225
rect 31435 5216 31447 5219
rect 29043 5188 31447 5216
rect 29043 5185 29055 5188
rect 28997 5179 29055 5185
rect 31435 5185 31447 5188
rect 31481 5185 31493 5219
rect 31435 5179 31493 5185
rect 16206 5148 16212 5160
rect 16167 5120 16212 5148
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16669 5151 16727 5157
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 17126 5148 17132 5160
rect 16715 5120 17132 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 10918 5083 10976 5089
rect 10918 5080 10930 5083
rect 10704 5052 10930 5080
rect 10918 5049 10930 5052
rect 10964 5049 10976 5083
rect 13170 5080 13176 5092
rect 13131 5052 13176 5080
rect 10918 5043 10976 5049
rect 13170 5040 13176 5052
rect 13228 5040 13234 5092
rect 13265 5083 13323 5089
rect 13265 5049 13277 5083
rect 13311 5049 13323 5083
rect 14826 5080 14832 5092
rect 14787 5052 14832 5080
rect 13265 5043 13323 5049
rect 10042 5012 10048 5024
rect 3660 4984 4108 5012
rect 10003 4984 10048 5012
rect 3660 4972 3666 4984
rect 10042 4972 10048 4984
rect 10100 4972 10106 5024
rect 11517 5015 11575 5021
rect 11517 4981 11529 5015
rect 11563 5012 11575 5015
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 11563 4984 13001 5012
rect 11563 4981 11575 4984
rect 11517 4975 11575 4981
rect 12989 4981 13001 4984
rect 13035 5012 13047 5015
rect 13280 5012 13308 5043
rect 14826 5040 14832 5052
rect 14884 5040 14890 5092
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 16117 5083 16175 5089
rect 16117 5080 16129 5083
rect 15160 5052 16129 5080
rect 15160 5040 15166 5052
rect 16117 5049 16129 5052
rect 16163 5080 16175 5083
rect 16684 5080 16712 5111
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 18233 5151 18291 5157
rect 18233 5117 18245 5151
rect 18279 5148 18291 5151
rect 19705 5151 19763 5157
rect 18279 5120 19012 5148
rect 18279 5117 18291 5120
rect 18233 5111 18291 5117
rect 16163 5052 16712 5080
rect 18049 5083 18107 5089
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 18049 5049 18061 5083
rect 18095 5049 18107 5083
rect 18049 5043 18107 5049
rect 13722 5012 13728 5024
rect 13035 4984 13728 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13722 4972 13728 4984
rect 13780 4972 13786 5024
rect 15562 4972 15568 5024
rect 15620 5012 15626 5024
rect 15657 5015 15715 5021
rect 15657 5012 15669 5015
rect 15620 4984 15669 5012
rect 15620 4972 15626 4984
rect 15657 4981 15669 4984
rect 15703 4981 15715 5015
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 15657 4975 15715 4981
rect 17770 4972 17776 4984
rect 17828 5012 17834 5024
rect 18064 5012 18092 5043
rect 18984 5021 19012 5120
rect 19705 5117 19717 5151
rect 19751 5148 19763 5151
rect 19794 5148 19800 5160
rect 19751 5120 19800 5148
rect 19751 5117 19763 5120
rect 19705 5111 19763 5117
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20530 5148 20536 5160
rect 20027 5120 20536 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 19058 5040 19064 5092
rect 19116 5080 19122 5092
rect 19996 5080 20024 5111
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 21726 5148 21732 5160
rect 21687 5120 21732 5148
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 23290 5108 23296 5160
rect 23348 5148 23354 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23348 5120 23673 5148
rect 23348 5108 23354 5120
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23661 5111 23719 5117
rect 24213 5151 24271 5157
rect 24213 5117 24225 5151
rect 24259 5117 24271 5151
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 24213 5111 24271 5117
rect 19116 5052 20024 5080
rect 19116 5040 19122 5052
rect 20622 5040 20628 5092
rect 20680 5080 20686 5092
rect 21269 5083 21327 5089
rect 21269 5080 21281 5083
rect 20680 5052 21281 5080
rect 20680 5040 20686 5052
rect 21269 5049 21281 5052
rect 21315 5049 21327 5083
rect 21269 5043 21327 5049
rect 22554 5040 22560 5092
rect 22612 5080 22618 5092
rect 22925 5083 22983 5089
rect 22925 5080 22937 5083
rect 22612 5052 22937 5080
rect 22612 5040 22618 5052
rect 22925 5049 22937 5052
rect 22971 5080 22983 5083
rect 24026 5080 24032 5092
rect 22971 5052 24032 5080
rect 22971 5049 22983 5052
rect 22925 5043 22983 5049
rect 24026 5040 24032 5052
rect 24084 5080 24090 5092
rect 24228 5080 24256 5111
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 25777 5151 25835 5157
rect 25777 5117 25789 5151
rect 25823 5148 25835 5151
rect 26050 5148 26056 5160
rect 25823 5120 26056 5148
rect 25823 5117 25835 5120
rect 25777 5111 25835 5117
rect 25314 5080 25320 5092
rect 24084 5052 25320 5080
rect 24084 5040 24090 5052
rect 25314 5040 25320 5052
rect 25372 5080 25378 5092
rect 25792 5080 25820 5111
rect 26050 5108 26056 5120
rect 26108 5108 26114 5160
rect 29340 5151 29398 5157
rect 29340 5117 29352 5151
rect 29386 5148 29398 5151
rect 29730 5148 29736 5160
rect 29386 5120 29736 5148
rect 29386 5117 29398 5120
rect 29340 5111 29398 5117
rect 29730 5108 29736 5120
rect 29788 5108 29794 5160
rect 30352 5151 30410 5157
rect 30352 5117 30364 5151
rect 30398 5148 30410 5151
rect 30561 5151 30619 5157
rect 30561 5148 30573 5151
rect 30398 5120 30573 5148
rect 30398 5117 30410 5120
rect 30352 5111 30410 5117
rect 30561 5117 30573 5120
rect 30607 5117 30619 5151
rect 30561 5111 30619 5117
rect 31294 5108 31300 5160
rect 31352 5157 31358 5160
rect 31352 5151 31390 5157
rect 31378 5148 31390 5151
rect 34952 5151 35010 5157
rect 31378 5120 31800 5148
rect 31378 5117 31390 5120
rect 31352 5111 31390 5117
rect 31352 5108 31358 5111
rect 25372 5052 25820 5080
rect 27157 5083 27215 5089
rect 25372 5040 25378 5052
rect 27157 5049 27169 5083
rect 27203 5049 27215 5083
rect 27157 5043 27215 5049
rect 17828 4984 18092 5012
rect 18969 5015 19027 5021
rect 17828 4972 17834 4984
rect 18969 4981 18981 5015
rect 19015 5012 19027 5015
rect 19150 5012 19156 5024
rect 19015 4984 19156 5012
rect 19015 4981 19027 4984
rect 18969 4975 19027 4981
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 23293 5015 23351 5021
rect 23293 4981 23305 5015
rect 23339 5012 23351 5015
rect 23382 5012 23388 5024
rect 23339 4984 23388 5012
rect 23339 4981 23351 4984
rect 23293 4975 23351 4981
rect 23382 4972 23388 4984
rect 23440 4972 23446 5024
rect 23658 4972 23664 5024
rect 23716 5012 23722 5024
rect 23753 5015 23811 5021
rect 23753 5012 23765 5015
rect 23716 4984 23765 5012
rect 23716 4972 23722 4984
rect 23753 4981 23765 4984
rect 23799 4981 23811 5015
rect 27172 5012 27200 5043
rect 27246 5040 27252 5092
rect 27304 5080 27310 5092
rect 27304 5052 27349 5080
rect 27304 5040 27310 5052
rect 31772 5024 31800 5120
rect 34952 5117 34964 5151
rect 34998 5148 35010 5151
rect 34998 5120 35480 5148
rect 34998 5117 35010 5120
rect 34952 5111 35010 5117
rect 35452 5024 35480 5120
rect 28166 5012 28172 5024
rect 27172 4984 28172 5012
rect 23753 4975 23811 4981
rect 28166 4972 28172 4984
rect 28224 4972 28230 5024
rect 28534 5012 28540 5024
rect 28495 4984 28540 5012
rect 28534 4972 28540 4984
rect 28592 4972 28598 5024
rect 31754 4972 31760 5024
rect 31812 5012 31818 5024
rect 35434 5012 35440 5024
rect 31812 4984 31857 5012
rect 35395 4984 35440 5012
rect 31812 4972 31818 4984
rect 35434 4972 35440 4984
rect 35492 4972 35498 5024
rect 35986 5012 35992 5024
rect 35947 4984 35992 5012
rect 35986 4972 35992 4984
rect 36044 4972 36050 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2038 4808 2044 4820
rect 1995 4780 2044 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2038 4768 2044 4780
rect 2096 4808 2102 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 2096 4780 2237 4808
rect 2096 4768 2102 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 3789 4811 3847 4817
rect 3789 4808 3801 4811
rect 3752 4780 3801 4808
rect 3752 4768 3758 4780
rect 3789 4777 3801 4780
rect 3835 4808 3847 4811
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 3835 4780 4169 4808
rect 3835 4777 3847 4780
rect 3789 4771 3847 4777
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 6730 4768 6736 4820
rect 6788 4808 6794 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 6788 4780 7665 4808
rect 6788 4768 6794 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 10686 4808 10692 4820
rect 10647 4780 10692 4808
rect 7653 4771 7711 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12345 4811 12403 4817
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 12434 4808 12440 4820
rect 12391 4780 12440 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 13446 4808 13452 4820
rect 13407 4780 13452 4808
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14737 4811 14795 4817
rect 14737 4777 14749 4811
rect 14783 4808 14795 4811
rect 14826 4808 14832 4820
rect 14783 4780 14832 4808
rect 14783 4777 14795 4780
rect 14737 4771 14795 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 17034 4768 17040 4820
rect 17092 4808 17098 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17092 4780 17785 4808
rect 17092 4768 17098 4780
rect 17773 4777 17785 4780
rect 17819 4808 17831 4811
rect 17819 4780 18828 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 2682 4740 2688 4752
rect 2639 4712 2688 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 6362 4740 6368 4752
rect 6323 4712 6368 4740
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 8202 4700 8208 4752
rect 8260 4740 8266 4752
rect 8849 4743 8907 4749
rect 8849 4740 8861 4743
rect 8260 4712 8861 4740
rect 8260 4700 8266 4712
rect 8849 4709 8861 4712
rect 8895 4740 8907 4743
rect 9766 4740 9772 4752
rect 8895 4712 9772 4740
rect 8895 4709 8907 4712
rect 8849 4703 8907 4709
rect 9766 4700 9772 4712
rect 9824 4700 9830 4752
rect 13814 4740 13820 4752
rect 13775 4712 13820 4740
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14369 4743 14427 4749
rect 14369 4709 14381 4743
rect 14415 4740 14427 4743
rect 14918 4740 14924 4752
rect 14415 4712 14924 4740
rect 14415 4709 14427 4712
rect 14369 4703 14427 4709
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 15105 4743 15163 4749
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 16390 4740 16396 4752
rect 15151 4712 16396 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 1464 4675 1522 4681
rect 1464 4641 1476 4675
rect 1510 4672 1522 4675
rect 1670 4672 1676 4684
rect 1510 4644 1676 4672
rect 1510 4641 1522 4644
rect 1464 4635 1522 4641
rect 1670 4632 1676 4644
rect 1728 4672 1734 4684
rect 4341 4675 4399 4681
rect 1728 4644 2303 4672
rect 1728 4632 1734 4644
rect 2275 4536 2303 4644
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4522 4672 4528 4684
rect 4483 4644 4528 4672
rect 4341 4635 4399 4641
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2682 4604 2688 4616
rect 2547 4576 2688 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2958 4604 2964 4616
rect 2919 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 4356 4604 4384 4635
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 5534 4672 5540 4684
rect 5495 4644 5540 4672
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5902 4681 5908 4684
rect 5875 4675 5908 4681
rect 5684 4644 5729 4672
rect 5684 4632 5690 4644
rect 5875 4641 5887 4675
rect 5875 4635 5908 4641
rect 5902 4632 5908 4635
rect 5960 4632 5966 4684
rect 7190 4672 7196 4684
rect 7151 4644 7196 4672
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7466 4672 7472 4684
rect 7427 4644 7472 4672
rect 7466 4632 7472 4644
rect 7524 4632 7530 4684
rect 9677 4675 9735 4681
rect 9677 4641 9689 4675
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 4430 4604 4436 4616
rect 4356 4576 4436 4604
rect 4430 4564 4436 4576
rect 4488 4564 4494 4616
rect 9692 4604 9720 4635
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9916 4644 9965 4672
rect 9916 4632 9922 4644
rect 9953 4641 9965 4644
rect 9999 4672 10011 4675
rect 10962 4672 10968 4684
rect 9999 4644 10968 4672
rect 9999 4641 10011 4644
rect 9953 4635 10011 4641
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 12250 4672 12256 4684
rect 12211 4644 12256 4672
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12618 4672 12624 4684
rect 12579 4644 12624 4672
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 15286 4672 15292 4684
rect 15247 4644 15292 4672
rect 15286 4632 15292 4644
rect 15344 4632 15350 4684
rect 15488 4681 15516 4712
rect 16390 4700 16396 4712
rect 16448 4740 16454 4752
rect 16666 4740 16672 4752
rect 16448 4712 16672 4740
rect 16448 4700 16454 4712
rect 16666 4700 16672 4712
rect 16724 4700 16730 4752
rect 17494 4700 17500 4752
rect 17552 4740 17558 4752
rect 17552 4712 18276 4740
rect 17552 4700 17558 4712
rect 15473 4675 15531 4681
rect 15473 4641 15485 4675
rect 15519 4641 15531 4675
rect 15838 4672 15844 4684
rect 15799 4644 15844 4672
rect 15473 4635 15531 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 16298 4632 16304 4684
rect 16356 4672 16362 4684
rect 18248 4681 18276 4712
rect 16816 4675 16874 4681
rect 16816 4672 16828 4675
rect 16356 4644 16828 4672
rect 16356 4632 16362 4644
rect 16816 4641 16828 4644
rect 16862 4641 16874 4675
rect 18049 4675 18107 4681
rect 18049 4672 18061 4675
rect 16816 4635 16874 4641
rect 17052 4644 18061 4672
rect 10134 4604 10140 4616
rect 9692 4576 9904 4604
rect 10095 4576 10140 4604
rect 4890 4536 4896 4548
rect 2275 4508 4896 4536
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5258 4496 5264 4548
rect 5316 4536 5322 4548
rect 5721 4539 5779 4545
rect 5721 4536 5733 4539
rect 5316 4508 5733 4536
rect 5316 4496 5322 4508
rect 5721 4505 5733 4508
rect 5767 4536 5779 4539
rect 7009 4539 7067 4545
rect 7009 4536 7021 4539
rect 5767 4508 7021 4536
rect 5767 4505 5779 4508
rect 5721 4499 5779 4505
rect 7009 4505 7021 4508
rect 7055 4536 7067 4539
rect 7098 4536 7104 4548
rect 7055 4508 7104 4536
rect 7055 4505 7067 4508
rect 7009 4499 7067 4505
rect 7098 4496 7104 4508
rect 7156 4536 7162 4548
rect 7285 4539 7343 4545
rect 7285 4536 7297 4539
rect 7156 4508 7297 4536
rect 7156 4496 7162 4508
rect 7285 4505 7297 4508
rect 7331 4505 7343 4539
rect 7285 4499 7343 4505
rect 8478 4496 8484 4548
rect 8536 4536 8542 4548
rect 9769 4539 9827 4545
rect 9769 4536 9781 4539
rect 8536 4508 9781 4536
rect 8536 4496 8542 4508
rect 9769 4505 9781 4508
rect 9815 4505 9827 4539
rect 9876 4536 9904 4576
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 17052 4613 17080 4644
rect 18049 4641 18061 4644
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4641 18291 4675
rect 18233 4635 18291 4641
rect 18690 4632 18696 4684
rect 18748 4672 18754 4684
rect 18800 4681 18828 4780
rect 19242 4768 19248 4820
rect 19300 4808 19306 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 19300 4780 19349 4808
rect 19300 4768 19306 4780
rect 19337 4777 19349 4780
rect 19383 4777 19395 4811
rect 19978 4808 19984 4820
rect 19939 4780 19984 4808
rect 19337 4771 19395 4777
rect 19978 4768 19984 4780
rect 20036 4768 20042 4820
rect 20714 4808 20720 4820
rect 20675 4780 20720 4808
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 20806 4768 20812 4820
rect 20864 4808 20870 4820
rect 20901 4811 20959 4817
rect 20901 4808 20913 4811
rect 20864 4780 20913 4808
rect 20864 4768 20870 4780
rect 20901 4777 20913 4780
rect 20947 4777 20959 4811
rect 20901 4771 20959 4777
rect 23290 4768 23296 4820
rect 23348 4808 23354 4820
rect 23661 4811 23719 4817
rect 23661 4808 23673 4811
rect 23348 4780 23673 4808
rect 23348 4768 23354 4780
rect 23661 4777 23673 4780
rect 23707 4777 23719 4811
rect 23661 4771 23719 4777
rect 25130 4768 25136 4820
rect 25188 4808 25194 4820
rect 25777 4811 25835 4817
rect 25777 4808 25789 4811
rect 25188 4780 25789 4808
rect 25188 4768 25194 4780
rect 25777 4777 25789 4780
rect 25823 4777 25835 4811
rect 25777 4771 25835 4777
rect 27154 4768 27160 4820
rect 27212 4808 27218 4820
rect 27617 4811 27675 4817
rect 27617 4808 27629 4811
rect 27212 4780 27629 4808
rect 27212 4768 27218 4780
rect 27617 4777 27629 4780
rect 27663 4808 27675 4811
rect 28534 4808 28540 4820
rect 27663 4780 28540 4808
rect 27663 4777 27675 4780
rect 27617 4771 27675 4777
rect 28534 4768 28540 4780
rect 28592 4768 28598 4820
rect 29086 4768 29092 4820
rect 29144 4808 29150 4820
rect 29779 4811 29837 4817
rect 29779 4808 29791 4811
rect 29144 4780 29791 4808
rect 29144 4768 29150 4780
rect 29779 4777 29791 4780
rect 29825 4777 29837 4811
rect 29779 4771 29837 4777
rect 30193 4811 30251 4817
rect 30193 4777 30205 4811
rect 30239 4808 30251 4811
rect 30282 4808 30288 4820
rect 30239 4780 30288 4808
rect 30239 4777 30251 4780
rect 30193 4771 30251 4777
rect 18966 4740 18972 4752
rect 18927 4712 18972 4740
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 25501 4743 25559 4749
rect 25501 4709 25513 4743
rect 25547 4740 25559 4743
rect 26142 4740 26148 4752
rect 25547 4712 26148 4740
rect 25547 4709 25559 4712
rect 25501 4703 25559 4709
rect 26142 4700 26148 4712
rect 26200 4700 26206 4752
rect 28718 4700 28724 4752
rect 28776 4740 28782 4752
rect 28813 4743 28871 4749
rect 28813 4740 28825 4743
rect 28776 4712 28825 4740
rect 28776 4700 28782 4712
rect 28813 4709 28825 4712
rect 28859 4709 28871 4743
rect 30208 4740 30236 4771
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 28813 4703 28871 4709
rect 29564 4712 30236 4740
rect 18785 4675 18843 4681
rect 18785 4672 18797 4675
rect 18748 4644 18797 4672
rect 18748 4632 18754 4644
rect 18785 4641 18797 4644
rect 18831 4672 18843 4675
rect 19058 4672 19064 4684
rect 18831 4644 19064 4672
rect 18831 4641 18843 4644
rect 18785 4635 18843 4641
rect 19058 4632 19064 4644
rect 19116 4632 19122 4684
rect 19334 4632 19340 4684
rect 19392 4672 19398 4684
rect 19797 4675 19855 4681
rect 19797 4672 19809 4675
rect 19392 4644 19809 4672
rect 19392 4632 19398 4644
rect 19797 4641 19809 4644
rect 19843 4672 19855 4675
rect 20257 4675 20315 4681
rect 20257 4672 20269 4675
rect 19843 4644 20269 4672
rect 19843 4641 19855 4644
rect 19797 4635 19855 4641
rect 20257 4641 20269 4644
rect 20303 4641 20315 4675
rect 20257 4635 20315 4641
rect 22373 4675 22431 4681
rect 22373 4641 22385 4675
rect 22419 4672 22431 4675
rect 22738 4672 22744 4684
rect 22419 4644 22744 4672
rect 22419 4641 22431 4644
rect 22373 4635 22431 4641
rect 22738 4632 22744 4644
rect 22796 4632 22802 4684
rect 22922 4672 22928 4684
rect 22883 4644 22928 4672
rect 22922 4632 22928 4644
rect 22980 4632 22986 4684
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4641 25099 4675
rect 25314 4672 25320 4684
rect 25275 4644 25320 4672
rect 25041 4635 25099 4641
rect 17037 4607 17095 4613
rect 17037 4604 17049 4607
rect 16684 4576 17049 4604
rect 9950 4536 9956 4548
rect 9876 4508 9956 4536
rect 9769 4499 9827 4505
rect 1535 4471 1593 4477
rect 1535 4437 1547 4471
rect 1581 4468 1593 4471
rect 1946 4468 1952 4480
rect 1581 4440 1952 4468
rect 1581 4437 1593 4440
rect 1535 4431 1593 4437
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 8386 4468 8392 4480
rect 8347 4440 8392 4468
rect 8386 4428 8392 4440
rect 8444 4428 8450 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 9582 4468 9588 4480
rect 9539 4440 9588 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9784 4468 9812 4499
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 16684 4480 16712 4576
rect 17037 4573 17049 4576
rect 17083 4573 17095 4607
rect 17037 4567 17095 4573
rect 17126 4564 17132 4616
rect 17184 4604 17190 4616
rect 22833 4607 22891 4613
rect 22833 4604 22845 4607
rect 17184 4576 17229 4604
rect 22296 4576 22845 4604
rect 17184 4564 17190 4576
rect 22296 4480 22324 4576
rect 22833 4573 22845 4576
rect 22879 4573 22891 4607
rect 25056 4604 25084 4635
rect 25314 4632 25320 4644
rect 25372 4632 25378 4684
rect 27154 4672 27160 4684
rect 27115 4644 27160 4672
rect 27154 4632 27160 4644
rect 27212 4632 27218 4684
rect 28074 4672 28080 4684
rect 28035 4644 28080 4672
rect 28074 4632 28080 4644
rect 28132 4632 28138 4684
rect 28258 4632 28264 4684
rect 28316 4672 28322 4684
rect 28629 4675 28687 4681
rect 28629 4672 28641 4675
rect 28316 4644 28641 4672
rect 28316 4632 28322 4644
rect 28629 4641 28641 4644
rect 28675 4672 28687 4675
rect 29564 4672 29592 4712
rect 28675 4644 29592 4672
rect 29708 4675 29766 4681
rect 28675 4641 28687 4644
rect 28629 4635 28687 4641
rect 29708 4641 29720 4675
rect 29754 4672 29766 4675
rect 30190 4672 30196 4684
rect 29754 4644 30196 4672
rect 29754 4641 29766 4644
rect 29708 4635 29766 4641
rect 30190 4632 30196 4644
rect 30248 4632 30254 4684
rect 25774 4604 25780 4616
rect 25056 4576 25780 4604
rect 22833 4567 22891 4573
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 26510 4604 26516 4616
rect 26471 4576 26516 4604
rect 26510 4564 26516 4576
rect 26568 4564 26574 4616
rect 10870 4468 10876 4480
rect 9784 4440 10876 4468
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11882 4468 11888 4480
rect 11843 4440 11888 4468
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 12492 4440 13093 4468
rect 12492 4428 12498 4440
rect 13081 4437 13093 4440
rect 13127 4468 13139 4471
rect 13170 4468 13176 4480
rect 13127 4440 13176 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 16485 4471 16543 4477
rect 16485 4437 16497 4471
rect 16531 4468 16543 4471
rect 16666 4468 16672 4480
rect 16531 4440 16672 4468
rect 16531 4437 16543 4440
rect 16485 4431 16543 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 16942 4468 16948 4480
rect 16855 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4468 17006 4480
rect 18046 4468 18052 4480
rect 17000 4440 18052 4468
rect 17000 4428 17006 4440
rect 18046 4428 18052 4440
rect 18104 4428 18110 4480
rect 19705 4471 19763 4477
rect 19705 4437 19717 4471
rect 19751 4468 19763 4471
rect 19886 4468 19892 4480
rect 19751 4440 19892 4468
rect 19751 4437 19763 4440
rect 19705 4431 19763 4437
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 22278 4468 22284 4480
rect 21775 4440 22284 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 22278 4428 22284 4440
rect 22336 4428 22342 4480
rect 23198 4428 23204 4480
rect 23256 4468 23262 4480
rect 24486 4468 24492 4480
rect 23256 4440 23301 4468
rect 24447 4440 24492 4468
rect 23256 4428 23262 4440
rect 24486 4428 24492 4440
rect 24544 4428 24550 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4580 4236 4813 4264
rect 4580 4224 4586 4236
rect 4801 4233 4813 4236
rect 4847 4264 4859 4267
rect 4890 4264 4896 4276
rect 4847 4236 4896 4264
rect 4847 4233 4859 4236
rect 4801 4227 4859 4233
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5258 4264 5264 4276
rect 5219 4236 5264 4264
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 7098 4264 7104 4276
rect 7059 4236 7104 4264
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 12250 4264 12256 4276
rect 11931 4236 12256 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 13725 4267 13783 4273
rect 13725 4233 13737 4267
rect 13771 4264 13783 4267
rect 13814 4264 13820 4276
rect 13771 4236 13820 4264
rect 13771 4233 13783 4236
rect 13725 4227 13783 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 16301 4267 16359 4273
rect 16301 4264 16313 4267
rect 15396 4236 16313 4264
rect 2958 4196 2964 4208
rect 2700 4168 2964 4196
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2700 4128 2728 4168
rect 2958 4156 2964 4168
rect 3016 4156 3022 4208
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5902 4196 5908 4208
rect 5675 4168 5908 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5902 4156 5908 4168
rect 5960 4196 5966 4208
rect 7466 4196 7472 4208
rect 5960 4168 7472 4196
rect 5960 4156 5966 4168
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 2639 4100 2728 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 8220 4100 8708 4128
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3694 4060 3700 4072
rect 3655 4032 3700 4060
rect 3694 4020 3700 4032
rect 3752 4020 3758 4072
rect 3970 4060 3976 4072
rect 3931 4032 3976 4060
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 5718 4060 5724 4072
rect 5679 4032 5724 4060
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4060 6699 4063
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 6687 4032 7481 4060
rect 6687 4029 6699 4032
rect 6641 4023 6699 4029
rect 7469 4029 7481 4032
rect 7515 4060 7527 4063
rect 8110 4060 8116 4072
rect 7515 4032 8116 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 2096 3964 2141 3992
rect 2096 3952 2102 3964
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5626 3992 5632 4004
rect 5040 3964 5632 3992
rect 5040 3952 5046 3964
rect 5626 3952 5632 3964
rect 5684 3992 5690 4004
rect 6181 3995 6239 4001
rect 6181 3992 6193 3995
rect 5684 3964 6193 3992
rect 5684 3952 5690 3964
rect 6181 3961 6193 3964
rect 6227 3992 6239 3995
rect 7374 3992 7380 4004
rect 6227 3964 7380 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4430 3924 4436 3936
rect 4391 3896 4436 3924
rect 4430 3884 4436 3896
rect 4488 3884 4494 3936
rect 5902 3924 5908 3936
rect 5863 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3884 5966 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7834 3924 7840 3936
rect 7524 3896 7840 3924
rect 7524 3884 7530 3896
rect 7834 3884 7840 3896
rect 7892 3924 7898 3936
rect 8220 3933 8248 4100
rect 8386 4060 8392 4072
rect 8299 4032 8392 4060
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8478 4020 8484 4072
rect 8536 4060 8542 4072
rect 8680 4069 8708 4100
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11020 4100 11345 4128
rect 11020 4088 11026 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12161 4131 12219 4137
rect 12161 4128 12173 4131
rect 11848 4100 12173 4128
rect 11848 4088 11854 4100
rect 12161 4097 12173 4100
rect 12207 4128 12219 4131
rect 12986 4128 12992 4140
rect 12207 4100 12480 4128
rect 12947 4100 12992 4128
rect 12207 4097 12219 4100
rect 12161 4091 12219 4097
rect 8665 4063 8723 4069
rect 8536 4032 8581 4060
rect 8536 4020 8542 4032
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 8665 4023 8723 4029
rect 9769 4063 9827 4069
rect 9769 4029 9781 4063
rect 9815 4060 9827 4063
rect 9950 4060 9956 4072
rect 9815 4032 9956 4060
rect 9815 4029 9827 4032
rect 9769 4023 9827 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10134 4060 10140 4072
rect 10095 4032 10140 4060
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 10505 4063 10563 4069
rect 10505 4029 10517 4063
rect 10551 4060 10563 4063
rect 10686 4060 10692 4072
rect 10551 4032 10692 4060
rect 10551 4029 10563 4032
rect 10505 4023 10563 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 12452 4069 12480 4100
rect 12986 4088 12992 4100
rect 13044 4088 13050 4140
rect 15102 4128 15108 4140
rect 13096 4100 15108 4128
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 12710 4020 12716 4072
rect 12768 4060 12774 4072
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12768 4032 12909 4060
rect 12768 4020 12774 4032
rect 12897 4029 12909 4032
rect 12943 4060 12955 4063
rect 13096 4060 13124 4100
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 12943 4032 13124 4060
rect 14737 4063 14795 4069
rect 12943 4029 12955 4032
rect 12897 4023 12955 4029
rect 14737 4029 14749 4063
rect 14783 4060 14795 4063
rect 14918 4060 14924 4072
rect 14783 4032 14924 4060
rect 14783 4029 14795 4032
rect 14737 4023 14795 4029
rect 14918 4020 14924 4032
rect 14976 4060 14982 4072
rect 15396 4069 15424 4236
rect 16301 4233 16313 4236
rect 16347 4264 16359 4267
rect 16942 4264 16948 4276
rect 16347 4236 16948 4264
rect 16347 4233 16359 4236
rect 16301 4227 16359 4233
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 19886 4264 19892 4276
rect 18104 4236 19892 4264
rect 18104 4224 18110 4236
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 24026 4264 24032 4276
rect 23987 4236 24032 4264
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 25774 4264 25780 4276
rect 25735 4236 25780 4264
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 27154 4224 27160 4276
rect 27212 4264 27218 4276
rect 27249 4267 27307 4273
rect 27249 4264 27261 4267
rect 27212 4236 27261 4264
rect 27212 4224 27218 4236
rect 27249 4233 27261 4236
rect 27295 4233 27307 4267
rect 27249 4227 27307 4233
rect 27709 4267 27767 4273
rect 27709 4233 27721 4267
rect 27755 4264 27767 4267
rect 27985 4267 28043 4273
rect 27985 4264 27997 4267
rect 27755 4236 27997 4264
rect 27755 4233 27767 4236
rect 27709 4227 27767 4233
rect 27985 4233 27997 4236
rect 28031 4264 28043 4267
rect 28258 4264 28264 4276
rect 28031 4236 28264 4264
rect 28031 4233 28043 4236
rect 27985 4227 28043 4233
rect 28258 4224 28264 4236
rect 28316 4224 28322 4276
rect 30190 4264 30196 4276
rect 30103 4236 30196 4264
rect 30190 4224 30196 4236
rect 30248 4264 30254 4276
rect 35434 4264 35440 4276
rect 30248 4236 35440 4264
rect 30248 4224 30254 4236
rect 35434 4224 35440 4236
rect 35492 4224 35498 4276
rect 16574 4196 16580 4208
rect 15580 4168 16580 4196
rect 15580 4140 15608 4168
rect 16574 4156 16580 4168
rect 16632 4196 16638 4208
rect 16669 4199 16727 4205
rect 16669 4196 16681 4199
rect 16632 4168 16681 4196
rect 16632 4156 16638 4168
rect 16669 4165 16681 4168
rect 16715 4165 16727 4199
rect 16669 4159 16727 4165
rect 17589 4199 17647 4205
rect 17589 4165 17601 4199
rect 17635 4196 17647 4199
rect 19521 4199 19579 4205
rect 19521 4196 19533 4199
rect 17635 4168 19533 4196
rect 17635 4165 17647 4168
rect 17589 4159 17647 4165
rect 19521 4165 19533 4168
rect 19567 4196 19579 4199
rect 19751 4199 19809 4205
rect 19751 4196 19763 4199
rect 19567 4168 19763 4196
rect 19567 4165 19579 4168
rect 19521 4159 19579 4165
rect 19751 4165 19763 4168
rect 19797 4165 19809 4199
rect 25130 4196 25136 4208
rect 19751 4159 19809 4165
rect 24780 4168 25136 4196
rect 15562 4128 15568 4140
rect 15523 4100 15568 4128
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17034 4128 17040 4140
rect 16816 4100 16861 4128
rect 16995 4100 17040 4128
rect 16816 4088 16822 4100
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18138 4128 18144 4140
rect 17911 4100 18144 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 19981 4131 20039 4137
rect 19981 4128 19993 4131
rect 19076 4100 19993 4128
rect 15381 4063 15439 4069
rect 15381 4060 15393 4063
rect 14976 4032 15393 4060
rect 14976 4020 14982 4032
rect 15381 4029 15393 4032
rect 15427 4029 15439 4063
rect 16390 4060 16396 4072
rect 16351 4032 16396 4060
rect 15381 4023 15439 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 16482 4020 16488 4072
rect 16540 4069 16546 4072
rect 16540 4063 16598 4069
rect 16540 4029 16552 4063
rect 16586 4060 16598 4063
rect 17954 4060 17960 4072
rect 16586 4032 17960 4060
rect 16586 4029 16598 4032
rect 16540 4023 16598 4029
rect 16540 4020 16546 4023
rect 17954 4020 17960 4032
rect 18012 4060 18018 4072
rect 19076 4069 19104 4100
rect 19981 4097 19993 4100
rect 20027 4097 20039 4131
rect 19981 4091 20039 4097
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 18012 4032 18061 4060
rect 18012 4020 18018 4032
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18279 4063 18337 4069
rect 18279 4060 18291 4063
rect 18049 4023 18107 4029
rect 18156 4032 18291 4060
rect 8404 3992 8432 4020
rect 9030 3992 9036 4004
rect 8404 3964 9036 3992
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 16298 3952 16304 4004
rect 16356 3992 16362 4004
rect 17405 3995 17463 4001
rect 17405 3992 17417 3995
rect 16356 3964 17417 3992
rect 16356 3952 16362 3964
rect 17405 3961 17417 3964
rect 17451 3992 17463 3995
rect 17589 3995 17647 4001
rect 17589 3992 17601 3995
rect 17451 3964 17601 3992
rect 17451 3961 17463 3964
rect 17405 3955 17463 3961
rect 17589 3961 17601 3964
rect 17635 3961 17647 3995
rect 17589 3955 17647 3961
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 18156 3992 18184 4032
rect 18279 4029 18291 4032
rect 18325 4060 18337 4063
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 18325 4032 19073 4060
rect 18325 4029 18337 4032
rect 18279 4023 18337 4029
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 20088 4060 20116 4091
rect 22830 4088 22836 4140
rect 22888 4128 22894 4140
rect 23477 4131 23535 4137
rect 23477 4128 23489 4131
rect 22888 4100 23489 4128
rect 22888 4088 22894 4100
rect 23477 4097 23489 4100
rect 23523 4128 23535 4131
rect 24780 4128 24808 4168
rect 25130 4156 25136 4168
rect 25188 4156 25194 4208
rect 28166 4156 28172 4208
rect 28224 4196 28230 4208
rect 28224 4168 28948 4196
rect 28224 4156 28230 4168
rect 26145 4131 26203 4137
rect 26145 4128 26157 4131
rect 23523 4100 24808 4128
rect 25424 4100 26157 4128
rect 23523 4097 23535 4100
rect 23477 4091 23535 4097
rect 19300 4032 20116 4060
rect 19300 4020 19306 4032
rect 20898 4020 20904 4072
rect 20956 4060 20962 4072
rect 21453 4063 21511 4069
rect 21453 4060 21465 4063
rect 20956 4032 21465 4060
rect 20956 4020 20962 4032
rect 21453 4029 21465 4032
rect 21499 4060 21511 4063
rect 21634 4060 21640 4072
rect 21499 4032 21640 4060
rect 21499 4029 21511 4032
rect 21453 4023 21511 4029
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 22278 4060 22284 4072
rect 22239 4032 22284 4060
rect 22278 4020 22284 4032
rect 22336 4020 22342 4072
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22922 4060 22928 4072
rect 22511 4032 22928 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 18782 3992 18788 4004
rect 17828 3964 18184 3992
rect 18743 3964 18788 3992
rect 17828 3952 17834 3964
rect 18782 3952 18788 3964
rect 18840 3952 18846 4004
rect 19613 3995 19671 4001
rect 19613 3961 19625 3995
rect 19659 3992 19671 3995
rect 20625 3995 20683 4001
rect 20625 3992 20637 3995
rect 19659 3964 20637 3992
rect 19659 3961 19671 3964
rect 19613 3955 19671 3961
rect 20625 3961 20637 3964
rect 20671 3992 20683 3995
rect 20714 3992 20720 4004
rect 20671 3964 20720 3992
rect 20671 3961 20683 3964
rect 20625 3955 20683 3961
rect 20714 3952 20720 3964
rect 20772 3952 20778 4004
rect 22480 3992 22508 4023
rect 22922 4020 22928 4032
rect 22980 4060 22986 4072
rect 23017 4063 23075 4069
rect 23017 4060 23029 4063
rect 22980 4032 23029 4060
rect 22980 4020 22986 4032
rect 23017 4029 23029 4032
rect 23063 4029 23075 4063
rect 23017 4023 23075 4029
rect 23934 4020 23940 4072
rect 23992 4060 23998 4072
rect 24486 4060 24492 4072
rect 23992 4032 24492 4060
rect 23992 4020 23998 4032
rect 24486 4020 24492 4032
rect 24544 4020 24550 4072
rect 25424 4069 25452 4100
rect 26145 4097 26157 4100
rect 26191 4128 26203 4131
rect 26418 4128 26424 4140
rect 26191 4100 26424 4128
rect 26191 4097 26203 4100
rect 26145 4091 26203 4097
rect 26418 4088 26424 4100
rect 26476 4088 26482 4140
rect 28074 4088 28080 4140
rect 28132 4128 28138 4140
rect 28261 4131 28319 4137
rect 28261 4128 28273 4131
rect 28132 4100 28273 4128
rect 28132 4088 28138 4100
rect 28261 4097 28273 4100
rect 28307 4097 28319 4131
rect 28920 4128 28948 4168
rect 29411 4131 29469 4137
rect 29411 4128 29423 4131
rect 28920 4100 29423 4128
rect 28261 4091 28319 4097
rect 29411 4097 29423 4100
rect 29457 4097 29469 4131
rect 29411 4091 29469 4097
rect 25409 4063 25467 4069
rect 25409 4029 25421 4063
rect 25455 4029 25467 4063
rect 27798 4060 27804 4072
rect 27759 4032 27804 4060
rect 25409 4023 25467 4029
rect 27798 4020 27804 4032
rect 27856 4060 27862 4072
rect 28629 4063 28687 4069
rect 28629 4060 28641 4063
rect 27856 4032 28641 4060
rect 27856 4020 27862 4032
rect 28629 4029 28641 4032
rect 28675 4029 28687 4063
rect 28629 4023 28687 4029
rect 29324 4063 29382 4069
rect 29324 4029 29336 4063
rect 29370 4060 29382 4063
rect 29822 4060 29828 4072
rect 29370 4032 29828 4060
rect 29370 4029 29382 4032
rect 29324 4023 29382 4029
rect 29822 4020 29828 4032
rect 29880 4020 29886 4072
rect 30282 4060 30288 4072
rect 30243 4032 30288 4060
rect 30282 4020 30288 4032
rect 30340 4060 30346 4072
rect 30745 4063 30803 4069
rect 30745 4060 30757 4063
rect 30340 4032 30757 4060
rect 30340 4020 30346 4032
rect 30745 4029 30757 4032
rect 30791 4029 30803 4063
rect 30745 4023 30803 4029
rect 21100 3964 22508 3992
rect 21100 3936 21128 3964
rect 23382 3952 23388 4004
rect 23440 3992 23446 4004
rect 24397 3995 24455 4001
rect 24397 3992 24409 3995
rect 23440 3964 24409 3992
rect 23440 3952 23446 3964
rect 24397 3961 24409 3964
rect 24443 3992 24455 3995
rect 24851 3995 24909 4001
rect 24851 3992 24863 3995
rect 24443 3964 24863 3992
rect 24443 3961 24455 3964
rect 24397 3955 24455 3961
rect 24851 3961 24863 3964
rect 24897 3992 24909 3995
rect 25038 3992 25044 4004
rect 24897 3964 25044 3992
rect 24897 3961 24909 3964
rect 24851 3955 24909 3961
rect 25038 3952 25044 3964
rect 25096 3952 25102 4004
rect 26329 3995 26387 4001
rect 26329 3992 26341 3995
rect 26252 3964 26341 3992
rect 26252 3936 26280 3964
rect 26329 3961 26341 3964
rect 26375 3961 26387 3995
rect 26329 3955 26387 3961
rect 26418 3952 26424 4004
rect 26476 3992 26482 4004
rect 26970 3992 26976 4004
rect 26476 3964 26569 3992
rect 26931 3964 26976 3992
rect 26476 3952 26482 3964
rect 26970 3952 26976 3964
rect 27028 3952 27034 4004
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7892 3896 8217 3924
rect 7892 3884 7898 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 8205 3887 8263 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 10226 3924 10232 3936
rect 10187 3896 10232 3924
rect 10226 3884 10232 3896
rect 10284 3884 10290 3936
rect 10870 3884 10876 3936
rect 10928 3924 10934 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10928 3896 11069 3924
rect 10928 3884 10934 3896
rect 11057 3893 11069 3896
rect 11103 3924 11115 3927
rect 11606 3924 11612 3936
rect 11103 3896 11612 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13998 3924 14004 3936
rect 13780 3896 14004 3924
rect 13780 3884 13786 3896
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15252 3896 15853 3924
rect 15252 3884 15258 3896
rect 15841 3893 15853 3896
rect 15887 3924 15899 3927
rect 16758 3924 16764 3936
rect 15887 3896 16764 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 21082 3924 21088 3936
rect 21043 3896 21088 3924
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21634 3884 21640 3936
rect 21692 3924 21698 3936
rect 22002 3924 22008 3936
rect 21692 3896 22008 3924
rect 21692 3884 21698 3896
rect 22002 3884 22008 3896
rect 22060 3924 22066 3936
rect 22646 3924 22652 3936
rect 22060 3896 22652 3924
rect 22060 3884 22066 3896
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 22741 3927 22799 3933
rect 22741 3893 22753 3927
rect 22787 3924 22799 3927
rect 23290 3924 23296 3936
rect 22787 3896 23296 3924
rect 22787 3893 22799 3896
rect 22741 3887 22799 3893
rect 23290 3884 23296 3896
rect 23348 3884 23354 3936
rect 26234 3884 26240 3936
rect 26292 3884 26298 3936
rect 26436 3924 26464 3952
rect 27154 3924 27160 3936
rect 26436 3896 27160 3924
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 30466 3924 30472 3936
rect 30427 3896 30472 3924
rect 30466 3884 30472 3896
rect 30524 3884 30530 3936
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1762 3720 1768 3732
rect 1723 3692 1768 3720
rect 1762 3680 1768 3692
rect 1820 3680 1826 3732
rect 1946 3680 1952 3732
rect 2004 3720 2010 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2004 3692 2697 3720
rect 2004 3680 2010 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3053 3723 3111 3729
rect 3053 3720 3065 3723
rect 2832 3692 3065 3720
rect 2832 3680 2838 3692
rect 3053 3689 3065 3692
rect 3099 3689 3111 3723
rect 3053 3683 3111 3689
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3694 3720 3700 3732
rect 3559 3692 3700 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 3528 3584 3556 3683
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 4203 3723 4261 3729
rect 4203 3689 4215 3723
rect 4249 3720 4261 3723
rect 5350 3720 5356 3732
rect 4249 3692 5356 3720
rect 4249 3689 4261 3692
rect 4203 3683 4261 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6546 3720 6552 3732
rect 6507 3692 6552 3720
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 8110 3680 8116 3732
rect 8168 3720 8174 3732
rect 8478 3720 8484 3732
rect 8168 3692 8484 3720
rect 8168 3680 8174 3692
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 9214 3720 9220 3732
rect 9175 3692 9220 3720
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9674 3680 9680 3732
rect 9732 3720 9738 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9732 3692 9781 3720
rect 9732 3680 9738 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10192 3692 10701 3720
rect 10192 3680 10198 3692
rect 10689 3689 10701 3692
rect 10735 3720 10747 3723
rect 12618 3720 12624 3732
rect 10735 3692 12624 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 12618 3680 12624 3692
rect 12676 3720 12682 3732
rect 12897 3723 12955 3729
rect 12897 3720 12909 3723
rect 12676 3692 12909 3720
rect 12676 3680 12682 3692
rect 12897 3689 12909 3692
rect 12943 3689 12955 3723
rect 12897 3683 12955 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15838 3720 15844 3732
rect 15344 3692 15844 3720
rect 15344 3680 15350 3692
rect 15838 3680 15844 3692
rect 15896 3680 15902 3732
rect 16482 3720 16488 3732
rect 16443 3692 16488 3720
rect 16482 3680 16488 3692
rect 16540 3720 16546 3732
rect 17037 3723 17095 3729
rect 17037 3720 17049 3723
rect 16540 3692 17049 3720
rect 16540 3680 16546 3692
rect 17037 3689 17049 3692
rect 17083 3689 17095 3723
rect 17586 3720 17592 3732
rect 17547 3692 17592 3720
rect 17037 3683 17095 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17862 3720 17868 3732
rect 17788 3692 17868 3720
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 5215 3655 5273 3661
rect 5215 3652 5227 3655
rect 4396 3624 5227 3652
rect 4396 3612 4402 3624
rect 5215 3621 5227 3624
rect 5261 3621 5273 3655
rect 5215 3615 5273 3621
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 7285 3655 7343 3661
rect 7285 3652 7297 3655
rect 7248 3624 7297 3652
rect 7248 3612 7254 3624
rect 7285 3621 7297 3624
rect 7331 3652 7343 3655
rect 8386 3652 8392 3664
rect 7331 3624 8392 3652
rect 7331 3621 7343 3624
rect 7285 3615 7343 3621
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 9950 3612 9956 3664
rect 10008 3652 10014 3664
rect 12250 3652 12256 3664
rect 10008 3624 11652 3652
rect 12211 3624 12256 3652
rect 10008 3612 10014 3624
rect 4154 3593 4160 3596
rect 2271 3556 3556 3584
rect 4132 3587 4160 3593
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 4132 3553 4144 3587
rect 4132 3547 4160 3553
rect 4154 3544 4160 3547
rect 4212 3544 4218 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 5112 3587 5170 3593
rect 5112 3584 5124 3587
rect 4856 3556 5124 3584
rect 4856 3544 4862 3556
rect 5112 3553 5124 3556
rect 5158 3553 5170 3587
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 5112 3547 5170 3553
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 7374 3584 7380 3596
rect 7335 3556 7380 3584
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3584 7711 3587
rect 7834 3584 7840 3596
rect 7699 3556 7840 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7668 3516 7696 3547
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 10318 3593 10324 3596
rect 10275 3587 10324 3593
rect 10275 3553 10287 3587
rect 10321 3553 10324 3587
rect 10275 3547 10324 3553
rect 10318 3544 10324 3547
rect 10376 3584 10382 3596
rect 11624 3593 11652 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 14826 3652 14832 3664
rect 14016 3624 14832 3652
rect 11609 3587 11667 3593
rect 10376 3556 11560 3584
rect 10376 3544 10382 3556
rect 7156 3488 7696 3516
rect 8113 3519 8171 3525
rect 7156 3476 7162 3488
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 8202 3516 8208 3528
rect 8159 3488 8208 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 11532 3516 11560 3556
rect 11609 3553 11621 3587
rect 11655 3584 11667 3587
rect 11790 3584 11796 3596
rect 11655 3556 11796 3584
rect 11655 3553 11667 3556
rect 11609 3547 11667 3553
rect 11790 3544 11796 3556
rect 11848 3544 11854 3596
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 12710 3584 12716 3596
rect 12667 3556 12716 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 12636 3516 12664 3547
rect 12710 3544 12716 3556
rect 12768 3544 12774 3596
rect 14016 3593 14044 3624
rect 14826 3612 14832 3624
rect 14884 3652 14890 3664
rect 17788 3661 17816 3692
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18417 3723 18475 3729
rect 18417 3689 18429 3723
rect 18463 3720 18475 3723
rect 18874 3720 18880 3732
rect 18463 3692 18880 3720
rect 18463 3689 18475 3692
rect 18417 3683 18475 3689
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 20993 3723 21051 3729
rect 20993 3720 21005 3723
rect 20864 3692 21005 3720
rect 20864 3680 20870 3692
rect 20993 3689 21005 3692
rect 21039 3689 21051 3723
rect 23934 3720 23940 3732
rect 23895 3692 23940 3720
rect 20993 3683 21051 3689
rect 15565 3655 15623 3661
rect 15565 3652 15577 3655
rect 14884 3624 15577 3652
rect 14884 3612 14890 3624
rect 15565 3621 15577 3624
rect 15611 3652 15623 3655
rect 17773 3655 17831 3661
rect 17773 3652 17785 3655
rect 15611 3624 17785 3652
rect 15611 3621 15623 3624
rect 15565 3615 15623 3621
rect 17773 3621 17785 3624
rect 17819 3621 17831 3655
rect 19886 3652 19892 3664
rect 19847 3624 19892 3652
rect 17773 3615 17831 3621
rect 19886 3612 19892 3624
rect 19944 3612 19950 3664
rect 21008 3652 21036 3683
rect 23934 3680 23940 3692
rect 23992 3680 23998 3732
rect 28629 3723 28687 3729
rect 28629 3689 28641 3723
rect 28675 3720 28687 3723
rect 29086 3720 29092 3732
rect 28675 3692 29092 3720
rect 28675 3689 28687 3692
rect 28629 3683 28687 3689
rect 29086 3680 29092 3692
rect 29144 3720 29150 3732
rect 29144 3692 29684 3720
rect 29144 3680 29150 3692
rect 24213 3655 24271 3661
rect 24213 3652 24225 3655
rect 21008 3624 24225 3652
rect 24213 3621 24225 3624
rect 24259 3621 24271 3655
rect 24213 3615 24271 3621
rect 25038 3612 25044 3664
rect 25096 3652 25102 3664
rect 28071 3655 28129 3661
rect 28071 3652 28083 3655
rect 25096 3624 28083 3652
rect 25096 3612 25102 3624
rect 28071 3621 28083 3624
rect 28117 3652 28129 3655
rect 28350 3652 28356 3664
rect 28117 3624 28356 3652
rect 28117 3621 28129 3624
rect 28071 3615 28129 3621
rect 28350 3612 28356 3624
rect 28408 3612 28414 3664
rect 29656 3661 29684 3692
rect 29641 3655 29699 3661
rect 29641 3621 29653 3655
rect 29687 3621 29699 3655
rect 29641 3615 29699 3621
rect 13909 3587 13967 3593
rect 13909 3553 13921 3587
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14001 3587 14059 3593
rect 14001 3553 14013 3587
rect 14047 3553 14059 3587
rect 14366 3584 14372 3596
rect 14327 3556 14372 3584
rect 14001 3547 14059 3553
rect 11532 3488 12664 3516
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13924 3516 13952 3547
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 16298 3584 16304 3596
rect 16259 3556 16304 3584
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 17954 3593 17960 3596
rect 17920 3587 17960 3593
rect 17920 3553 17932 3587
rect 18012 3584 18018 3596
rect 18506 3584 18512 3596
rect 18012 3556 18512 3584
rect 17920 3547 17960 3553
rect 17954 3544 17960 3547
rect 18012 3544 18018 3556
rect 18506 3544 18512 3556
rect 18564 3584 18570 3596
rect 18785 3587 18843 3593
rect 18785 3584 18797 3587
rect 18564 3556 18797 3584
rect 18564 3544 18570 3556
rect 18785 3553 18797 3556
rect 18831 3553 18843 3587
rect 19334 3584 19340 3596
rect 19295 3556 19340 3584
rect 18785 3547 18843 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 19518 3584 19524 3596
rect 19479 3556 19524 3584
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 20898 3584 20904 3596
rect 20859 3556 20904 3584
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 21361 3587 21419 3593
rect 21361 3553 21373 3587
rect 21407 3553 21419 3587
rect 21361 3547 21419 3553
rect 21729 3587 21787 3593
rect 21729 3553 21741 3587
rect 21775 3584 21787 3587
rect 21818 3584 21824 3596
rect 21775 3556 21824 3584
rect 21775 3553 21787 3556
rect 21729 3547 21787 3553
rect 14642 3516 14648 3528
rect 13228 3488 14648 3516
rect 13228 3476 13234 3488
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17828 3488 18153 3516
rect 17828 3476 17834 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18141 3479 18199 3485
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21376 3516 21404 3547
rect 21818 3544 21824 3556
rect 21876 3544 21882 3596
rect 22741 3587 22799 3593
rect 22741 3553 22753 3587
rect 22787 3584 22799 3587
rect 22830 3584 22836 3596
rect 22787 3556 22836 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 23106 3544 23112 3596
rect 23164 3584 23170 3596
rect 23661 3587 23719 3593
rect 23661 3584 23673 3587
rect 23164 3556 23673 3584
rect 23164 3544 23170 3556
rect 23661 3553 23673 3556
rect 23707 3553 23719 3587
rect 23842 3584 23848 3596
rect 23803 3556 23848 3584
rect 23661 3547 23719 3553
rect 23842 3544 23848 3556
rect 23900 3544 23906 3596
rect 24854 3584 24860 3596
rect 24815 3556 24860 3584
rect 24854 3544 24860 3556
rect 24912 3544 24918 3596
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 26548 3587 26606 3593
rect 26548 3584 26560 3587
rect 26476 3556 26560 3584
rect 26476 3544 26482 3556
rect 26548 3553 26560 3556
rect 26594 3553 26606 3587
rect 26548 3547 26606 3553
rect 22278 3516 22284 3528
rect 20772 3488 22284 3516
rect 20772 3476 20778 3488
rect 22278 3476 22284 3488
rect 22336 3476 22342 3528
rect 27709 3519 27767 3525
rect 27709 3485 27721 3519
rect 27755 3516 27767 3519
rect 27982 3516 27988 3528
rect 27755 3488 27988 3516
rect 27755 3485 27767 3488
rect 27709 3479 27767 3485
rect 27982 3476 27988 3488
rect 28040 3476 28046 3528
rect 29546 3516 29552 3528
rect 29507 3488 29552 3516
rect 29546 3476 29552 3488
rect 29604 3476 29610 3528
rect 7469 3451 7527 3457
rect 7469 3417 7481 3451
rect 7515 3417 7527 3451
rect 7469 3411 7527 3417
rect 7484 3380 7512 3411
rect 16574 3408 16580 3460
rect 16632 3448 16638 3460
rect 17954 3448 17960 3460
rect 16632 3420 17960 3448
rect 16632 3408 16638 3420
rect 17954 3408 17960 3420
rect 18012 3448 18018 3460
rect 18049 3451 18107 3457
rect 18049 3448 18061 3451
rect 18012 3420 18061 3448
rect 18012 3408 18018 3420
rect 18049 3417 18061 3420
rect 18095 3417 18107 3451
rect 18049 3411 18107 3417
rect 8110 3380 8116 3392
rect 7484 3352 8116 3380
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 14921 3383 14979 3389
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15194 3380 15200 3392
rect 14967 3352 15200 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15194 3340 15200 3352
rect 15252 3340 15258 3392
rect 18064 3380 18092 3411
rect 18322 3408 18328 3460
rect 18380 3448 18386 3460
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 18380 3420 20177 3448
rect 18380 3408 18386 3420
rect 20165 3417 20177 3420
rect 20211 3417 20223 3451
rect 20165 3411 20223 3417
rect 22296 3389 22324 3476
rect 30098 3448 30104 3460
rect 30059 3420 30104 3448
rect 30098 3408 30104 3420
rect 30156 3408 30162 3460
rect 19153 3383 19211 3389
rect 19153 3380 19165 3383
rect 18064 3352 19165 3380
rect 19153 3349 19165 3352
rect 19199 3349 19211 3383
rect 19153 3343 19211 3349
rect 22281 3383 22339 3389
rect 22281 3349 22293 3383
rect 22327 3380 22339 3383
rect 22462 3380 22468 3392
rect 22327 3352 22468 3380
rect 22327 3349 22339 3352
rect 22281 3343 22339 3349
rect 22462 3340 22468 3352
rect 22520 3340 22526 3392
rect 24578 3380 24584 3392
rect 24539 3352 24584 3380
rect 24578 3340 24584 3352
rect 24636 3340 24642 3392
rect 25222 3380 25228 3392
rect 25183 3352 25228 3380
rect 25222 3340 25228 3352
rect 25280 3340 25286 3392
rect 26234 3380 26240 3392
rect 26195 3352 26240 3380
rect 26234 3340 26240 3352
rect 26292 3340 26298 3392
rect 26326 3340 26332 3392
rect 26384 3380 26390 3392
rect 26651 3383 26709 3389
rect 26651 3380 26663 3383
rect 26384 3352 26663 3380
rect 26384 3340 26390 3352
rect 26651 3349 26663 3352
rect 26697 3380 26709 3383
rect 26973 3383 27031 3389
rect 26973 3380 26985 3383
rect 26697 3352 26985 3380
rect 26697 3349 26709 3352
rect 26651 3343 26709 3349
rect 26973 3349 26985 3352
rect 27019 3349 27031 3383
rect 26973 3343 27031 3349
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3835 3179 3893 3185
rect 3835 3176 3847 3179
rect 3292 3148 3847 3176
rect 3292 3136 3298 3148
rect 3835 3145 3847 3148
rect 3881 3145 3893 3179
rect 4154 3176 4160 3188
rect 4115 3148 4160 3176
rect 3835 3139 3893 3145
rect 4154 3136 4160 3148
rect 4212 3136 4218 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 4856 3148 5089 3176
rect 4856 3136 4862 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6362 3176 6368 3188
rect 5675 3148 6368 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 8110 3176 8116 3188
rect 7760 3148 8116 3176
rect 3421 3111 3479 3117
rect 3421 3077 3433 3111
rect 3467 3108 3479 3111
rect 3694 3108 3700 3120
rect 3467 3080 3700 3108
rect 3467 3077 3479 3080
rect 3421 3071 3479 3077
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 5905 3111 5963 3117
rect 5905 3077 5917 3111
rect 5951 3108 5963 3111
rect 5994 3108 6000 3120
rect 5951 3080 6000 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 6270 3108 6276 3120
rect 6231 3080 6276 3108
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 7760 3117 7788 3148
rect 8110 3136 8116 3148
rect 8168 3136 8174 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 9858 3176 9864 3188
rect 8803 3148 9864 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 6641 3111 6699 3117
rect 6641 3077 6653 3111
rect 6687 3108 6699 3111
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 6687 3080 7757 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 7745 3071 7803 3077
rect 2590 3040 2596 3052
rect 2551 3012 2596 3040
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 3936 3012 4537 3040
rect 3936 3000 3942 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2972 1823 2975
rect 1946 2972 1952 2984
rect 1811 2944 1952 2972
rect 1811 2941 1823 2944
rect 1765 2935 1823 2941
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 2501 2975 2559 2981
rect 2501 2972 2513 2975
rect 2188 2944 2513 2972
rect 2188 2932 2194 2944
rect 2501 2941 2513 2944
rect 2547 2972 2559 2975
rect 2958 2972 2964 2984
rect 2547 2944 2964 2972
rect 2547 2941 2559 2944
rect 2501 2935 2559 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3764 2975 3822 2981
rect 3764 2941 3776 2975
rect 3810 2972 3822 2975
rect 3896 2972 3924 3000
rect 3810 2944 3924 2972
rect 5721 2975 5779 2981
rect 3810 2941 3822 2944
rect 3764 2935 3822 2941
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6288 2972 6316 3068
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 6972 3012 8125 3040
rect 6972 3000 6978 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 7374 2972 7380 2984
rect 5767 2944 6316 2972
rect 7335 2944 7380 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2941 7711 2975
rect 7653 2935 7711 2941
rect 7668 2904 7696 2935
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7892 2944 7941 2972
rect 7892 2932 7898 2944
rect 7929 2941 7941 2944
rect 7975 2972 7987 2975
rect 8772 2972 8800 3139
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10318 3176 10324 3188
rect 10091 3148 10324 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 11471 3179 11529 3185
rect 11471 3145 11483 3179
rect 11517 3176 11529 3179
rect 12342 3176 12348 3188
rect 11517 3148 12348 3176
rect 11517 3145 11529 3148
rect 11471 3139 11529 3145
rect 12342 3136 12348 3148
rect 12400 3136 12406 3188
rect 13170 3176 13176 3188
rect 13131 3148 13176 3176
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 13403 3179 13461 3185
rect 13403 3145 13415 3179
rect 13449 3176 13461 3179
rect 13998 3176 14004 3188
rect 13449 3148 14004 3176
rect 13449 3145 13461 3148
rect 13403 3139 13461 3145
rect 13998 3136 14004 3148
rect 14056 3136 14062 3188
rect 14918 3136 14924 3188
rect 14976 3176 14982 3188
rect 15105 3179 15163 3185
rect 15105 3176 15117 3179
rect 14976 3148 15117 3176
rect 14976 3136 14982 3148
rect 15105 3145 15117 3148
rect 15151 3145 15163 3179
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15105 3139 15163 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17770 3176 17776 3188
rect 16816 3148 17776 3176
rect 16816 3136 16822 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18506 3176 18512 3188
rect 18467 3148 18512 3176
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 20257 3179 20315 3185
rect 20257 3176 20269 3179
rect 19392 3148 20269 3176
rect 19392 3136 19398 3148
rect 20257 3145 20269 3148
rect 20303 3145 20315 3179
rect 20257 3139 20315 3145
rect 21726 3136 21732 3188
rect 21784 3176 21790 3188
rect 22094 3176 22100 3188
rect 21784 3148 22100 3176
rect 21784 3136 21790 3148
rect 22094 3136 22100 3148
rect 22152 3136 22158 3188
rect 23106 3176 23112 3188
rect 23067 3148 23112 3176
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 23201 3179 23259 3185
rect 23201 3145 23213 3179
rect 23247 3176 23259 3179
rect 23474 3176 23480 3188
rect 23247 3148 23480 3176
rect 23247 3145 23259 3148
rect 23201 3139 23259 3145
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 26418 3136 26424 3188
rect 26476 3176 26482 3188
rect 27246 3176 27252 3188
rect 26476 3148 27252 3176
rect 26476 3136 26482 3148
rect 27246 3136 27252 3148
rect 27304 3136 27310 3188
rect 27709 3179 27767 3185
rect 27709 3145 27721 3179
rect 27755 3176 27767 3179
rect 27982 3176 27988 3188
rect 27755 3148 27988 3176
rect 27755 3145 27767 3148
rect 27709 3139 27767 3145
rect 27982 3136 27988 3148
rect 28040 3136 28046 3188
rect 29546 3136 29552 3188
rect 29604 3176 29610 3188
rect 30745 3179 30803 3185
rect 30745 3176 30757 3179
rect 29604 3148 30757 3176
rect 29604 3136 29610 3148
rect 30745 3145 30757 3148
rect 30791 3145 30803 3179
rect 30745 3139 30803 3145
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 9732 3080 10609 3108
rect 9732 3068 9738 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 11790 3108 11796 3120
rect 11751 3080 11796 3108
rect 10597 3071 10655 3077
rect 11790 3068 11796 3080
rect 11848 3108 11854 3120
rect 11974 3108 11980 3120
rect 11848 3080 11980 3108
rect 11848 3068 11854 3080
rect 11974 3068 11980 3080
rect 12032 3068 12038 3120
rect 12158 3108 12164 3120
rect 12119 3080 12164 3108
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 13817 3111 13875 3117
rect 13817 3077 13829 3111
rect 13863 3108 13875 3111
rect 14366 3108 14372 3120
rect 13863 3080 14372 3108
rect 13863 3077 13875 3080
rect 13817 3071 13875 3077
rect 14366 3068 14372 3080
rect 14424 3068 14430 3120
rect 16485 3111 16543 3117
rect 16485 3077 16497 3111
rect 16531 3108 16543 3111
rect 16574 3108 16580 3120
rect 16531 3080 16580 3108
rect 16531 3077 16543 3080
rect 16485 3071 16543 3077
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 22462 3108 22468 3120
rect 22375 3080 22468 3108
rect 22462 3068 22468 3080
rect 22520 3108 22526 3120
rect 23842 3108 23848 3120
rect 22520 3080 23848 3108
rect 22520 3068 22526 3080
rect 23842 3068 23848 3080
rect 23900 3068 23906 3120
rect 29472 3080 30972 3108
rect 9125 3043 9183 3049
rect 9125 3009 9137 3043
rect 9171 3040 9183 3043
rect 9766 3040 9772 3052
rect 9171 3012 9628 3040
rect 9727 3012 9772 3040
rect 9171 3009 9183 3012
rect 9125 3003 9183 3009
rect 9600 2984 9628 3012
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 9214 2972 9220 2984
rect 7975 2944 8800 2972
rect 9175 2944 9220 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9677 2975 9735 2981
rect 9677 2972 9689 2975
rect 9640 2944 9689 2972
rect 9640 2932 9646 2944
rect 9677 2941 9689 2944
rect 9723 2972 9735 2975
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9723 2944 10057 2972
rect 9723 2941 9735 2944
rect 9677 2935 9735 2941
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 11400 2975 11458 2981
rect 11400 2941 11412 2975
rect 11446 2972 11458 2975
rect 12176 2972 12204 3068
rect 29472 3052 29500 3080
rect 14182 3040 14188 3052
rect 14143 3012 14188 3040
rect 14182 3000 14188 3012
rect 14240 3000 14246 3052
rect 15194 3040 15200 3052
rect 15155 3012 15200 3040
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 17862 3040 17868 3052
rect 17543 3012 17868 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 19337 3043 19395 3049
rect 19337 3009 19349 3043
rect 19383 3040 19395 3043
rect 22695 3043 22753 3049
rect 22695 3040 22707 3043
rect 19383 3012 22707 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 22695 3009 22707 3012
rect 22741 3040 22753 3043
rect 25593 3043 25651 3049
rect 25593 3040 25605 3043
rect 22741 3012 25605 3040
rect 22741 3009 22753 3012
rect 22695 3003 22753 3009
rect 25593 3009 25605 3012
rect 25639 3009 25651 3043
rect 26326 3040 26332 3052
rect 26287 3012 26332 3040
rect 25593 3003 25651 3009
rect 26326 3000 26332 3012
rect 26384 3000 26390 3052
rect 26970 3040 26976 3052
rect 26931 3012 26976 3040
rect 26970 3000 26976 3012
rect 27028 3000 27034 3052
rect 29454 3040 29460 3052
rect 29367 3012 29460 3040
rect 29454 3000 29460 3012
rect 29512 3000 29518 3052
rect 30098 3040 30104 3052
rect 30059 3012 30104 3040
rect 30098 3000 30104 3012
rect 30156 3000 30162 3052
rect 30944 3049 30972 3080
rect 30929 3043 30987 3049
rect 30929 3009 30941 3043
rect 30975 3009 30987 3043
rect 30929 3003 30987 3009
rect 11446 2944 12204 2972
rect 13332 2975 13390 2981
rect 11446 2941 11458 2944
rect 11400 2935 11458 2941
rect 13332 2941 13344 2975
rect 13378 2972 13390 2975
rect 14200 2972 14228 3000
rect 15010 2981 15016 2984
rect 13378 2944 14228 2972
rect 14737 2975 14795 2981
rect 13378 2941 13390 2944
rect 13332 2935 13390 2941
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 14976 2975 15016 2981
rect 14976 2972 14988 2975
rect 14783 2944 14988 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 14976 2941 14988 2944
rect 15068 2972 15074 2984
rect 16025 2975 16083 2981
rect 16025 2972 16037 2975
rect 15068 2944 16037 2972
rect 14976 2935 15016 2941
rect 15010 2932 15016 2935
rect 15068 2932 15074 2944
rect 16025 2941 16037 2944
rect 16071 2972 16083 2975
rect 16298 2972 16304 2984
rect 16071 2944 16304 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 16298 2932 16304 2944
rect 16356 2972 16362 2984
rect 16393 2975 16451 2981
rect 16393 2972 16405 2975
rect 16356 2944 16405 2972
rect 16356 2932 16362 2944
rect 16393 2941 16405 2944
rect 16439 2941 16451 2975
rect 16666 2972 16672 2984
rect 16627 2944 16672 2972
rect 16393 2935 16451 2941
rect 16666 2932 16672 2944
rect 16724 2932 16730 2984
rect 17129 2975 17187 2981
rect 17129 2941 17141 2975
rect 17175 2972 17187 2975
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17175 2944 18061 2972
rect 17175 2941 17187 2944
rect 17129 2935 17187 2941
rect 18049 2941 18061 2944
rect 18095 2972 18107 2975
rect 18322 2972 18328 2984
rect 18095 2944 18328 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20254 2972 20260 2984
rect 20027 2944 20260 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20254 2932 20260 2944
rect 20312 2932 20318 2984
rect 20806 2972 20812 2984
rect 20767 2944 20812 2972
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 21726 2972 21732 2984
rect 21008 2944 21732 2972
rect 8386 2904 8392 2916
rect 7668 2876 8392 2904
rect 8386 2864 8392 2876
rect 8444 2864 8450 2916
rect 14826 2904 14832 2916
rect 14787 2876 14832 2904
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 19429 2907 19487 2913
rect 19429 2873 19441 2907
rect 19475 2904 19487 2907
rect 21008 2904 21036 2944
rect 21726 2932 21732 2944
rect 21784 2932 21790 2984
rect 22002 2972 22008 2984
rect 21963 2944 22008 2972
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 22554 2972 22560 2984
rect 22518 2944 22560 2972
rect 22554 2932 22560 2944
rect 22612 2981 22618 2984
rect 22612 2975 22666 2981
rect 22612 2941 22620 2975
rect 22654 2972 22666 2975
rect 23201 2975 23259 2981
rect 23201 2972 23213 2975
rect 22654 2944 23213 2972
rect 22654 2941 22666 2944
rect 22612 2935 22666 2941
rect 23201 2941 23213 2944
rect 23247 2941 23259 2975
rect 23201 2935 23259 2941
rect 22612 2932 22618 2935
rect 23290 2932 23296 2984
rect 23348 2972 23354 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23348 2944 23673 2972
rect 23348 2932 23354 2944
rect 23661 2941 23673 2944
rect 23707 2972 23719 2975
rect 24578 2972 24584 2984
rect 23707 2944 24584 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24578 2932 24584 2944
rect 24636 2932 24642 2984
rect 27062 2932 27068 2984
rect 27120 2972 27126 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27120 2944 27813 2972
rect 27120 2932 27126 2944
rect 27801 2941 27813 2944
rect 27847 2972 27859 2975
rect 28629 2975 28687 2981
rect 28629 2972 28641 2975
rect 27847 2944 28641 2972
rect 27847 2941 27859 2944
rect 27801 2935 27859 2941
rect 28629 2941 28641 2944
rect 28675 2941 28687 2975
rect 28629 2935 28687 2941
rect 19475 2876 21036 2904
rect 19475 2873 19487 2876
rect 19429 2867 19487 2873
rect 21082 2864 21088 2916
rect 21140 2913 21146 2916
rect 21140 2907 21188 2913
rect 21140 2873 21142 2907
rect 21176 2873 21188 2907
rect 21818 2904 21824 2916
rect 21140 2867 21188 2873
rect 21259 2876 21824 2904
rect 21140 2864 21146 2867
rect 7098 2836 7104 2848
rect 7059 2808 7104 2836
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 18233 2839 18291 2845
rect 18233 2805 18245 2839
rect 18279 2836 18291 2839
rect 18414 2836 18420 2848
rect 18279 2808 18420 2836
rect 18279 2805 18291 2808
rect 18233 2799 18291 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 19150 2836 19156 2848
rect 19111 2808 19156 2836
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 20990 2836 20996 2848
rect 20763 2808 20996 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 20990 2796 20996 2808
rect 21048 2836 21054 2848
rect 21259 2836 21287 2876
rect 21818 2864 21824 2876
rect 21876 2904 21882 2916
rect 23106 2904 23112 2916
rect 21876 2876 23112 2904
rect 21876 2864 21882 2876
rect 23106 2864 23112 2876
rect 23164 2864 23170 2916
rect 23750 2864 23756 2916
rect 23808 2904 23814 2916
rect 24023 2907 24081 2913
rect 24023 2904 24035 2907
rect 23808 2876 24035 2904
rect 23808 2864 23814 2876
rect 24023 2873 24035 2876
rect 24069 2904 24081 2907
rect 25038 2904 25044 2916
rect 24069 2876 25044 2904
rect 24069 2873 24081 2876
rect 24023 2867 24081 2873
rect 25038 2864 25044 2876
rect 25096 2864 25102 2916
rect 26145 2907 26203 2913
rect 26145 2873 26157 2907
rect 26191 2904 26203 2907
rect 26421 2907 26479 2913
rect 26421 2904 26433 2907
rect 26191 2876 26433 2904
rect 26191 2873 26203 2876
rect 26145 2867 26203 2873
rect 26421 2873 26433 2876
rect 26467 2904 26479 2907
rect 26510 2904 26516 2916
rect 26467 2876 26516 2904
rect 26467 2873 26479 2876
rect 26421 2867 26479 2873
rect 26510 2864 26516 2876
rect 26568 2864 26574 2916
rect 27614 2864 27620 2916
rect 27672 2864 27678 2916
rect 29089 2907 29147 2913
rect 29089 2873 29101 2907
rect 29135 2904 29147 2907
rect 29546 2904 29552 2916
rect 29135 2876 29552 2904
rect 29135 2873 29147 2876
rect 29089 2867 29147 2873
rect 29546 2864 29552 2876
rect 29604 2864 29610 2916
rect 21048 2808 21287 2836
rect 21048 2796 21054 2808
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24581 2839 24639 2845
rect 24581 2836 24593 2839
rect 23532 2808 24593 2836
rect 23532 2796 23538 2808
rect 24581 2805 24593 2808
rect 24627 2836 24639 2839
rect 24854 2836 24860 2848
rect 24627 2808 24860 2836
rect 24627 2805 24639 2808
rect 24581 2799 24639 2805
rect 24854 2796 24860 2808
rect 24912 2836 24918 2848
rect 25225 2839 25283 2845
rect 25225 2836 25237 2839
rect 24912 2808 25237 2836
rect 24912 2796 24918 2808
rect 25225 2805 25237 2808
rect 25271 2805 25283 2839
rect 27632 2836 27660 2864
rect 27985 2839 28043 2845
rect 27985 2836 27997 2839
rect 27632 2808 27997 2836
rect 25225 2799 25283 2805
rect 27985 2805 27997 2808
rect 28031 2805 28043 2839
rect 28350 2836 28356 2848
rect 28311 2808 28356 2836
rect 27985 2799 28043 2805
rect 28350 2796 28356 2808
rect 28408 2796 28414 2848
rect 29822 2796 29828 2848
rect 29880 2836 29886 2848
rect 30377 2839 30435 2845
rect 30377 2836 30389 2839
rect 29880 2808 30389 2836
rect 29880 2796 29886 2808
rect 30377 2805 30389 2808
rect 30423 2805 30435 2839
rect 30377 2799 30435 2805
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2363 2635 2421 2641
rect 2363 2601 2375 2635
rect 2409 2632 2421 2635
rect 2682 2632 2688 2644
rect 2409 2604 2688 2632
rect 2409 2601 2421 2604
rect 2363 2595 2421 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 8110 2632 8116 2644
rect 8071 2604 8116 2632
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8444 2604 8493 2632
rect 8444 2592 8450 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8846 2632 8852 2644
rect 8807 2604 8852 2632
rect 8481 2595 8539 2601
rect 8846 2592 8852 2604
rect 8904 2592 8910 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 11655 2635 11713 2641
rect 11655 2601 11667 2635
rect 11701 2632 11713 2635
rect 11882 2632 11888 2644
rect 11701 2604 11888 2632
rect 11701 2601 11713 2604
rect 11655 2595 11713 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 12943 2635 13001 2641
rect 12943 2601 12955 2635
rect 12989 2632 13001 2635
rect 13630 2632 13636 2644
rect 12989 2604 13636 2632
rect 12989 2601 13001 2604
rect 12943 2595 13001 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14918 2632 14924 2644
rect 14879 2604 14924 2632
rect 14918 2592 14924 2604
rect 14976 2592 14982 2644
rect 16298 2592 16304 2644
rect 16356 2632 16362 2644
rect 16577 2635 16635 2641
rect 16577 2632 16589 2635
rect 16356 2604 16589 2632
rect 16356 2592 16362 2604
rect 16577 2601 16589 2604
rect 16623 2601 16635 2635
rect 16577 2595 16635 2601
rect 16758 2592 16764 2644
rect 16816 2632 16822 2644
rect 17313 2635 17371 2641
rect 17313 2632 17325 2635
rect 16816 2604 17325 2632
rect 16816 2592 16822 2604
rect 17313 2601 17325 2604
rect 17359 2601 17371 2635
rect 17954 2632 17960 2644
rect 17915 2604 17960 2632
rect 17313 2595 17371 2601
rect 17954 2592 17960 2604
rect 18012 2592 18018 2644
rect 18690 2632 18696 2644
rect 18651 2604 18696 2632
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 19061 2635 19119 2641
rect 19061 2601 19073 2635
rect 19107 2632 19119 2635
rect 19242 2632 19248 2644
rect 19107 2604 19248 2632
rect 19107 2601 19119 2604
rect 19061 2595 19119 2601
rect 7834 2564 7840 2576
rect 7795 2536 7840 2564
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8864 2564 8892 2592
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 8864 2536 10793 2564
rect 2222 2456 2228 2508
rect 2280 2505 2286 2508
rect 2280 2499 2318 2505
rect 2306 2496 2318 2499
rect 2685 2499 2743 2505
rect 2685 2496 2697 2499
rect 2306 2468 2697 2496
rect 2306 2465 2318 2468
rect 2280 2459 2318 2465
rect 2685 2465 2697 2468
rect 2731 2496 2743 2499
rect 6086 2496 6092 2508
rect 2731 2468 6092 2496
rect 2731 2465 2743 2468
rect 2685 2459 2743 2465
rect 2280 2456 2286 2459
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7098 2496 7104 2508
rect 6779 2468 7104 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7098 2456 7104 2468
rect 7156 2496 7162 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7156 2468 7757 2496
rect 7156 2456 7162 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 7745 2459 7803 2465
rect 7760 2428 7788 2459
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 9784 2505 9812 2536
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 14553 2567 14611 2573
rect 14553 2533 14565 2567
rect 14599 2564 14611 2567
rect 14642 2564 14648 2576
rect 14599 2536 14648 2564
rect 14599 2533 14611 2536
rect 14553 2527 14611 2533
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8352 2468 8677 2496
rect 8352 2456 8358 2468
rect 8665 2465 8677 2468
rect 8711 2496 8723 2499
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8711 2468 9137 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2465 9827 2499
rect 10226 2496 10232 2508
rect 10187 2468 10232 2496
rect 9769 2459 9827 2465
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 11514 2456 11520 2508
rect 11572 2505 11578 2508
rect 12894 2505 12900 2508
rect 11572 2499 11610 2505
rect 11598 2496 11610 2499
rect 11977 2499 12035 2505
rect 11977 2496 11989 2499
rect 11598 2468 11989 2496
rect 11598 2465 11610 2468
rect 11572 2459 11610 2465
rect 11977 2465 11989 2468
rect 12023 2465 12035 2499
rect 11977 2459 12035 2465
rect 12856 2499 12900 2505
rect 12856 2465 12868 2499
rect 12952 2496 12958 2508
rect 13354 2496 13360 2508
rect 12952 2468 13360 2496
rect 12856 2459 12900 2465
rect 11572 2456 11578 2459
rect 12894 2456 12900 2459
rect 12952 2456 12958 2468
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 14461 2499 14519 2505
rect 14461 2496 14473 2499
rect 13771 2468 14473 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 14461 2465 14473 2468
rect 14507 2496 14519 2499
rect 14734 2496 14740 2508
rect 14507 2468 14740 2496
rect 14507 2465 14519 2468
rect 14461 2459 14519 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 15657 2499 15715 2505
rect 15657 2465 15669 2499
rect 15703 2465 15715 2499
rect 15657 2459 15715 2465
rect 17129 2499 17187 2505
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17129 2459 17187 2465
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 19076 2496 19104 2595
rect 19242 2592 19248 2604
rect 19300 2592 19306 2644
rect 22094 2632 22100 2644
rect 22055 2604 22100 2632
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 23750 2632 23756 2644
rect 22204 2604 23756 2632
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 19475 2536 19717 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 19705 2533 19717 2536
rect 19751 2564 19763 2567
rect 20622 2564 20628 2576
rect 19751 2536 20628 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 20901 2567 20959 2573
rect 20901 2533 20913 2567
rect 20947 2564 20959 2567
rect 21082 2564 21088 2576
rect 20947 2536 21088 2564
rect 20947 2533 20959 2536
rect 20901 2527 20959 2533
rect 21082 2524 21088 2536
rect 21140 2564 21146 2576
rect 22204 2564 22232 2604
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 25222 2632 25228 2644
rect 24320 2604 25228 2632
rect 21140 2536 22232 2564
rect 22557 2567 22615 2573
rect 21140 2524 21146 2536
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 23382 2564 23388 2576
rect 22603 2536 23388 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 23382 2524 23388 2536
rect 23440 2524 23446 2576
rect 24320 2573 24348 2604
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 26234 2592 26240 2644
rect 26292 2632 26298 2644
rect 27019 2635 27077 2641
rect 27019 2632 27031 2635
rect 26292 2604 27031 2632
rect 26292 2592 26298 2604
rect 27019 2601 27031 2604
rect 27065 2601 27077 2635
rect 29086 2632 29092 2644
rect 29047 2604 29092 2632
rect 27019 2595 27077 2601
rect 29086 2592 29092 2604
rect 29144 2592 29150 2644
rect 29454 2632 29460 2644
rect 29415 2604 29460 2632
rect 29454 2592 29460 2604
rect 29512 2592 29518 2644
rect 24305 2567 24363 2573
rect 24305 2533 24317 2567
rect 24351 2533 24363 2567
rect 24305 2527 24363 2533
rect 21266 2505 21272 2508
rect 21244 2499 21272 2505
rect 21244 2496 21256 2499
rect 18555 2468 19104 2496
rect 21179 2468 21256 2496
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 21244 2465 21256 2468
rect 21324 2496 21330 2508
rect 21637 2499 21695 2505
rect 21637 2496 21649 2499
rect 21324 2468 21649 2496
rect 21244 2459 21272 2465
rect 15194 2428 15200 2440
rect 7760 2400 8340 2428
rect 15155 2400 15200 2428
rect 8312 2372 8340 2400
rect 15194 2388 15200 2400
rect 15252 2428 15258 2440
rect 15672 2428 15700 2459
rect 15252 2400 15700 2428
rect 16301 2431 16359 2437
rect 15252 2388 15258 2400
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16666 2428 16672 2440
rect 16347 2400 16672 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16666 2388 16672 2400
rect 16724 2428 16730 2440
rect 16945 2431 17003 2437
rect 16945 2428 16957 2431
rect 16724 2400 16957 2428
rect 16724 2388 16730 2400
rect 16945 2397 16957 2400
rect 16991 2428 17003 2431
rect 17144 2428 17172 2459
rect 21266 2456 21272 2459
rect 21324 2456 21330 2468
rect 21637 2465 21649 2468
rect 21683 2465 21695 2499
rect 21637 2459 21695 2465
rect 26326 2456 26332 2508
rect 26384 2496 26390 2508
rect 26948 2499 27006 2505
rect 26948 2496 26960 2499
rect 26384 2468 26960 2496
rect 26384 2456 26390 2468
rect 26948 2465 26960 2468
rect 26994 2496 27006 2499
rect 27430 2496 27436 2508
rect 26994 2468 27436 2496
rect 26994 2465 27006 2468
rect 26948 2459 27006 2465
rect 27430 2456 27436 2468
rect 27488 2456 27494 2508
rect 27890 2456 27896 2508
rect 27948 2505 27954 2508
rect 27948 2499 27986 2505
rect 27974 2496 27986 2499
rect 28353 2499 28411 2505
rect 28353 2496 28365 2499
rect 27974 2468 28365 2496
rect 27974 2465 27986 2468
rect 27948 2459 27986 2465
rect 28353 2465 28365 2468
rect 28399 2465 28411 2499
rect 29104 2496 29132 2592
rect 29546 2524 29552 2576
rect 29604 2564 29610 2576
rect 29733 2567 29791 2573
rect 29733 2564 29745 2567
rect 29604 2536 29745 2564
rect 29604 2524 29610 2536
rect 29733 2533 29745 2536
rect 29779 2533 29791 2567
rect 29733 2527 29791 2533
rect 29822 2496 29828 2508
rect 29104 2468 29828 2496
rect 28353 2459 28411 2465
rect 27948 2456 27954 2459
rect 29822 2456 29828 2468
rect 29880 2456 29886 2508
rect 30374 2456 30380 2508
rect 30432 2496 30438 2508
rect 31332 2499 31390 2505
rect 31332 2496 31344 2499
rect 30432 2468 31344 2496
rect 30432 2456 30438 2468
rect 31332 2465 31344 2468
rect 31378 2496 31390 2499
rect 31757 2499 31815 2505
rect 31757 2496 31769 2499
rect 31378 2468 31769 2496
rect 31378 2465 31390 2468
rect 31332 2459 31390 2465
rect 31757 2465 31769 2468
rect 31803 2465 31815 2499
rect 31757 2459 31815 2465
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 16991 2400 17601 2428
rect 16991 2397 17003 2400
rect 16945 2391 17003 2397
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 19613 2431 19671 2437
rect 19613 2397 19625 2431
rect 19659 2428 19671 2431
rect 22462 2428 22468 2440
rect 19659 2400 21173 2428
rect 22423 2400 22468 2428
rect 19659 2397 19671 2400
rect 19613 2391 19671 2397
rect 8294 2320 8300 2372
rect 8352 2320 8358 2372
rect 20165 2363 20223 2369
rect 20165 2329 20177 2363
rect 20211 2360 20223 2363
rect 20254 2360 20260 2372
rect 20211 2332 20260 2360
rect 20211 2329 20223 2332
rect 20165 2323 20223 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 21145 2360 21173 2400
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 24213 2431 24271 2437
rect 24213 2397 24225 2431
rect 24259 2428 24271 2431
rect 25501 2431 25559 2437
rect 25501 2428 25513 2431
rect 24259 2400 25513 2428
rect 24259 2397 24271 2400
rect 24213 2391 24271 2397
rect 25501 2397 25513 2400
rect 25547 2428 25559 2431
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25547 2400 25697 2428
rect 25547 2397 25559 2400
rect 25501 2391 25559 2397
rect 25685 2397 25697 2400
rect 25731 2397 25743 2431
rect 25685 2391 25743 2397
rect 21358 2369 21364 2372
rect 21315 2363 21364 2369
rect 21315 2360 21327 2363
rect 21145 2332 21327 2360
rect 21315 2329 21327 2332
rect 21361 2329 21364 2363
rect 21315 2323 21364 2329
rect 21358 2320 21364 2323
rect 21416 2360 21422 2372
rect 23017 2363 23075 2369
rect 21416 2332 21463 2360
rect 21416 2320 21422 2332
rect 23017 2329 23029 2363
rect 23063 2360 23075 2363
rect 24762 2360 24768 2372
rect 23063 2332 24768 2360
rect 23063 2329 23075 2332
rect 23017 2323 23075 2329
rect 24762 2320 24768 2332
rect 24820 2320 24826 2372
rect 26234 2320 26240 2372
rect 26292 2360 26298 2372
rect 26292 2332 26337 2360
rect 26292 2320 26298 2332
rect 26510 2292 26516 2304
rect 26471 2264 26516 2292
rect 26510 2252 26516 2264
rect 26568 2252 26574 2304
rect 27430 2292 27436 2304
rect 27391 2264 27436 2292
rect 27430 2252 27436 2264
rect 27488 2252 27494 2304
rect 28031 2295 28089 2301
rect 28031 2261 28043 2295
rect 28077 2292 28089 2295
rect 28902 2292 28908 2304
rect 28077 2264 28908 2292
rect 28077 2261 28089 2264
rect 28031 2255 28089 2261
rect 28902 2252 28908 2264
rect 28960 2252 28966 2304
rect 31435 2295 31493 2301
rect 31435 2261 31447 2295
rect 31481 2292 31493 2295
rect 31662 2292 31668 2304
rect 31481 2264 31668 2292
rect 31481 2261 31493 2264
rect 31435 2255 31493 2261
rect 31662 2252 31668 2264
rect 31720 2252 31726 2304
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 18046 552 18052 604
rect 18104 592 18110 604
rect 18322 592 18328 604
rect 18104 564 18328 592
rect 18104 552 18110 564
rect 18322 552 18328 564
rect 18380 552 18386 604
<< via1 >>
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 1676 13336 1728 13388
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 1492 12928 1544 12980
rect 1676 12928 1728 12980
rect 9128 12928 9180 12980
rect 2136 12588 2188 12640
rect 3792 12588 3844 12640
rect 5816 12588 5868 12640
rect 24584 12588 24636 12640
rect 24952 12588 25004 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 35624 12427 35676 12436
rect 35624 12393 35633 12427
rect 35633 12393 35667 12427
rect 35667 12393 35676 12427
rect 35624 12384 35676 12393
rect 2044 12248 2096 12300
rect 3148 12248 3200 12300
rect 11336 12248 11388 12300
rect 19432 12248 19484 12300
rect 24124 12291 24176 12300
rect 24124 12257 24142 12291
rect 24142 12257 24176 12291
rect 24124 12248 24176 12257
rect 25228 12248 25280 12300
rect 34612 12248 34664 12300
rect 35440 12291 35492 12300
rect 35440 12257 35449 12291
rect 35449 12257 35483 12291
rect 35483 12257 35492 12291
rect 35440 12248 35492 12257
rect 29552 12223 29604 12232
rect 29552 12189 29561 12223
rect 29561 12189 29595 12223
rect 29595 12189 29604 12223
rect 29552 12180 29604 12189
rect 2320 12044 2372 12096
rect 2780 12044 2832 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 11428 12044 11480 12096
rect 19340 12087 19392 12096
rect 19340 12053 19349 12087
rect 19349 12053 19383 12087
rect 19383 12053 19392 12087
rect 19340 12044 19392 12053
rect 24400 12044 24452 12096
rect 24860 12044 24912 12096
rect 34152 12044 34204 12096
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 22468 11840 22520 11892
rect 2044 11815 2096 11824
rect 2044 11781 2053 11815
rect 2053 11781 2087 11815
rect 2087 11781 2096 11815
rect 2044 11772 2096 11781
rect 19524 11772 19576 11824
rect 2228 11704 2280 11756
rect 9680 11704 9732 11756
rect 10140 11704 10192 11756
rect 10968 11704 11020 11756
rect 18604 11679 18656 11688
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 2412 11500 2464 11509
rect 2596 11500 2648 11552
rect 3148 11500 3200 11552
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 10784 11611 10836 11620
rect 10784 11577 10793 11611
rect 10793 11577 10827 11611
rect 10827 11577 10836 11611
rect 10784 11568 10836 11577
rect 10692 11500 10744 11552
rect 11336 11500 11388 11552
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 19708 11543 19760 11552
rect 19708 11509 19717 11543
rect 19717 11509 19751 11543
rect 19751 11509 19760 11543
rect 19708 11500 19760 11509
rect 24308 11636 24360 11688
rect 30104 11679 30156 11688
rect 30104 11645 30122 11679
rect 30122 11645 30156 11679
rect 30104 11636 30156 11645
rect 35440 11840 35492 11892
rect 35716 11840 35768 11892
rect 37188 11840 37240 11892
rect 33416 11772 33468 11824
rect 33876 11679 33928 11688
rect 33876 11645 33894 11679
rect 33894 11645 33928 11679
rect 33876 11636 33928 11645
rect 35348 11636 35400 11688
rect 36544 11679 36596 11688
rect 36544 11645 36588 11679
rect 36588 11645 36596 11679
rect 36544 11636 36596 11645
rect 21640 11500 21692 11552
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 24676 11500 24728 11552
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 25412 11543 25464 11552
rect 25412 11509 25421 11543
rect 25421 11509 25455 11543
rect 25455 11509 25464 11543
rect 25412 11500 25464 11509
rect 30288 11500 30340 11552
rect 31484 11500 31536 11552
rect 32036 11568 32088 11620
rect 34612 11611 34664 11620
rect 34612 11577 34621 11611
rect 34621 11577 34655 11611
rect 34655 11577 34664 11611
rect 34612 11568 34664 11577
rect 33784 11500 33836 11552
rect 34060 11500 34112 11552
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 10140 11339 10192 11348
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 27436 11296 27488 11348
rect 31484 11339 31536 11348
rect 31484 11305 31493 11339
rect 31493 11305 31527 11339
rect 31527 11305 31536 11339
rect 31484 11296 31536 11305
rect 35624 11339 35676 11348
rect 35624 11305 35633 11339
rect 35633 11305 35667 11339
rect 35667 11305 35676 11339
rect 35624 11296 35676 11305
rect 11612 11271 11664 11280
rect 11612 11237 11621 11271
rect 11621 11237 11655 11271
rect 11655 11237 11664 11271
rect 11612 11228 11664 11237
rect 20812 11228 20864 11280
rect 24400 11271 24452 11280
rect 24400 11237 24409 11271
rect 24409 11237 24443 11271
rect 24443 11237 24452 11271
rect 24400 11228 24452 11237
rect 24492 11271 24544 11280
rect 24492 11237 24501 11271
rect 24501 11237 24535 11271
rect 24535 11237 24544 11271
rect 24492 11228 24544 11237
rect 29552 11228 29604 11280
rect 29920 11271 29972 11280
rect 29920 11237 29929 11271
rect 29929 11237 29963 11271
rect 29963 11237 29972 11271
rect 30472 11271 30524 11280
rect 29920 11228 29972 11237
rect 30472 11237 30481 11271
rect 30481 11237 30515 11271
rect 30515 11237 30524 11271
rect 30472 11228 30524 11237
rect 33508 11228 33560 11280
rect 1676 11160 1728 11212
rect 4804 11160 4856 11212
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10692 11160 10744 11212
rect 13452 11160 13504 11212
rect 11520 11135 11572 11144
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 11520 11101 11529 11135
rect 11529 11101 11563 11135
rect 11563 11101 11572 11135
rect 11520 11092 11572 11101
rect 15568 11160 15620 11212
rect 18236 11203 18288 11212
rect 18236 11169 18254 11203
rect 18254 11169 18288 11203
rect 18236 11160 18288 11169
rect 19340 11203 19392 11212
rect 19340 11169 19349 11203
rect 19349 11169 19383 11203
rect 19383 11169 19392 11203
rect 19340 11160 19392 11169
rect 19524 11160 19576 11212
rect 23388 11203 23440 11212
rect 23388 11169 23406 11203
rect 23406 11169 23440 11203
rect 23388 11160 23440 11169
rect 27068 11160 27120 11212
rect 28080 11203 28132 11212
rect 28080 11169 28089 11203
rect 28089 11169 28123 11203
rect 28123 11169 28132 11203
rect 28080 11160 28132 11169
rect 4252 11024 4304 11076
rect 10048 11024 10100 11076
rect 11152 11024 11204 11076
rect 16120 11092 16172 11144
rect 13176 11067 13228 11076
rect 13176 11033 13185 11067
rect 13185 11033 13219 11067
rect 13219 11033 13228 11067
rect 13176 11024 13228 11033
rect 17960 11024 18012 11076
rect 21456 11092 21508 11144
rect 21640 11135 21692 11144
rect 21640 11101 21649 11135
rect 21649 11101 21683 11135
rect 21683 11101 21692 11135
rect 21640 11092 21692 11101
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 31760 11160 31812 11212
rect 32404 11160 32456 11212
rect 33968 11160 34020 11212
rect 35440 11203 35492 11212
rect 35440 11169 35449 11203
rect 35449 11169 35483 11203
rect 35483 11169 35492 11203
rect 35440 11160 35492 11169
rect 35900 11160 35952 11212
rect 37004 11160 37056 11212
rect 21272 11024 21324 11076
rect 28908 11092 28960 11144
rect 32680 11135 32732 11144
rect 32680 11101 32689 11135
rect 32689 11101 32723 11135
rect 32723 11101 32732 11135
rect 32680 11092 32732 11101
rect 35072 11092 35124 11144
rect 36728 11067 36780 11076
rect 36728 11033 36737 11067
rect 36737 11033 36771 11067
rect 36771 11033 36780 11067
rect 36728 11024 36780 11033
rect 3424 10956 3476 11008
rect 10232 10956 10284 11008
rect 12716 10956 12768 11008
rect 20168 10999 20220 11008
rect 20168 10965 20177 10999
rect 20177 10965 20211 10999
rect 20211 10965 20220 10999
rect 20168 10956 20220 10965
rect 23204 10956 23256 11008
rect 27620 10999 27672 11008
rect 27620 10965 27629 10999
rect 27629 10965 27663 10999
rect 27663 10965 27672 10999
rect 27620 10956 27672 10965
rect 34796 10956 34848 11008
rect 34980 10956 35032 11008
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 4804 10795 4856 10804
rect 4804 10761 4813 10795
rect 4813 10761 4847 10795
rect 4847 10761 4856 10795
rect 4804 10752 4856 10761
rect 8576 10752 8628 10804
rect 11612 10752 11664 10804
rect 17500 10752 17552 10804
rect 19340 10752 19392 10804
rect 21364 10752 21416 10804
rect 21732 10795 21784 10804
rect 21732 10761 21741 10795
rect 21741 10761 21775 10795
rect 21775 10761 21784 10795
rect 21732 10752 21784 10761
rect 23112 10795 23164 10804
rect 23112 10761 23121 10795
rect 23121 10761 23155 10795
rect 23155 10761 23164 10795
rect 23112 10752 23164 10761
rect 24400 10752 24452 10804
rect 27068 10795 27120 10804
rect 27068 10761 27077 10795
rect 27077 10761 27111 10795
rect 27111 10761 27120 10795
rect 27068 10752 27120 10761
rect 29552 10752 29604 10804
rect 33232 10752 33284 10804
rect 33968 10752 34020 10804
rect 35900 10795 35952 10804
rect 35900 10761 35909 10795
rect 35909 10761 35943 10795
rect 35943 10761 35952 10795
rect 35900 10752 35952 10761
rect 36636 10795 36688 10804
rect 36636 10761 36645 10795
rect 36645 10761 36679 10795
rect 36679 10761 36688 10795
rect 36636 10752 36688 10761
rect 37004 10795 37056 10804
rect 37004 10761 37013 10795
rect 37013 10761 37047 10795
rect 37047 10761 37056 10795
rect 37004 10752 37056 10761
rect 9588 10684 9640 10736
rect 29460 10684 29512 10736
rect 29920 10684 29972 10736
rect 31484 10684 31536 10736
rect 34060 10684 34112 10736
rect 11520 10616 11572 10668
rect 14924 10616 14976 10668
rect 16212 10616 16264 10668
rect 19708 10616 19760 10668
rect 20076 10659 20128 10668
rect 20076 10625 20085 10659
rect 20085 10625 20119 10659
rect 20119 10625 20128 10659
rect 20076 10616 20128 10625
rect 21640 10616 21692 10668
rect 24584 10659 24636 10668
rect 24584 10625 24593 10659
rect 24593 10625 24627 10659
rect 24627 10625 24636 10659
rect 24584 10616 24636 10625
rect 2136 10548 2188 10600
rect 3056 10591 3108 10600
rect 3056 10557 3065 10591
rect 3065 10557 3099 10591
rect 3099 10557 3108 10591
rect 3056 10548 3108 10557
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2688 10412 2740 10464
rect 3424 10455 3476 10464
rect 3424 10421 3433 10455
rect 3433 10421 3467 10455
rect 3467 10421 3476 10455
rect 3424 10412 3476 10421
rect 4068 10412 4120 10464
rect 4712 10412 4764 10464
rect 6552 10412 6604 10464
rect 9128 10548 9180 10600
rect 9956 10548 10008 10600
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 10232 10523 10284 10532
rect 10232 10489 10241 10523
rect 10241 10489 10275 10523
rect 10275 10489 10284 10523
rect 10232 10480 10284 10489
rect 10324 10523 10376 10532
rect 10324 10489 10333 10523
rect 10333 10489 10367 10523
rect 10367 10489 10376 10523
rect 10324 10480 10376 10489
rect 11152 10480 11204 10532
rect 14188 10548 14240 10600
rect 17684 10548 17736 10600
rect 21548 10591 21600 10600
rect 15108 10523 15160 10532
rect 9220 10412 9272 10464
rect 10692 10412 10744 10464
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 16120 10523 16172 10532
rect 15200 10480 15252 10489
rect 16120 10489 16129 10523
rect 16129 10489 16163 10523
rect 16163 10489 16172 10523
rect 16120 10480 16172 10489
rect 12348 10412 12400 10464
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 14832 10412 14884 10464
rect 18236 10455 18288 10464
rect 18236 10421 18245 10455
rect 18245 10421 18279 10455
rect 18279 10421 18288 10455
rect 18236 10412 18288 10421
rect 21548 10557 21557 10591
rect 21557 10557 21591 10591
rect 21591 10557 21600 10591
rect 21548 10548 21600 10557
rect 22192 10548 22244 10600
rect 23112 10548 23164 10600
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26148 10548 26200 10600
rect 29276 10616 29328 10668
rect 30472 10659 30524 10668
rect 30472 10625 30481 10659
rect 30481 10625 30515 10659
rect 30515 10625 30524 10659
rect 30472 10616 30524 10625
rect 32404 10616 32456 10668
rect 27712 10548 27764 10600
rect 27988 10548 28040 10600
rect 19156 10523 19208 10532
rect 19156 10489 19165 10523
rect 19165 10489 19199 10523
rect 19199 10489 19208 10523
rect 19156 10480 19208 10489
rect 20168 10523 20220 10532
rect 20168 10489 20177 10523
rect 20177 10489 20211 10523
rect 20211 10489 20220 10523
rect 20168 10480 20220 10489
rect 24584 10480 24636 10532
rect 25044 10480 25096 10532
rect 28356 10523 28408 10532
rect 28356 10489 28365 10523
rect 28365 10489 28399 10523
rect 28399 10489 28408 10523
rect 28356 10480 28408 10489
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 20812 10412 20864 10464
rect 21456 10455 21508 10464
rect 21456 10421 21465 10455
rect 21465 10421 21499 10455
rect 21499 10421 21508 10455
rect 21456 10412 21508 10421
rect 22928 10412 22980 10464
rect 23572 10412 23624 10464
rect 24400 10455 24452 10464
rect 24400 10421 24409 10455
rect 24409 10421 24443 10455
rect 24443 10421 24452 10455
rect 24400 10412 24452 10421
rect 26240 10412 26292 10464
rect 28080 10412 28132 10464
rect 30104 10523 30156 10532
rect 30104 10489 30113 10523
rect 30113 10489 30147 10523
rect 30147 10489 30156 10523
rect 30104 10480 30156 10489
rect 30472 10480 30524 10532
rect 31116 10412 31168 10464
rect 31576 10480 31628 10532
rect 32220 10523 32272 10532
rect 32220 10489 32229 10523
rect 32229 10489 32263 10523
rect 32263 10489 32272 10523
rect 32220 10480 32272 10489
rect 34060 10480 34112 10532
rect 34980 10523 35032 10532
rect 34980 10489 34989 10523
rect 34989 10489 35023 10523
rect 35023 10489 35032 10523
rect 34980 10480 35032 10489
rect 35072 10523 35124 10532
rect 35072 10489 35081 10523
rect 35081 10489 35115 10523
rect 35115 10489 35124 10523
rect 35072 10480 35124 10489
rect 35808 10480 35860 10532
rect 31760 10412 31812 10464
rect 32404 10412 32456 10464
rect 32864 10455 32916 10464
rect 32864 10421 32873 10455
rect 32873 10421 32907 10455
rect 32907 10421 32916 10455
rect 32864 10412 32916 10421
rect 36084 10412 36136 10464
rect 37280 10412 37332 10464
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 1768 10208 1820 10260
rect 4160 10208 4212 10260
rect 10048 10208 10100 10260
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 10968 10208 11020 10260
rect 11612 10208 11664 10260
rect 10600 10183 10652 10192
rect 10600 10149 10609 10183
rect 10609 10149 10643 10183
rect 10643 10149 10652 10183
rect 10600 10140 10652 10149
rect 11428 10140 11480 10192
rect 13084 10208 13136 10260
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15568 10251 15620 10260
rect 15568 10217 15577 10251
rect 15577 10217 15611 10251
rect 15611 10217 15620 10251
rect 15568 10208 15620 10217
rect 19156 10208 19208 10260
rect 19432 10251 19484 10260
rect 19432 10217 19441 10251
rect 19441 10217 19475 10251
rect 19475 10217 19484 10251
rect 19432 10208 19484 10217
rect 20076 10208 20128 10260
rect 26148 10251 26200 10260
rect 26148 10217 26157 10251
rect 26157 10217 26191 10251
rect 26191 10217 26200 10251
rect 26148 10208 26200 10217
rect 26516 10208 26568 10260
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 5172 10072 5224 10124
rect 7380 10072 7432 10124
rect 8392 10072 8444 10124
rect 14188 10115 14240 10124
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 6736 10004 6788 10056
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 14188 10081 14197 10115
rect 14197 10081 14231 10115
rect 14231 10081 14240 10115
rect 15660 10140 15712 10192
rect 16580 10140 16632 10192
rect 21916 10140 21968 10192
rect 23204 10183 23256 10192
rect 23204 10149 23213 10183
rect 23213 10149 23247 10183
rect 23247 10149 23256 10183
rect 23204 10140 23256 10149
rect 23296 10183 23348 10192
rect 23296 10149 23305 10183
rect 23305 10149 23339 10183
rect 23339 10149 23348 10183
rect 23296 10140 23348 10149
rect 24584 10140 24636 10192
rect 24768 10183 24820 10192
rect 24768 10149 24777 10183
rect 24777 10149 24811 10183
rect 24811 10149 24820 10183
rect 24768 10140 24820 10149
rect 24952 10140 25004 10192
rect 26608 10183 26660 10192
rect 26608 10149 26617 10183
rect 26617 10149 26651 10183
rect 26651 10149 26660 10183
rect 26608 10140 26660 10149
rect 27988 10208 28040 10260
rect 29460 10251 29512 10260
rect 29460 10217 29469 10251
rect 29469 10217 29503 10251
rect 29503 10217 29512 10251
rect 29460 10208 29512 10217
rect 30380 10208 30432 10260
rect 31576 10251 31628 10260
rect 28816 10140 28868 10192
rect 29000 10140 29052 10192
rect 31576 10217 31585 10251
rect 31585 10217 31619 10251
rect 31619 10217 31628 10251
rect 31576 10208 31628 10217
rect 32680 10251 32732 10260
rect 32680 10217 32689 10251
rect 32689 10217 32723 10251
rect 32723 10217 32732 10251
rect 32680 10208 32732 10217
rect 30564 10183 30616 10192
rect 30564 10149 30573 10183
rect 30573 10149 30607 10183
rect 30607 10149 30616 10183
rect 33140 10183 33192 10192
rect 30564 10140 30616 10149
rect 33140 10149 33149 10183
rect 33149 10149 33183 10183
rect 33183 10149 33192 10183
rect 33140 10140 33192 10149
rect 33692 10183 33744 10192
rect 33692 10149 33701 10183
rect 33701 10149 33735 10183
rect 33735 10149 33744 10183
rect 33692 10140 33744 10149
rect 17592 10115 17644 10124
rect 14188 10072 14240 10081
rect 17592 10081 17601 10115
rect 17601 10081 17635 10115
rect 17635 10081 17644 10115
rect 17592 10072 17644 10081
rect 17868 10072 17920 10124
rect 19340 10115 19392 10124
rect 14096 10004 14148 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 16212 10047 16264 10056
rect 16212 10013 16221 10047
rect 16221 10013 16255 10047
rect 16255 10013 16264 10047
rect 16212 10004 16264 10013
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19524 10072 19576 10124
rect 19984 10072 20036 10124
rect 21640 10115 21692 10124
rect 21640 10081 21649 10115
rect 21649 10081 21683 10115
rect 21683 10081 21692 10115
rect 21640 10072 21692 10081
rect 19248 10004 19300 10056
rect 20720 10004 20772 10056
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 25044 10047 25096 10056
rect 25044 10013 25053 10047
rect 25053 10013 25087 10047
rect 25087 10013 25096 10047
rect 25044 10004 25096 10013
rect 26884 10047 26936 10056
rect 26884 10013 26893 10047
rect 26893 10013 26927 10047
rect 26927 10013 26936 10047
rect 26884 10004 26936 10013
rect 28540 10047 28592 10056
rect 28540 10013 28549 10047
rect 28549 10013 28583 10047
rect 28583 10013 28592 10047
rect 28540 10004 28592 10013
rect 31116 10047 31168 10056
rect 31116 10013 31125 10047
rect 31125 10013 31159 10047
rect 31159 10013 31168 10047
rect 31116 10004 31168 10013
rect 32220 10004 32272 10056
rect 35808 10208 35860 10260
rect 36360 10208 36412 10260
rect 36452 10208 36504 10260
rect 34704 10183 34756 10192
rect 34704 10149 34713 10183
rect 34713 10149 34747 10183
rect 34747 10149 34756 10183
rect 34704 10140 34756 10149
rect 36084 10115 36136 10124
rect 36084 10081 36093 10115
rect 36093 10081 36127 10115
rect 36127 10081 36136 10115
rect 36084 10072 36136 10081
rect 34612 10047 34664 10056
rect 34612 10013 34621 10047
rect 34621 10013 34655 10047
rect 34655 10013 34664 10047
rect 34612 10004 34664 10013
rect 34888 10047 34940 10056
rect 34888 10013 34897 10047
rect 34897 10013 34931 10047
rect 34931 10013 34940 10047
rect 34888 10004 34940 10013
rect 9680 9936 9732 9988
rect 18788 9936 18840 9988
rect 8208 9868 8260 9920
rect 8852 9868 8904 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 24124 9911 24176 9920
rect 24124 9877 24133 9911
rect 24133 9877 24167 9911
rect 24167 9877 24176 9911
rect 24124 9868 24176 9877
rect 30104 9911 30156 9920
rect 30104 9877 30113 9911
rect 30113 9877 30147 9911
rect 30147 9877 30156 9911
rect 30104 9868 30156 9877
rect 32404 9911 32456 9920
rect 32404 9877 32413 9911
rect 32413 9877 32447 9911
rect 32447 9877 32456 9911
rect 32404 9868 32456 9877
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 5172 9707 5224 9716
rect 5172 9673 5181 9707
rect 5181 9673 5215 9707
rect 5215 9673 5224 9707
rect 5172 9664 5224 9673
rect 8852 9664 8904 9716
rect 10508 9664 10560 9716
rect 11428 9707 11480 9716
rect 11428 9673 11437 9707
rect 11437 9673 11471 9707
rect 11471 9673 11480 9707
rect 11428 9664 11480 9673
rect 11612 9664 11664 9716
rect 14188 9664 14240 9716
rect 15660 9664 15712 9716
rect 18788 9707 18840 9716
rect 18788 9673 18797 9707
rect 18797 9673 18831 9707
rect 18831 9673 18840 9707
rect 18788 9664 18840 9673
rect 20168 9707 20220 9716
rect 20168 9673 20177 9707
rect 20177 9673 20211 9707
rect 20211 9673 20220 9707
rect 20168 9664 20220 9673
rect 21916 9707 21968 9716
rect 21916 9673 21925 9707
rect 21925 9673 21959 9707
rect 21959 9673 21968 9707
rect 21916 9664 21968 9673
rect 23204 9664 23256 9716
rect 23480 9664 23532 9716
rect 24952 9707 25004 9716
rect 2412 9596 2464 9648
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 5908 9596 5960 9648
rect 11060 9639 11112 9648
rect 11060 9605 11069 9639
rect 11069 9605 11103 9639
rect 11103 9605 11112 9639
rect 11060 9596 11112 9605
rect 12624 9596 12676 9648
rect 13084 9639 13136 9648
rect 13084 9605 13093 9639
rect 13093 9605 13127 9639
rect 13127 9605 13136 9639
rect 13084 9596 13136 9605
rect 15200 9596 15252 9648
rect 16580 9639 16632 9648
rect 16580 9605 16589 9639
rect 16589 9605 16623 9639
rect 16623 9605 16632 9639
rect 16580 9596 16632 9605
rect 17132 9596 17184 9648
rect 17868 9639 17920 9648
rect 17868 9605 17877 9639
rect 17877 9605 17911 9639
rect 17911 9605 17920 9639
rect 17868 9596 17920 9605
rect 9036 9528 9088 9580
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 14372 9528 14424 9580
rect 15016 9571 15068 9580
rect 15016 9537 15025 9571
rect 15025 9537 15059 9571
rect 15059 9537 15068 9571
rect 15016 9528 15068 9537
rect 19156 9528 19208 9580
rect 21272 9528 21324 9580
rect 23296 9596 23348 9648
rect 24952 9673 24961 9707
rect 24961 9673 24995 9707
rect 24995 9673 25004 9707
rect 24952 9664 25004 9673
rect 26884 9664 26936 9716
rect 30380 9664 30432 9716
rect 33140 9664 33192 9716
rect 24676 9528 24728 9580
rect 25504 9571 25556 9580
rect 25504 9537 25513 9571
rect 25513 9537 25547 9571
rect 25547 9537 25556 9571
rect 25504 9528 25556 9537
rect 27988 9596 28040 9648
rect 28816 9596 28868 9648
rect 4528 9460 4580 9512
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 5632 9503 5684 9512
rect 4620 9460 4672 9469
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 3332 9392 3384 9444
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 13544 9460 13596 9512
rect 16948 9503 17000 9512
rect 16948 9469 16992 9503
rect 16992 9469 17000 9503
rect 17408 9503 17460 9512
rect 16948 9460 17000 9469
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 18788 9460 18840 9512
rect 23020 9460 23072 9512
rect 24124 9460 24176 9512
rect 28540 9528 28592 9580
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 2136 9324 2188 9376
rect 4160 9324 4212 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6828 9324 6880 9376
rect 7380 9324 7432 9376
rect 7840 9367 7892 9376
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 9772 9324 9824 9376
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 15936 9392 15988 9444
rect 13912 9324 13964 9376
rect 17316 9324 17368 9376
rect 18696 9324 18748 9376
rect 19156 9367 19208 9376
rect 19156 9333 19165 9367
rect 19165 9333 19199 9367
rect 19199 9333 19208 9367
rect 19156 9324 19208 9333
rect 19340 9324 19392 9376
rect 19800 9324 19852 9376
rect 21456 9324 21508 9376
rect 23664 9324 23716 9376
rect 24952 9324 25004 9376
rect 28172 9392 28224 9444
rect 30564 9639 30616 9648
rect 30564 9605 30573 9639
rect 30573 9605 30607 9639
rect 30607 9605 30616 9639
rect 30564 9596 30616 9605
rect 31484 9596 31536 9648
rect 34612 9664 34664 9716
rect 34888 9596 34940 9648
rect 29000 9528 29052 9580
rect 32680 9528 32732 9580
rect 34152 9528 34204 9580
rect 35164 9528 35216 9580
rect 35900 9528 35952 9580
rect 30748 9460 30800 9512
rect 33048 9460 33100 9512
rect 36084 9503 36136 9512
rect 36084 9469 36093 9503
rect 36093 9469 36127 9503
rect 36127 9469 36136 9503
rect 36084 9460 36136 9469
rect 29184 9392 29236 9444
rect 32680 9435 32732 9444
rect 32680 9401 32683 9435
rect 32683 9401 32717 9435
rect 32717 9401 32732 9435
rect 32680 9392 32732 9401
rect 35072 9435 35124 9444
rect 35072 9401 35081 9435
rect 35081 9401 35115 9435
rect 35115 9401 35124 9435
rect 35072 9392 35124 9401
rect 36360 9392 36412 9444
rect 36544 9435 36596 9444
rect 36544 9401 36553 9435
rect 36553 9401 36587 9435
rect 36587 9401 36596 9435
rect 36544 9392 36596 9401
rect 36728 9392 36780 9444
rect 26516 9367 26568 9376
rect 26516 9333 26525 9367
rect 26525 9333 26559 9367
rect 26559 9333 26568 9367
rect 26516 9324 26568 9333
rect 34336 9367 34388 9376
rect 34336 9333 34345 9367
rect 34345 9333 34379 9367
rect 34379 9333 34388 9367
rect 34336 9324 34388 9333
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 6920 9120 6972 9172
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 10784 9120 10836 9172
rect 11612 9120 11664 9172
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 16580 9120 16632 9172
rect 17592 9163 17644 9172
rect 17592 9129 17601 9163
rect 17601 9129 17635 9163
rect 17635 9129 17644 9163
rect 17592 9120 17644 9129
rect 18696 9163 18748 9172
rect 18696 9129 18705 9163
rect 18705 9129 18739 9163
rect 18739 9129 18748 9163
rect 20720 9163 20772 9172
rect 18696 9120 18748 9129
rect 2596 9095 2648 9104
rect 2596 9061 2605 9095
rect 2605 9061 2639 9095
rect 2639 9061 2648 9095
rect 2596 9052 2648 9061
rect 5080 9095 5132 9104
rect 5080 9061 5089 9095
rect 5089 9061 5123 9095
rect 5123 9061 5132 9095
rect 5080 9052 5132 9061
rect 6552 9095 6604 9104
rect 6552 9061 6561 9095
rect 6561 9061 6595 9095
rect 6595 9061 6604 9095
rect 6552 9052 6604 9061
rect 6644 9095 6696 9104
rect 6644 9061 6653 9095
rect 6653 9061 6687 9095
rect 6687 9061 6696 9095
rect 6644 9052 6696 9061
rect 10232 9052 10284 9104
rect 11244 9052 11296 9104
rect 13820 9095 13872 9104
rect 13820 9061 13829 9095
rect 13829 9061 13863 9095
rect 13863 9061 13872 9095
rect 13820 9052 13872 9061
rect 14924 9052 14976 9104
rect 15936 9052 15988 9104
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 21272 9120 21324 9172
rect 24860 9120 24912 9172
rect 25136 9120 25188 9172
rect 28540 9163 28592 9172
rect 28540 9129 28549 9163
rect 28549 9129 28583 9163
rect 28583 9129 28592 9163
rect 28540 9120 28592 9129
rect 30104 9120 30156 9172
rect 35164 9120 35216 9172
rect 36360 9163 36412 9172
rect 36360 9129 36369 9163
rect 36369 9129 36403 9163
rect 36403 9129 36412 9163
rect 36360 9120 36412 9129
rect 36728 9163 36780 9172
rect 36728 9129 36737 9163
rect 36737 9129 36771 9163
rect 36771 9129 36780 9163
rect 36728 9120 36780 9129
rect 19064 9095 19116 9104
rect 19064 9061 19073 9095
rect 19073 9061 19107 9095
rect 19107 9061 19116 9095
rect 23020 9095 23072 9104
rect 19064 9052 19116 9061
rect 23020 9061 23029 9095
rect 23029 9061 23063 9095
rect 23063 9061 23072 9095
rect 23020 9052 23072 9061
rect 23664 9052 23716 9104
rect 25504 9095 25556 9104
rect 25504 9061 25513 9095
rect 25513 9061 25547 9095
rect 25547 9061 25556 9095
rect 25504 9052 25556 9061
rect 29184 9052 29236 9104
rect 32772 9052 32824 9104
rect 34152 9052 34204 9104
rect 35900 9052 35952 9104
rect 1492 9027 1544 9036
rect 1492 8993 1510 9027
rect 1510 8993 1544 9027
rect 1492 8984 1544 8993
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8116 8984 8168 8993
rect 8300 8984 8352 9036
rect 9680 9027 9732 9036
rect 9680 8993 9724 9027
rect 9724 8993 9732 9027
rect 9680 8984 9732 8993
rect 12348 8984 12400 9036
rect 15752 9027 15804 9036
rect 15752 8993 15761 9027
rect 15761 8993 15795 9027
rect 15795 8993 15804 9027
rect 15752 8984 15804 8993
rect 17868 9027 17920 9036
rect 17868 8993 17912 9027
rect 17912 8993 17920 9027
rect 17868 8984 17920 8993
rect 20720 8984 20772 9036
rect 21272 8984 21324 9036
rect 22560 9027 22612 9036
rect 22560 8993 22569 9027
rect 22569 8993 22603 9027
rect 22603 8993 22612 9027
rect 22560 8984 22612 8993
rect 22744 9027 22796 9036
rect 22744 8993 22753 9027
rect 22753 8993 22787 9027
rect 22787 8993 22796 9027
rect 22744 8984 22796 8993
rect 24952 8984 25004 9036
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 26976 9027 27028 9036
rect 26976 8993 26985 9027
rect 26985 8993 27019 9027
rect 27019 8993 27028 9027
rect 26976 8984 27028 8993
rect 28356 8984 28408 9036
rect 30472 9027 30524 9036
rect 30472 8993 30481 9027
rect 30481 8993 30515 9027
rect 30515 8993 30524 9027
rect 30472 8984 30524 8993
rect 30932 9027 30984 9036
rect 30932 8993 30941 9027
rect 30941 8993 30975 9027
rect 30975 8993 30984 9027
rect 30932 8984 30984 8993
rect 32128 9027 32180 9036
rect 32128 8993 32137 9027
rect 32137 8993 32171 9027
rect 32171 8993 32180 9027
rect 32128 8984 32180 8993
rect 32404 8984 32456 9036
rect 34336 8984 34388 9036
rect 34704 8984 34756 9036
rect 2688 8916 2740 8968
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 4804 8916 4856 8968
rect 5172 8916 5224 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 25136 8916 25188 8968
rect 26608 8916 26660 8968
rect 34060 8916 34112 8968
rect 36268 8916 36320 8968
rect 18972 8848 19024 8900
rect 19524 8891 19576 8900
rect 19524 8857 19533 8891
rect 19533 8857 19567 8891
rect 19567 8857 19576 8891
rect 19524 8848 19576 8857
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 8760 8780 8812 8832
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 14096 8780 14148 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 20720 8780 20772 8832
rect 21548 8823 21600 8832
rect 21548 8789 21557 8823
rect 21557 8789 21591 8823
rect 21591 8789 21600 8823
rect 21548 8780 21600 8789
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 27712 8823 27764 8832
rect 27712 8789 27721 8823
rect 27721 8789 27755 8823
rect 27755 8789 27764 8823
rect 27712 8780 27764 8789
rect 30196 8780 30248 8832
rect 34704 8780 34756 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1492 8576 1544 8628
rect 2596 8576 2648 8628
rect 3148 8576 3200 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 6552 8576 6604 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8300 8576 8352 8628
rect 9036 8576 9088 8628
rect 9680 8576 9732 8628
rect 10600 8576 10652 8628
rect 12348 8576 12400 8628
rect 13820 8576 13872 8628
rect 15752 8576 15804 8628
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 19432 8576 19484 8628
rect 20812 8576 20864 8628
rect 21364 8619 21416 8628
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 22744 8576 22796 8628
rect 23480 8576 23532 8628
rect 24400 8576 24452 8628
rect 25136 8576 25188 8628
rect 25412 8576 25464 8628
rect 2872 8551 2924 8560
rect 2872 8517 2881 8551
rect 2881 8517 2915 8551
rect 2915 8517 2924 8551
rect 2872 8508 2924 8517
rect 5172 8508 5224 8560
rect 1860 8440 1912 8492
rect 2688 8440 2740 8492
rect 5356 8440 5408 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 10784 8440 10836 8492
rect 12808 8483 12860 8492
rect 12808 8449 12817 8483
rect 12817 8449 12851 8483
rect 12851 8449 12860 8483
rect 12808 8440 12860 8449
rect 16028 8508 16080 8560
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 8852 8372 8904 8424
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 14648 8372 14700 8424
rect 16028 8372 16080 8424
rect 16948 8372 17000 8424
rect 2320 8304 2372 8356
rect 2688 8304 2740 8356
rect 3332 8304 3384 8356
rect 4896 8236 4948 8288
rect 5356 8347 5408 8356
rect 5356 8313 5365 8347
rect 5365 8313 5399 8347
rect 5399 8313 5408 8347
rect 5356 8304 5408 8313
rect 7196 8304 7248 8356
rect 9772 8304 9824 8356
rect 11244 8347 11296 8356
rect 11244 8313 11253 8347
rect 11253 8313 11287 8347
rect 11287 8313 11296 8347
rect 11244 8304 11296 8313
rect 17040 8347 17092 8356
rect 17040 8313 17049 8347
rect 17049 8313 17083 8347
rect 17083 8313 17092 8347
rect 17040 8304 17092 8313
rect 17316 8440 17368 8492
rect 18512 8440 18564 8492
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 21272 8508 21324 8560
rect 18604 8440 18656 8449
rect 26976 8576 27028 8628
rect 28356 8576 28408 8628
rect 31668 8576 31720 8628
rect 31852 8576 31904 8628
rect 32128 8619 32180 8628
rect 32128 8585 32137 8619
rect 32137 8585 32171 8619
rect 32171 8585 32180 8619
rect 32128 8576 32180 8585
rect 34152 8576 34204 8628
rect 35900 8619 35952 8628
rect 35900 8585 35909 8619
rect 35909 8585 35943 8619
rect 35943 8585 35952 8619
rect 35900 8576 35952 8585
rect 36268 8619 36320 8628
rect 36268 8585 36277 8619
rect 36277 8585 36311 8619
rect 36311 8585 36320 8619
rect 36268 8576 36320 8585
rect 36636 8619 36688 8628
rect 36636 8585 36645 8619
rect 36645 8585 36679 8619
rect 36679 8585 36688 8619
rect 36636 8576 36688 8585
rect 26516 8508 26568 8560
rect 27068 8440 27120 8492
rect 19156 8372 19208 8424
rect 18420 8304 18472 8356
rect 18696 8304 18748 8356
rect 19064 8304 19116 8356
rect 21364 8372 21416 8424
rect 21548 8372 21600 8424
rect 24216 8372 24268 8424
rect 20536 8304 20588 8356
rect 22560 8347 22612 8356
rect 22560 8313 22569 8347
rect 22569 8313 22603 8347
rect 22603 8313 22612 8347
rect 22560 8304 22612 8313
rect 5540 8236 5592 8288
rect 6092 8236 6144 8288
rect 7380 8236 7432 8288
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 15936 8236 15988 8288
rect 18052 8236 18104 8288
rect 19432 8236 19484 8288
rect 19616 8279 19668 8288
rect 19616 8245 19625 8279
rect 19625 8245 19659 8279
rect 19659 8245 19668 8279
rect 19616 8236 19668 8245
rect 21548 8279 21600 8288
rect 21548 8245 21557 8279
rect 21557 8245 21591 8279
rect 21591 8245 21600 8279
rect 21548 8236 21600 8245
rect 23664 8236 23716 8288
rect 25872 8347 25924 8356
rect 25872 8313 25881 8347
rect 25881 8313 25915 8347
rect 25915 8313 25924 8347
rect 25872 8304 25924 8313
rect 26056 8304 26108 8356
rect 26516 8304 26568 8356
rect 28080 8508 28132 8560
rect 27712 8372 27764 8424
rect 30380 8440 30432 8492
rect 30932 8440 30984 8492
rect 32772 8483 32824 8492
rect 32772 8449 32781 8483
rect 32781 8449 32815 8483
rect 32815 8449 32824 8483
rect 32772 8440 32824 8449
rect 34704 8440 34756 8492
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35256 8440 35308 8449
rect 29000 8372 29052 8424
rect 31576 8415 31628 8424
rect 24676 8236 24728 8288
rect 28908 8304 28960 8356
rect 28080 8236 28132 8288
rect 30196 8347 30248 8356
rect 30196 8313 30205 8347
rect 30205 8313 30239 8347
rect 30239 8313 30248 8347
rect 31576 8381 31620 8415
rect 31620 8381 31628 8415
rect 31576 8372 31628 8381
rect 30196 8304 30248 8313
rect 32680 8347 32732 8356
rect 32680 8313 32689 8347
rect 32689 8313 32723 8347
rect 32723 8313 32732 8347
rect 32680 8304 32732 8313
rect 34152 8304 34204 8356
rect 36084 8372 36136 8424
rect 30656 8236 30708 8288
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 4160 8032 4212 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 5816 8075 5868 8084
rect 5816 8041 5825 8075
rect 5825 8041 5859 8075
rect 5859 8041 5868 8075
rect 5816 8032 5868 8041
rect 6644 8032 6696 8084
rect 8944 8032 8996 8084
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 13728 8032 13780 8084
rect 2320 7964 2372 8016
rect 4436 7964 4488 8016
rect 4804 8007 4856 8016
rect 4804 7973 4813 8007
rect 4813 7973 4847 8007
rect 4847 7973 4856 8007
rect 4804 7964 4856 7973
rect 7196 8007 7248 8016
rect 7196 7973 7199 8007
rect 7199 7973 7233 8007
rect 7233 7973 7248 8007
rect 7196 7964 7248 7973
rect 14740 8032 14792 8084
rect 17040 8032 17092 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 19064 8032 19116 8084
rect 23480 8032 23532 8084
rect 24124 8032 24176 8084
rect 25872 8032 25924 8084
rect 30196 8032 30248 8084
rect 30472 8075 30524 8084
rect 30472 8041 30481 8075
rect 30481 8041 30515 8075
rect 30515 8041 30524 8075
rect 30472 8032 30524 8041
rect 30656 8075 30708 8084
rect 30656 8041 30665 8075
rect 30665 8041 30699 8075
rect 30699 8041 30708 8075
rect 30656 8032 30708 8041
rect 32404 8075 32456 8084
rect 32404 8041 32413 8075
rect 32413 8041 32447 8075
rect 32447 8041 32456 8075
rect 32404 8032 32456 8041
rect 1768 7939 1820 7948
rect 1768 7905 1777 7939
rect 1777 7905 1811 7939
rect 1811 7905 1820 7939
rect 1768 7896 1820 7905
rect 5724 7896 5776 7948
rect 9036 7896 9088 7948
rect 10784 7939 10836 7948
rect 10784 7905 10793 7939
rect 10793 7905 10827 7939
rect 10827 7905 10836 7939
rect 10784 7896 10836 7905
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 11152 7896 11204 7948
rect 12164 7896 12216 7948
rect 14648 8007 14700 8016
rect 14648 7973 14657 8007
rect 14657 7973 14691 8007
rect 14691 7973 14700 8007
rect 14648 7964 14700 7973
rect 15752 7964 15804 8016
rect 4252 7828 4304 7880
rect 6920 7828 6972 7880
rect 9956 7828 10008 7880
rect 12716 7896 12768 7948
rect 13820 7939 13872 7948
rect 13820 7905 13829 7939
rect 13829 7905 13863 7939
rect 13863 7905 13872 7939
rect 13820 7896 13872 7905
rect 14004 7896 14056 7948
rect 17592 7964 17644 8016
rect 19156 7964 19208 8016
rect 22008 7964 22060 8016
rect 24676 7964 24728 8016
rect 26884 8007 26936 8016
rect 26884 7973 26887 8007
rect 26887 7973 26921 8007
rect 26921 7973 26936 8007
rect 26884 7964 26936 7973
rect 29184 7964 29236 8016
rect 34152 7964 34204 8016
rect 35440 8007 35492 8016
rect 35440 7973 35449 8007
rect 35449 7973 35483 8007
rect 35483 7973 35492 8007
rect 35440 7964 35492 7973
rect 35992 8007 36044 8016
rect 35992 7973 36001 8007
rect 36001 7973 36035 8007
rect 36035 7973 36044 8007
rect 35992 7964 36044 7973
rect 18696 7896 18748 7948
rect 22652 7896 22704 7948
rect 23388 7896 23440 7948
rect 29000 7896 29052 7948
rect 30104 7939 30156 7948
rect 30104 7905 30113 7939
rect 30113 7905 30147 7939
rect 30147 7905 30156 7939
rect 30104 7896 30156 7905
rect 30564 7896 30616 7948
rect 32772 7896 32824 7948
rect 35164 7896 35216 7948
rect 14556 7828 14608 7880
rect 17960 7828 18012 7880
rect 18604 7828 18656 7880
rect 18972 7828 19024 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 12624 7760 12676 7812
rect 19064 7760 19116 7812
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 25044 7828 25096 7880
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 28724 7828 28776 7880
rect 33508 7871 33560 7880
rect 33508 7837 33517 7871
rect 33517 7837 33551 7871
rect 33551 7837 33560 7871
rect 33508 7828 33560 7837
rect 35348 7871 35400 7880
rect 35348 7837 35357 7871
rect 35357 7837 35391 7871
rect 35391 7837 35400 7871
rect 35348 7828 35400 7837
rect 22100 7760 22152 7769
rect 24860 7760 24912 7812
rect 31024 7760 31076 7812
rect 33600 7760 33652 7812
rect 3516 7692 3568 7744
rect 9772 7692 9824 7744
rect 13636 7692 13688 7744
rect 14004 7692 14056 7744
rect 16948 7692 17000 7744
rect 18420 7692 18472 7744
rect 19248 7692 19300 7744
rect 20812 7692 20864 7744
rect 22560 7692 22612 7744
rect 23296 7692 23348 7744
rect 24216 7735 24268 7744
rect 24216 7701 24225 7735
rect 24225 7701 24259 7735
rect 24259 7701 24268 7735
rect 24216 7692 24268 7701
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 27712 7735 27764 7744
rect 27712 7701 27721 7735
rect 27721 7701 27755 7735
rect 27755 7701 27764 7735
rect 27712 7692 27764 7701
rect 33140 7692 33192 7744
rect 34888 7735 34940 7744
rect 34888 7701 34897 7735
rect 34897 7701 34931 7735
rect 34931 7701 34940 7735
rect 34888 7692 34940 7701
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 8760 7531 8812 7540
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 10232 7488 10284 7540
rect 10784 7488 10836 7540
rect 12624 7488 12676 7540
rect 13728 7488 13780 7540
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 15292 7531 15344 7540
rect 15292 7497 15301 7531
rect 15301 7497 15335 7531
rect 15335 7497 15344 7531
rect 15292 7488 15344 7497
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 9956 7463 10008 7472
rect 9956 7429 9965 7463
rect 9965 7429 9999 7463
rect 9999 7429 10008 7463
rect 9956 7420 10008 7429
rect 12164 7463 12216 7472
rect 12164 7429 12173 7463
rect 12173 7429 12207 7463
rect 12207 7429 12216 7463
rect 12164 7420 12216 7429
rect 13544 7420 13596 7472
rect 18788 7420 18840 7472
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 9036 7352 9088 7404
rect 10968 7352 11020 7404
rect 13820 7352 13872 7404
rect 17040 7352 17092 7404
rect 20628 7488 20680 7540
rect 22008 7488 22060 7540
rect 26884 7488 26936 7540
rect 31024 7531 31076 7540
rect 31024 7497 31033 7531
rect 31033 7497 31067 7531
rect 31067 7497 31076 7531
rect 31024 7488 31076 7497
rect 32772 7531 32824 7540
rect 32772 7497 32781 7531
rect 32781 7497 32815 7531
rect 32815 7497 32824 7531
rect 32772 7488 32824 7497
rect 34152 7488 34204 7540
rect 35440 7488 35492 7540
rect 36636 7531 36688 7540
rect 36636 7497 36645 7531
rect 36645 7497 36679 7531
rect 36679 7497 36688 7531
rect 36636 7488 36688 7497
rect 19524 7420 19576 7472
rect 34888 7420 34940 7472
rect 19156 7352 19208 7404
rect 21548 7352 21600 7404
rect 24216 7395 24268 7404
rect 24216 7361 24225 7395
rect 24225 7361 24259 7395
rect 24259 7361 24268 7395
rect 24216 7352 24268 7361
rect 26148 7352 26200 7404
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 27988 7352 28040 7404
rect 28080 7395 28132 7404
rect 28080 7361 28089 7395
rect 28089 7361 28123 7395
rect 28123 7361 28132 7395
rect 30104 7395 30156 7404
rect 28080 7352 28132 7361
rect 30104 7361 30113 7395
rect 30113 7361 30147 7395
rect 30147 7361 30156 7395
rect 30104 7352 30156 7361
rect 3516 7284 3568 7336
rect 6736 7284 6788 7336
rect 8024 7284 8076 7336
rect 12624 7327 12676 7336
rect 12624 7293 12642 7327
rect 12642 7293 12676 7327
rect 12624 7284 12676 7293
rect 2320 7148 2372 7200
rect 3608 7148 3660 7200
rect 5540 7216 5592 7268
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 6920 7148 6972 7200
rect 7104 7148 7156 7200
rect 7196 7148 7248 7200
rect 10232 7259 10284 7268
rect 10232 7225 10241 7259
rect 10241 7225 10275 7259
rect 10275 7225 10284 7259
rect 10232 7216 10284 7225
rect 13636 7259 13688 7268
rect 13636 7225 13645 7259
rect 13645 7225 13679 7259
rect 13679 7225 13688 7259
rect 13636 7216 13688 7225
rect 13728 7259 13780 7268
rect 13728 7225 13737 7259
rect 13737 7225 13771 7259
rect 13771 7225 13780 7259
rect 13728 7216 13780 7225
rect 15752 7216 15804 7268
rect 16580 7259 16632 7268
rect 16580 7225 16583 7259
rect 16583 7225 16617 7259
rect 16617 7225 16632 7259
rect 16580 7216 16632 7225
rect 10600 7148 10652 7200
rect 12808 7148 12860 7200
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 20168 7327 20220 7336
rect 20168 7293 20212 7327
rect 20212 7293 20220 7327
rect 20168 7284 20220 7293
rect 22192 7284 22244 7336
rect 23388 7284 23440 7336
rect 23940 7327 23992 7336
rect 23940 7293 23949 7327
rect 23949 7293 23983 7327
rect 23983 7293 23992 7327
rect 23940 7284 23992 7293
rect 24124 7327 24176 7336
rect 24124 7293 24133 7327
rect 24133 7293 24167 7327
rect 24167 7293 24176 7327
rect 24124 7284 24176 7293
rect 21364 7259 21416 7268
rect 18604 7148 18656 7200
rect 21364 7225 21373 7259
rect 21373 7225 21407 7259
rect 21407 7225 21416 7259
rect 21364 7216 21416 7225
rect 26884 7216 26936 7268
rect 19248 7148 19300 7200
rect 22652 7191 22704 7200
rect 22652 7157 22661 7191
rect 22661 7157 22695 7191
rect 22695 7157 22704 7191
rect 22652 7148 22704 7157
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 25044 7191 25096 7200
rect 25044 7157 25053 7191
rect 25053 7157 25087 7191
rect 25087 7157 25096 7191
rect 25044 7148 25096 7157
rect 28724 7216 28776 7268
rect 32680 7352 32732 7404
rect 33140 7352 33192 7404
rect 35348 7395 35400 7404
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 32036 7284 32088 7336
rect 34428 7284 34480 7336
rect 36452 7327 36504 7336
rect 36452 7293 36461 7327
rect 36461 7293 36495 7327
rect 36495 7293 36504 7327
rect 36452 7284 36504 7293
rect 33600 7216 33652 7268
rect 33232 7148 33284 7200
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 1768 6987 1820 6996
rect 1768 6953 1777 6987
rect 1777 6953 1811 6987
rect 1811 6953 1820 6987
rect 1768 6944 1820 6953
rect 10600 6987 10652 6996
rect 10600 6953 10609 6987
rect 10609 6953 10643 6987
rect 10643 6953 10652 6987
rect 10600 6944 10652 6953
rect 14004 6944 14056 6996
rect 17960 6944 18012 6996
rect 22008 6987 22060 6996
rect 22008 6953 22017 6987
rect 22017 6953 22051 6987
rect 22051 6953 22060 6987
rect 22008 6944 22060 6953
rect 26148 6944 26200 6996
rect 33140 6944 33192 6996
rect 2320 6876 2372 6928
rect 3608 6876 3660 6928
rect 4160 6808 4212 6860
rect 4436 6876 4488 6928
rect 5080 6876 5132 6928
rect 6644 6808 6696 6860
rect 7196 6876 7248 6928
rect 9772 6876 9824 6928
rect 8668 6808 8720 6860
rect 12072 6808 12124 6860
rect 16304 6876 16356 6928
rect 15016 6808 15068 6860
rect 16672 6851 16724 6860
rect 16672 6817 16681 6851
rect 16681 6817 16715 6851
rect 16715 6817 16724 6851
rect 16672 6808 16724 6817
rect 17776 6851 17828 6860
rect 2596 6740 2648 6792
rect 4068 6740 4120 6792
rect 5264 6740 5316 6792
rect 6828 6740 6880 6792
rect 10232 6740 10284 6792
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 14832 6740 14884 6792
rect 16856 6740 16908 6792
rect 3332 6672 3384 6724
rect 8760 6715 8812 6724
rect 8760 6681 8769 6715
rect 8769 6681 8803 6715
rect 8803 6681 8812 6715
rect 8760 6672 8812 6681
rect 14188 6672 14240 6724
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 19156 6808 19208 6860
rect 19248 6808 19300 6860
rect 19616 6808 19668 6860
rect 20812 6808 20864 6860
rect 18144 6783 18196 6792
rect 18144 6749 18153 6783
rect 18153 6749 18187 6783
rect 18187 6749 18196 6783
rect 18144 6740 18196 6749
rect 20720 6783 20772 6792
rect 18420 6672 18472 6724
rect 20720 6749 20729 6783
rect 20729 6749 20763 6783
rect 20763 6749 20772 6783
rect 20720 6740 20772 6749
rect 21640 6783 21692 6792
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 22100 6740 22152 6792
rect 21272 6672 21324 6724
rect 21824 6672 21876 6724
rect 23940 6876 23992 6928
rect 25044 6876 25096 6928
rect 27436 6876 27488 6928
rect 28080 6876 28132 6928
rect 28816 6919 28868 6928
rect 28816 6885 28825 6919
rect 28825 6885 28859 6919
rect 28859 6885 28868 6919
rect 28816 6876 28868 6885
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 24860 6808 24912 6860
rect 25320 6851 25372 6860
rect 25320 6817 25329 6851
rect 25329 6817 25363 6851
rect 25363 6817 25372 6851
rect 25320 6808 25372 6817
rect 30380 6851 30432 6860
rect 30380 6817 30389 6851
rect 30389 6817 30423 6851
rect 30423 6817 30432 6851
rect 30380 6808 30432 6817
rect 30564 6808 30616 6860
rect 32680 6876 32732 6928
rect 34612 6919 34664 6928
rect 34612 6885 34621 6919
rect 34621 6885 34655 6919
rect 34655 6885 34664 6919
rect 34612 6876 34664 6885
rect 35348 6944 35400 6996
rect 36176 6919 36228 6928
rect 36176 6885 36185 6919
rect 36185 6885 36219 6919
rect 36219 6885 36228 6919
rect 36176 6876 36228 6885
rect 26332 6740 26384 6792
rect 28908 6740 28960 6792
rect 29092 6783 29144 6792
rect 29092 6749 29101 6783
rect 29101 6749 29135 6783
rect 29135 6749 29144 6783
rect 29092 6740 29144 6749
rect 31576 6808 31628 6860
rect 31116 6740 31168 6792
rect 33876 6740 33928 6792
rect 34152 6740 34204 6792
rect 36084 6783 36136 6792
rect 36084 6749 36093 6783
rect 36093 6749 36127 6783
rect 36127 6749 36136 6783
rect 36084 6740 36136 6749
rect 36360 6783 36412 6792
rect 36360 6749 36369 6783
rect 36369 6749 36403 6783
rect 36403 6749 36412 6783
rect 36360 6740 36412 6749
rect 24952 6672 25004 6724
rect 26056 6672 26108 6724
rect 2780 6604 2832 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 7012 6604 7064 6656
rect 8024 6604 8076 6656
rect 8484 6604 8536 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 12900 6647 12952 6656
rect 12900 6613 12909 6647
rect 12909 6613 12943 6647
rect 12943 6613 12952 6647
rect 12900 6604 12952 6613
rect 14004 6647 14056 6656
rect 14004 6613 14013 6647
rect 14013 6613 14047 6647
rect 14047 6613 14056 6647
rect 14004 6604 14056 6613
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18972 6604 19024 6656
rect 21548 6604 21600 6656
rect 23388 6604 23440 6656
rect 26240 6604 26292 6656
rect 26516 6604 26568 6656
rect 33048 6647 33100 6656
rect 33048 6613 33057 6647
rect 33057 6613 33091 6647
rect 33091 6613 33100 6647
rect 33048 6604 33100 6613
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2228 6400 2280 6452
rect 4160 6443 4212 6452
rect 4160 6409 4169 6443
rect 4169 6409 4203 6443
rect 4203 6409 4212 6443
rect 4160 6400 4212 6409
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 5540 6400 5592 6452
rect 6644 6400 6696 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 12072 6443 12124 6452
rect 12072 6409 12081 6443
rect 12081 6409 12115 6443
rect 12115 6409 12124 6443
rect 12072 6400 12124 6409
rect 13728 6400 13780 6452
rect 14004 6400 14056 6452
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 16580 6443 16632 6452
rect 16580 6409 16589 6443
rect 16589 6409 16623 6443
rect 16623 6409 16632 6443
rect 16580 6400 16632 6409
rect 16856 6400 16908 6452
rect 17776 6400 17828 6452
rect 20812 6400 20864 6452
rect 21824 6443 21876 6452
rect 21824 6409 21833 6443
rect 21833 6409 21867 6443
rect 21867 6409 21876 6443
rect 21824 6400 21876 6409
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 24032 6400 24084 6452
rect 24952 6443 25004 6452
rect 24952 6409 24961 6443
rect 24961 6409 24995 6443
rect 24995 6409 25004 6443
rect 24952 6400 25004 6409
rect 25320 6443 25372 6452
rect 25320 6409 25329 6443
rect 25329 6409 25363 6443
rect 25363 6409 25372 6443
rect 25320 6400 25372 6409
rect 27436 6400 27488 6452
rect 28816 6400 28868 6452
rect 30564 6443 30616 6452
rect 30564 6409 30573 6443
rect 30573 6409 30607 6443
rect 30607 6409 30616 6443
rect 30564 6400 30616 6409
rect 32680 6400 32732 6452
rect 33876 6443 33928 6452
rect 33876 6409 33885 6443
rect 33885 6409 33919 6443
rect 33919 6409 33928 6443
rect 33876 6400 33928 6409
rect 36084 6400 36136 6452
rect 36452 6400 36504 6452
rect 3332 6375 3384 6384
rect 3332 6341 3341 6375
rect 3341 6341 3375 6375
rect 3375 6341 3384 6375
rect 3332 6332 3384 6341
rect 24584 6375 24636 6384
rect 24584 6341 24593 6375
rect 24593 6341 24627 6375
rect 24627 6341 24636 6375
rect 24584 6332 24636 6341
rect 2504 6264 2556 6316
rect 3424 6264 3476 6316
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 4620 6307 4672 6316
rect 4620 6273 4629 6307
rect 4629 6273 4663 6307
rect 4663 6273 4672 6307
rect 4620 6264 4672 6273
rect 7012 6264 7064 6316
rect 9036 6264 9088 6316
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 18696 6264 18748 6316
rect 28080 6332 28132 6384
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 29092 6264 29144 6316
rect 31116 6264 31168 6316
rect 33048 6332 33100 6384
rect 34612 6332 34664 6384
rect 36176 6332 36228 6384
rect 35348 6307 35400 6316
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 1676 6128 1728 6180
rect 2320 6171 2372 6180
rect 2320 6137 2329 6171
rect 2329 6137 2363 6171
rect 2363 6137 2372 6171
rect 2320 6128 2372 6137
rect 3148 6128 3200 6180
rect 2780 6060 2832 6112
rect 4620 6128 4672 6180
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 8300 6128 8352 6180
rect 12992 6196 13044 6248
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 15384 6239 15436 6248
rect 15384 6205 15393 6239
rect 15393 6205 15427 6239
rect 15427 6205 15436 6239
rect 15384 6196 15436 6205
rect 20168 6196 20220 6248
rect 21824 6196 21876 6248
rect 22560 6239 22612 6248
rect 22560 6205 22569 6239
rect 22569 6205 22603 6239
rect 22603 6205 22612 6239
rect 22560 6196 22612 6205
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 25872 6239 25924 6248
rect 25872 6205 25881 6239
rect 25881 6205 25915 6239
rect 25915 6205 25924 6239
rect 25872 6196 25924 6205
rect 31392 6239 31444 6248
rect 31392 6205 31401 6239
rect 31401 6205 31435 6239
rect 31435 6205 31444 6239
rect 31392 6196 31444 6205
rect 32680 6239 32732 6248
rect 32680 6205 32689 6239
rect 32689 6205 32723 6239
rect 32723 6205 32732 6239
rect 32680 6196 32732 6205
rect 10784 6171 10836 6180
rect 10784 6137 10793 6171
rect 10793 6137 10827 6171
rect 10827 6137 10836 6171
rect 10784 6128 10836 6137
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 12072 6128 12124 6180
rect 13176 6128 13228 6180
rect 15752 6171 15804 6180
rect 15752 6137 15755 6171
rect 15755 6137 15789 6171
rect 15789 6137 15804 6171
rect 15752 6128 15804 6137
rect 18604 6171 18656 6180
rect 18604 6137 18613 6171
rect 18613 6137 18647 6171
rect 18647 6137 18656 6171
rect 18604 6128 18656 6137
rect 19616 6128 19668 6180
rect 21364 6128 21416 6180
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 10232 6060 10284 6112
rect 14188 6060 14240 6112
rect 15016 6060 15068 6112
rect 18420 6060 18472 6112
rect 20720 6060 20772 6112
rect 22284 6103 22336 6112
rect 22284 6069 22293 6103
rect 22293 6069 22327 6103
rect 22327 6069 22336 6103
rect 22284 6060 22336 6069
rect 23388 6103 23440 6112
rect 23388 6069 23397 6103
rect 23397 6069 23431 6103
rect 23431 6069 23440 6103
rect 23388 6060 23440 6069
rect 24676 6060 24728 6112
rect 28816 6128 28868 6180
rect 29368 6171 29420 6180
rect 29368 6137 29377 6171
rect 29377 6137 29411 6171
rect 29411 6137 29420 6171
rect 29368 6128 29420 6137
rect 35348 6273 35357 6307
rect 35357 6273 35391 6307
rect 35391 6273 35400 6307
rect 35348 6264 35400 6273
rect 34612 6239 34664 6248
rect 34612 6205 34621 6239
rect 34621 6205 34655 6239
rect 34655 6205 34664 6239
rect 34612 6196 34664 6205
rect 35900 6196 35952 6248
rect 34980 6171 35032 6180
rect 29184 6060 29236 6112
rect 34980 6137 34989 6171
rect 34989 6137 35023 6171
rect 35023 6137 35032 6171
rect 34980 6128 35032 6137
rect 34612 6060 34664 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 3148 5856 3200 5908
rect 4344 5856 4396 5908
rect 6828 5856 6880 5908
rect 6920 5856 6972 5908
rect 8668 5856 8720 5908
rect 9128 5856 9180 5908
rect 9588 5856 9640 5908
rect 11980 5899 12032 5908
rect 2044 5831 2096 5840
rect 2044 5797 2053 5831
rect 2053 5797 2087 5831
rect 2087 5797 2096 5831
rect 2044 5788 2096 5797
rect 5816 5831 5868 5840
rect 5816 5797 5825 5831
rect 5825 5797 5859 5831
rect 5859 5797 5868 5831
rect 5816 5788 5868 5797
rect 7104 5831 7156 5840
rect 7104 5797 7113 5831
rect 7113 5797 7147 5831
rect 7147 5797 7156 5831
rect 7104 5788 7156 5797
rect 9496 5788 9548 5840
rect 9772 5788 9824 5840
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 12348 5856 12400 5908
rect 13176 5899 13228 5908
rect 13176 5865 13185 5899
rect 13185 5865 13219 5899
rect 13219 5865 13228 5899
rect 13176 5856 13228 5865
rect 13912 5856 13964 5908
rect 16672 5856 16724 5908
rect 17776 5856 17828 5908
rect 18604 5856 18656 5908
rect 19892 5899 19944 5908
rect 19892 5865 19901 5899
rect 19901 5865 19935 5899
rect 19935 5865 19944 5899
rect 19892 5856 19944 5865
rect 22560 5856 22612 5908
rect 23664 5856 23716 5908
rect 26332 5899 26384 5908
rect 26332 5865 26341 5899
rect 26341 5865 26375 5899
rect 26375 5865 26384 5899
rect 26332 5856 26384 5865
rect 31116 5899 31168 5908
rect 31116 5865 31125 5899
rect 31125 5865 31159 5899
rect 31159 5865 31168 5899
rect 31116 5856 31168 5865
rect 32680 5899 32732 5908
rect 32680 5865 32689 5899
rect 32689 5865 32723 5899
rect 32723 5865 32732 5899
rect 32680 5856 32732 5865
rect 34152 5856 34204 5908
rect 34980 5856 35032 5908
rect 36452 5899 36504 5908
rect 36452 5865 36461 5899
rect 36461 5865 36495 5899
rect 36495 5865 36504 5899
rect 36452 5856 36504 5865
rect 12164 5788 12216 5840
rect 12808 5788 12860 5840
rect 13452 5788 13504 5840
rect 14096 5788 14148 5840
rect 16396 5788 16448 5840
rect 16948 5831 17000 5840
rect 16948 5797 16957 5831
rect 16957 5797 16991 5831
rect 16991 5797 17000 5831
rect 16948 5788 17000 5797
rect 4160 5695 4212 5704
rect 4160 5661 4169 5695
rect 4169 5661 4203 5695
rect 4203 5661 4212 5695
rect 4160 5652 4212 5661
rect 4620 5652 4672 5704
rect 5540 5652 5592 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6828 5652 6880 5704
rect 8300 5720 8352 5772
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 11888 5652 11940 5704
rect 14924 5652 14976 5704
rect 15200 5652 15252 5704
rect 10876 5627 10928 5636
rect 10876 5593 10885 5627
rect 10885 5593 10919 5627
rect 10919 5593 10928 5627
rect 10876 5584 10928 5593
rect 13728 5584 13780 5636
rect 16764 5652 16816 5704
rect 19616 5788 19668 5840
rect 20720 5788 20772 5840
rect 21640 5831 21692 5840
rect 21640 5797 21649 5831
rect 21649 5797 21683 5831
rect 21683 5797 21692 5831
rect 21640 5788 21692 5797
rect 23388 5788 23440 5840
rect 27160 5831 27212 5840
rect 27160 5797 27169 5831
rect 27169 5797 27203 5831
rect 27203 5797 27212 5831
rect 27160 5788 27212 5797
rect 27988 5788 28040 5840
rect 28632 5788 28684 5840
rect 30840 5831 30892 5840
rect 30840 5797 30849 5831
rect 30849 5797 30883 5831
rect 30883 5797 30892 5831
rect 30840 5788 30892 5797
rect 18328 5720 18380 5772
rect 19248 5720 19300 5772
rect 24860 5720 24912 5772
rect 25136 5763 25188 5772
rect 25136 5729 25145 5763
rect 25145 5729 25179 5763
rect 25179 5729 25188 5763
rect 25136 5720 25188 5729
rect 29276 5720 29328 5772
rect 30104 5763 30156 5772
rect 30104 5729 30113 5763
rect 30113 5729 30147 5763
rect 30147 5729 30156 5763
rect 30104 5720 30156 5729
rect 30380 5720 30432 5772
rect 34612 5831 34664 5840
rect 34612 5797 34621 5831
rect 34621 5797 34655 5831
rect 34655 5797 34664 5831
rect 34612 5788 34664 5797
rect 34704 5788 34756 5840
rect 36360 5788 36412 5840
rect 32220 5763 32272 5772
rect 32220 5729 32238 5763
rect 32238 5729 32272 5763
rect 32220 5720 32272 5729
rect 33416 5763 33468 5772
rect 33416 5729 33460 5763
rect 33460 5729 33468 5763
rect 33416 5720 33468 5729
rect 35992 5763 36044 5772
rect 35992 5729 36036 5763
rect 36036 5729 36044 5763
rect 35992 5720 36044 5729
rect 20812 5652 20864 5704
rect 22284 5652 22336 5704
rect 25504 5695 25556 5704
rect 25504 5661 25513 5695
rect 25513 5661 25547 5695
rect 25547 5661 25556 5695
rect 25504 5652 25556 5661
rect 27068 5695 27120 5704
rect 27068 5661 27077 5695
rect 27077 5661 27111 5695
rect 27111 5661 27120 5695
rect 27068 5652 27120 5661
rect 28908 5652 28960 5704
rect 29092 5695 29144 5704
rect 29092 5661 29101 5695
rect 29101 5661 29135 5695
rect 29135 5661 29144 5695
rect 29092 5652 29144 5661
rect 34152 5652 34204 5704
rect 24124 5627 24176 5636
rect 24124 5593 24133 5627
rect 24133 5593 24167 5627
rect 24167 5593 24176 5627
rect 24124 5584 24176 5593
rect 29368 5584 29420 5636
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 2596 5516 2648 5568
rect 4344 5516 4396 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 15384 5516 15436 5568
rect 16488 5516 16540 5568
rect 18144 5516 18196 5568
rect 19340 5516 19392 5568
rect 20168 5559 20220 5568
rect 20168 5525 20177 5559
rect 20177 5525 20211 5559
rect 20211 5525 20220 5559
rect 20168 5516 20220 5525
rect 21732 5516 21784 5568
rect 25872 5559 25924 5568
rect 25872 5525 25881 5559
rect 25881 5525 25915 5559
rect 25915 5525 25924 5559
rect 25872 5516 25924 5525
rect 28080 5559 28132 5568
rect 28080 5525 28089 5559
rect 28089 5525 28123 5559
rect 28123 5525 28132 5559
rect 28080 5516 28132 5525
rect 29092 5516 29144 5568
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 2044 5312 2096 5364
rect 5816 5312 5868 5364
rect 5908 5355 5960 5364
rect 5908 5321 5917 5355
rect 5917 5321 5951 5355
rect 5951 5321 5960 5355
rect 6644 5355 6696 5364
rect 5908 5312 5960 5321
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 6828 5312 6880 5364
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 9128 5355 9180 5364
rect 9128 5321 9137 5355
rect 9137 5321 9171 5355
rect 9171 5321 9180 5355
rect 9128 5312 9180 5321
rect 9772 5312 9824 5364
rect 12164 5355 12216 5364
rect 7196 5244 7248 5296
rect 1768 5108 1820 5160
rect 3700 5151 3752 5160
rect 3700 5117 3709 5151
rect 3709 5117 3743 5151
rect 3743 5117 3752 5151
rect 3700 5108 3752 5117
rect 1676 5040 1728 5092
rect 4160 5108 4212 5160
rect 6368 5108 6420 5160
rect 3240 5015 3292 5024
rect 3240 4981 3249 5015
rect 3249 4981 3283 5015
rect 3283 4981 3292 5015
rect 3240 4972 3292 4981
rect 3608 5015 3660 5024
rect 3608 4981 3617 5015
rect 3617 4981 3651 5015
rect 3651 4981 3660 5015
rect 6828 5040 6880 5092
rect 12164 5321 12173 5355
rect 12173 5321 12207 5355
rect 12207 5321 12216 5355
rect 12164 5312 12216 5321
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 17776 5312 17828 5364
rect 19616 5312 19668 5364
rect 20536 5355 20588 5364
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 20812 5312 20864 5364
rect 22284 5312 22336 5364
rect 23480 5312 23532 5364
rect 24768 5355 24820 5364
rect 24768 5321 24777 5355
rect 24777 5321 24811 5355
rect 24811 5321 24820 5355
rect 24768 5312 24820 5321
rect 25228 5312 25280 5364
rect 26056 5312 26108 5364
rect 26884 5355 26936 5364
rect 26884 5321 26893 5355
rect 26893 5321 26927 5355
rect 26927 5321 26936 5355
rect 26884 5312 26936 5321
rect 27252 5312 27304 5364
rect 29000 5312 29052 5364
rect 29736 5355 29788 5364
rect 29736 5321 29745 5355
rect 29745 5321 29779 5355
rect 29779 5321 29788 5355
rect 29736 5312 29788 5321
rect 30104 5355 30156 5364
rect 30104 5321 30113 5355
rect 30113 5321 30147 5355
rect 30147 5321 30156 5355
rect 30104 5312 30156 5321
rect 30380 5312 30432 5364
rect 32220 5355 32272 5364
rect 32220 5321 32229 5355
rect 32229 5321 32263 5355
rect 32263 5321 32272 5355
rect 32220 5312 32272 5321
rect 33416 5355 33468 5364
rect 33416 5321 33425 5355
rect 33425 5321 33459 5355
rect 33459 5321 33468 5355
rect 33416 5312 33468 5321
rect 34152 5355 34204 5364
rect 34152 5321 34161 5355
rect 34161 5321 34195 5355
rect 34195 5321 34204 5355
rect 34152 5312 34204 5321
rect 34612 5312 34664 5364
rect 34980 5312 35032 5364
rect 13728 5287 13780 5296
rect 13728 5253 13737 5287
rect 13737 5253 13771 5287
rect 13771 5253 13780 5287
rect 13728 5244 13780 5253
rect 32772 5244 32824 5296
rect 8208 5151 8260 5160
rect 8208 5117 8217 5151
rect 8217 5117 8251 5151
rect 8251 5117 8260 5151
rect 8208 5108 8260 5117
rect 9772 5040 9824 5092
rect 13820 5176 13872 5228
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 14924 5176 14976 5228
rect 16396 5176 16448 5228
rect 16580 5176 16632 5228
rect 20168 5219 20220 5228
rect 20168 5185 20177 5219
rect 20177 5185 20211 5219
rect 20211 5185 20220 5219
rect 20168 5176 20220 5185
rect 25872 5219 25924 5228
rect 25872 5185 25881 5219
rect 25881 5185 25915 5219
rect 25915 5185 25924 5219
rect 25872 5176 25924 5185
rect 27988 5176 28040 5228
rect 28908 5176 28960 5228
rect 16212 5151 16264 5160
rect 16212 5117 16221 5151
rect 16221 5117 16255 5151
rect 16255 5117 16264 5151
rect 16212 5108 16264 5117
rect 13176 5083 13228 5092
rect 13176 5049 13185 5083
rect 13185 5049 13219 5083
rect 13219 5049 13228 5083
rect 13176 5040 13228 5049
rect 14832 5083 14884 5092
rect 10048 5015 10100 5024
rect 3608 4972 3660 4981
rect 10048 4981 10057 5015
rect 10057 4981 10091 5015
rect 10091 4981 10100 5015
rect 10048 4972 10100 4981
rect 14832 5049 14841 5083
rect 14841 5049 14875 5083
rect 14875 5049 14884 5083
rect 14832 5040 14884 5049
rect 15108 5040 15160 5092
rect 17132 5108 17184 5160
rect 13728 4972 13780 5024
rect 15568 4972 15620 5024
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 19800 5108 19852 5160
rect 19064 5040 19116 5092
rect 20536 5108 20588 5160
rect 21732 5151 21784 5160
rect 21732 5117 21741 5151
rect 21741 5117 21775 5151
rect 21775 5117 21784 5151
rect 21732 5108 21784 5117
rect 23296 5108 23348 5160
rect 25228 5151 25280 5160
rect 20628 5040 20680 5092
rect 22560 5040 22612 5092
rect 24032 5040 24084 5092
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 25320 5040 25372 5092
rect 26056 5108 26108 5160
rect 29736 5108 29788 5160
rect 31300 5151 31352 5160
rect 31300 5117 31344 5151
rect 31344 5117 31352 5151
rect 31300 5108 31352 5117
rect 17776 4972 17828 4981
rect 19156 4972 19208 5024
rect 23388 4972 23440 5024
rect 23664 4972 23716 5024
rect 27252 5083 27304 5092
rect 27252 5049 27261 5083
rect 27261 5049 27295 5083
rect 27295 5049 27304 5083
rect 27252 5040 27304 5049
rect 28172 5015 28224 5024
rect 28172 4981 28181 5015
rect 28181 4981 28215 5015
rect 28215 4981 28224 5015
rect 28172 4972 28224 4981
rect 28540 5015 28592 5024
rect 28540 4981 28549 5015
rect 28549 4981 28583 5015
rect 28583 4981 28592 5015
rect 28540 4972 28592 4981
rect 31760 5015 31812 5024
rect 31760 4981 31769 5015
rect 31769 4981 31803 5015
rect 31803 4981 31812 5015
rect 35440 5015 35492 5024
rect 31760 4972 31812 4981
rect 35440 4981 35449 5015
rect 35449 4981 35483 5015
rect 35483 4981 35492 5015
rect 35440 4972 35492 4981
rect 35992 5015 36044 5024
rect 35992 4981 36001 5015
rect 36001 4981 36035 5015
rect 36035 4981 36044 5015
rect 35992 4972 36044 4981
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2044 4768 2096 4820
rect 3700 4768 3752 4820
rect 6736 4768 6788 4820
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 12440 4768 12492 4820
rect 13452 4811 13504 4820
rect 13452 4777 13461 4811
rect 13461 4777 13495 4811
rect 13495 4777 13504 4811
rect 13452 4768 13504 4777
rect 14832 4768 14884 4820
rect 17040 4768 17092 4820
rect 2688 4700 2740 4752
rect 6368 4743 6420 4752
rect 6368 4709 6377 4743
rect 6377 4709 6411 4743
rect 6411 4709 6420 4743
rect 6368 4700 6420 4709
rect 8208 4700 8260 4752
rect 9772 4700 9824 4752
rect 13820 4743 13872 4752
rect 13820 4709 13829 4743
rect 13829 4709 13863 4743
rect 13863 4709 13872 4743
rect 13820 4700 13872 4709
rect 14924 4700 14976 4752
rect 1676 4632 1728 4684
rect 4528 4675 4580 4684
rect 2688 4564 2740 4616
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 4528 4641 4537 4675
rect 4537 4641 4571 4675
rect 4571 4641 4580 4675
rect 4528 4632 4580 4641
rect 5540 4675 5592 4684
rect 5540 4641 5549 4675
rect 5549 4641 5583 4675
rect 5583 4641 5592 4675
rect 5540 4632 5592 4641
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5908 4675 5960 4684
rect 5632 4632 5684 4641
rect 5908 4641 5921 4675
rect 5921 4641 5960 4675
rect 5908 4632 5960 4641
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 7472 4675 7524 4684
rect 7472 4641 7481 4675
rect 7481 4641 7515 4675
rect 7515 4641 7524 4675
rect 7472 4632 7524 4641
rect 4436 4564 4488 4616
rect 9864 4632 9916 4684
rect 10968 4632 11020 4684
rect 12256 4675 12308 4684
rect 12256 4641 12265 4675
rect 12265 4641 12299 4675
rect 12299 4641 12308 4675
rect 12256 4632 12308 4641
rect 12624 4675 12676 4684
rect 12624 4641 12633 4675
rect 12633 4641 12667 4675
rect 12667 4641 12676 4675
rect 12624 4632 12676 4641
rect 15292 4675 15344 4684
rect 15292 4641 15301 4675
rect 15301 4641 15335 4675
rect 15335 4641 15344 4675
rect 15292 4632 15344 4641
rect 16396 4700 16448 4752
rect 16672 4743 16724 4752
rect 16672 4709 16681 4743
rect 16681 4709 16715 4743
rect 16715 4709 16724 4743
rect 16672 4700 16724 4709
rect 17500 4700 17552 4752
rect 15844 4675 15896 4684
rect 15844 4641 15853 4675
rect 15853 4641 15887 4675
rect 15887 4641 15896 4675
rect 15844 4632 15896 4641
rect 16304 4632 16356 4684
rect 10140 4607 10192 4616
rect 4896 4496 4948 4548
rect 5264 4496 5316 4548
rect 7104 4496 7156 4548
rect 8484 4496 8536 4548
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 18696 4632 18748 4684
rect 19248 4768 19300 4820
rect 19984 4811 20036 4820
rect 19984 4777 19993 4811
rect 19993 4777 20027 4811
rect 20027 4777 20036 4811
rect 19984 4768 20036 4777
rect 20720 4811 20772 4820
rect 20720 4777 20729 4811
rect 20729 4777 20763 4811
rect 20763 4777 20772 4811
rect 20720 4768 20772 4777
rect 20812 4768 20864 4820
rect 23296 4768 23348 4820
rect 25136 4768 25188 4820
rect 27160 4768 27212 4820
rect 28540 4768 28592 4820
rect 29092 4768 29144 4820
rect 18972 4743 19024 4752
rect 18972 4709 18981 4743
rect 18981 4709 19015 4743
rect 19015 4709 19024 4743
rect 18972 4700 19024 4709
rect 26148 4700 26200 4752
rect 28724 4700 28776 4752
rect 30288 4768 30340 4820
rect 19064 4632 19116 4684
rect 19340 4632 19392 4684
rect 22744 4632 22796 4684
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 22928 4632 22980 4641
rect 25320 4675 25372 4684
rect 1952 4428 2004 4480
rect 8392 4471 8444 4480
rect 8392 4437 8401 4471
rect 8401 4437 8435 4471
rect 8435 4437 8444 4471
rect 8392 4428 8444 4437
rect 9588 4428 9640 4480
rect 9956 4496 10008 4548
rect 17132 4607 17184 4616
rect 17132 4573 17141 4607
rect 17141 4573 17175 4607
rect 17175 4573 17184 4607
rect 17132 4564 17184 4573
rect 25320 4641 25329 4675
rect 25329 4641 25363 4675
rect 25363 4641 25372 4675
rect 25320 4632 25372 4641
rect 27160 4675 27212 4684
rect 27160 4641 27169 4675
rect 27169 4641 27203 4675
rect 27203 4641 27212 4675
rect 27160 4632 27212 4641
rect 28080 4675 28132 4684
rect 28080 4641 28089 4675
rect 28089 4641 28123 4675
rect 28123 4641 28132 4675
rect 28080 4632 28132 4641
rect 28264 4632 28316 4684
rect 30196 4632 30248 4684
rect 25780 4564 25832 4616
rect 26516 4607 26568 4616
rect 26516 4573 26525 4607
rect 26525 4573 26559 4607
rect 26559 4573 26568 4607
rect 26516 4564 26568 4573
rect 10876 4428 10928 4480
rect 11888 4471 11940 4480
rect 11888 4437 11897 4471
rect 11897 4437 11931 4471
rect 11931 4437 11940 4471
rect 11888 4428 11940 4437
rect 12440 4428 12492 4480
rect 13176 4428 13228 4480
rect 16672 4428 16724 4480
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 18052 4428 18104 4480
rect 19892 4428 19944 4480
rect 22284 4428 22336 4480
rect 23204 4471 23256 4480
rect 23204 4437 23213 4471
rect 23213 4437 23247 4471
rect 23247 4437 23256 4471
rect 24492 4471 24544 4480
rect 23204 4428 23256 4437
rect 24492 4437 24501 4471
rect 24501 4437 24535 4471
rect 24535 4437 24544 4471
rect 24492 4428 24544 4437
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 4528 4224 4580 4276
rect 4896 4224 4948 4276
rect 5264 4267 5316 4276
rect 5264 4233 5273 4267
rect 5273 4233 5307 4267
rect 5307 4233 5316 4267
rect 5264 4224 5316 4233
rect 7104 4267 7156 4276
rect 7104 4233 7113 4267
rect 7113 4233 7147 4267
rect 7147 4233 7156 4267
rect 7104 4224 7156 4233
rect 12256 4224 12308 4276
rect 13820 4224 13872 4276
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2964 4156 3016 4208
rect 5908 4156 5960 4208
rect 7472 4156 7524 4208
rect 2780 4088 2832 4140
rect 3332 4063 3384 4072
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 3976 4063 4028 4072
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 5724 4020 5776 4029
rect 8116 4020 8168 4072
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 4988 3952 5040 4004
rect 5632 3952 5684 4004
rect 7380 3952 7432 4004
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 4436 3927 4488 3936
rect 4436 3893 4445 3927
rect 4445 3893 4479 3927
rect 4479 3893 4488 3927
rect 4436 3884 4488 3893
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 7472 3884 7524 3936
rect 7840 3927 7892 3936
rect 7840 3893 7849 3927
rect 7849 3893 7883 3927
rect 7883 3893 7892 3927
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 10968 4088 11020 4140
rect 11796 4088 11848 4140
rect 12992 4131 13044 4140
rect 8484 4020 8536 4029
rect 9956 4020 10008 4072
rect 10140 4063 10192 4072
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 10140 4020 10192 4029
rect 10692 4020 10744 4072
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 12716 4020 12768 4072
rect 15108 4088 15160 4140
rect 14924 4020 14976 4072
rect 16948 4224 17000 4276
rect 18052 4224 18104 4276
rect 19892 4267 19944 4276
rect 19892 4233 19901 4267
rect 19901 4233 19935 4267
rect 19935 4233 19944 4267
rect 19892 4224 19944 4233
rect 24032 4267 24084 4276
rect 24032 4233 24041 4267
rect 24041 4233 24075 4267
rect 24075 4233 24084 4267
rect 24032 4224 24084 4233
rect 25780 4267 25832 4276
rect 25780 4233 25789 4267
rect 25789 4233 25823 4267
rect 25823 4233 25832 4267
rect 25780 4224 25832 4233
rect 27160 4224 27212 4276
rect 28264 4224 28316 4276
rect 30196 4267 30248 4276
rect 30196 4233 30205 4267
rect 30205 4233 30239 4267
rect 30239 4233 30248 4267
rect 30196 4224 30248 4233
rect 35440 4224 35492 4276
rect 16580 4156 16632 4208
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 17040 4131 17092 4140
rect 16764 4088 16816 4097
rect 17040 4097 17049 4131
rect 17049 4097 17083 4131
rect 17083 4097 17092 4131
rect 17040 4088 17092 4097
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 16396 4063 16448 4072
rect 16396 4029 16405 4063
rect 16405 4029 16439 4063
rect 16439 4029 16448 4063
rect 16396 4020 16448 4029
rect 16488 4020 16540 4072
rect 17960 4020 18012 4072
rect 9036 3952 9088 4004
rect 16304 3952 16356 4004
rect 17776 3952 17828 4004
rect 19248 4020 19300 4072
rect 22836 4088 22888 4140
rect 25136 4156 25188 4208
rect 28172 4156 28224 4208
rect 20904 4020 20956 4072
rect 21640 4063 21692 4072
rect 21640 4029 21649 4063
rect 21649 4029 21683 4063
rect 21683 4029 21692 4063
rect 21640 4020 21692 4029
rect 22284 4063 22336 4072
rect 22284 4029 22293 4063
rect 22293 4029 22327 4063
rect 22327 4029 22336 4063
rect 22284 4020 22336 4029
rect 18788 3995 18840 4004
rect 18788 3961 18797 3995
rect 18797 3961 18831 3995
rect 18831 3961 18840 3995
rect 18788 3952 18840 3961
rect 20720 3952 20772 4004
rect 22928 4020 22980 4072
rect 23940 4020 23992 4072
rect 24492 4063 24544 4072
rect 24492 4029 24501 4063
rect 24501 4029 24535 4063
rect 24535 4029 24544 4063
rect 24492 4020 24544 4029
rect 26424 4088 26476 4140
rect 28080 4088 28132 4140
rect 27804 4063 27856 4072
rect 27804 4029 27813 4063
rect 27813 4029 27847 4063
rect 27847 4029 27856 4063
rect 27804 4020 27856 4029
rect 29828 4063 29880 4072
rect 29828 4029 29837 4063
rect 29837 4029 29871 4063
rect 29871 4029 29880 4063
rect 29828 4020 29880 4029
rect 30288 4063 30340 4072
rect 30288 4029 30297 4063
rect 30297 4029 30331 4063
rect 30331 4029 30340 4063
rect 30288 4020 30340 4029
rect 23388 3952 23440 4004
rect 25044 3952 25096 4004
rect 26424 3995 26476 4004
rect 26424 3961 26433 3995
rect 26433 3961 26467 3995
rect 26467 3961 26476 3995
rect 26976 3995 27028 4004
rect 26424 3952 26476 3961
rect 26976 3961 26985 3995
rect 26985 3961 27019 3995
rect 27019 3961 27028 3995
rect 26976 3952 27028 3961
rect 7840 3884 7892 3893
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 10876 3884 10928 3936
rect 11612 3884 11664 3936
rect 13728 3884 13780 3936
rect 14004 3927 14056 3936
rect 14004 3893 14013 3927
rect 14013 3893 14047 3927
rect 14047 3893 14056 3927
rect 14004 3884 14056 3893
rect 15200 3884 15252 3936
rect 16764 3884 16816 3936
rect 21088 3927 21140 3936
rect 21088 3893 21097 3927
rect 21097 3893 21131 3927
rect 21131 3893 21140 3927
rect 21088 3884 21140 3893
rect 21640 3884 21692 3936
rect 22008 3884 22060 3936
rect 22652 3884 22704 3936
rect 23296 3884 23348 3936
rect 26240 3884 26292 3936
rect 27160 3884 27212 3936
rect 30472 3927 30524 3936
rect 30472 3893 30481 3927
rect 30481 3893 30515 3927
rect 30515 3893 30524 3927
rect 30472 3884 30524 3893
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 1952 3680 2004 3732
rect 2780 3680 2832 3732
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 3700 3680 3752 3732
rect 5356 3680 5408 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6552 3723 6604 3732
rect 6552 3689 6561 3723
rect 6561 3689 6595 3723
rect 6595 3689 6604 3723
rect 6552 3680 6604 3689
rect 8116 3680 8168 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 9220 3723 9272 3732
rect 9220 3689 9229 3723
rect 9229 3689 9263 3723
rect 9263 3689 9272 3723
rect 9220 3680 9272 3689
rect 9680 3680 9732 3732
rect 10140 3680 10192 3732
rect 12624 3680 12676 3732
rect 15292 3680 15344 3732
rect 15844 3723 15896 3732
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17592 3723 17644 3732
rect 17592 3689 17601 3723
rect 17601 3689 17635 3723
rect 17635 3689 17644 3723
rect 17592 3680 17644 3689
rect 4344 3612 4396 3664
rect 7196 3612 7248 3664
rect 8392 3612 8444 3664
rect 9956 3612 10008 3664
rect 12256 3655 12308 3664
rect 4160 3587 4212 3596
rect 4160 3553 4178 3587
rect 4178 3553 4212 3587
rect 4160 3544 4212 3553
rect 4804 3544 4856 3596
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 7380 3587 7432 3596
rect 7380 3553 7389 3587
rect 7389 3553 7423 3587
rect 7423 3553 7432 3587
rect 7380 3544 7432 3553
rect 7104 3476 7156 3528
rect 7840 3544 7892 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 10324 3544 10376 3596
rect 12256 3621 12265 3655
rect 12265 3621 12299 3655
rect 12299 3621 12308 3655
rect 12256 3612 12308 3621
rect 8208 3476 8260 3528
rect 11796 3544 11848 3596
rect 12716 3544 12768 3596
rect 14832 3612 14884 3664
rect 17868 3680 17920 3732
rect 18880 3680 18932 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 20812 3680 20864 3732
rect 23940 3723 23992 3732
rect 19892 3655 19944 3664
rect 19892 3621 19901 3655
rect 19901 3621 19935 3655
rect 19935 3621 19944 3655
rect 19892 3612 19944 3621
rect 23940 3689 23949 3723
rect 23949 3689 23983 3723
rect 23983 3689 23992 3723
rect 23940 3680 23992 3689
rect 29092 3680 29144 3732
rect 25044 3612 25096 3664
rect 28356 3612 28408 3664
rect 14372 3587 14424 3596
rect 13176 3476 13228 3528
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 17960 3587 18012 3596
rect 17960 3553 17966 3587
rect 17966 3553 18012 3587
rect 17960 3544 18012 3553
rect 18512 3544 18564 3596
rect 19340 3587 19392 3596
rect 19340 3553 19349 3587
rect 19349 3553 19383 3587
rect 19383 3553 19392 3587
rect 19340 3544 19392 3553
rect 19524 3587 19576 3596
rect 19524 3553 19533 3587
rect 19533 3553 19567 3587
rect 19567 3553 19576 3587
rect 19524 3544 19576 3553
rect 20904 3587 20956 3596
rect 20904 3553 20913 3587
rect 20913 3553 20947 3587
rect 20947 3553 20956 3587
rect 20904 3544 20956 3553
rect 14648 3476 14700 3528
rect 17776 3476 17828 3528
rect 20720 3476 20772 3528
rect 21824 3544 21876 3596
rect 22836 3587 22888 3596
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 23112 3544 23164 3596
rect 23848 3587 23900 3596
rect 23848 3553 23857 3587
rect 23857 3553 23891 3587
rect 23891 3553 23900 3587
rect 23848 3544 23900 3553
rect 24860 3587 24912 3596
rect 24860 3553 24869 3587
rect 24869 3553 24903 3587
rect 24903 3553 24912 3587
rect 24860 3544 24912 3553
rect 26424 3544 26476 3596
rect 22284 3476 22336 3528
rect 27988 3476 28040 3528
rect 29552 3519 29604 3528
rect 29552 3485 29561 3519
rect 29561 3485 29595 3519
rect 29595 3485 29604 3519
rect 29552 3476 29604 3485
rect 16580 3408 16632 3460
rect 17960 3408 18012 3460
rect 8116 3340 8168 3392
rect 15200 3340 15252 3392
rect 18328 3408 18380 3460
rect 30104 3451 30156 3460
rect 30104 3417 30113 3451
rect 30113 3417 30147 3451
rect 30147 3417 30156 3451
rect 30104 3408 30156 3417
rect 22468 3340 22520 3392
rect 24584 3383 24636 3392
rect 24584 3349 24593 3383
rect 24593 3349 24627 3383
rect 24627 3349 24636 3383
rect 24584 3340 24636 3349
rect 25228 3383 25280 3392
rect 25228 3349 25237 3383
rect 25237 3349 25271 3383
rect 25271 3349 25280 3383
rect 25228 3340 25280 3349
rect 26240 3383 26292 3392
rect 26240 3349 26249 3383
rect 26249 3349 26283 3383
rect 26283 3349 26292 3383
rect 26240 3340 26292 3349
rect 26332 3340 26384 3392
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 3240 3136 3292 3188
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 4804 3136 4856 3188
rect 6368 3136 6420 3188
rect 3700 3068 3752 3120
rect 6000 3068 6052 3120
rect 6276 3111 6328 3120
rect 6276 3077 6285 3111
rect 6285 3077 6319 3111
rect 6319 3077 6328 3111
rect 6276 3068 6328 3077
rect 8116 3136 8168 3188
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 3884 3000 3936 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 2136 2932 2188 2984
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 6920 3000 6972 3052
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 7840 2932 7892 2984
rect 9864 3136 9916 3188
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 12348 3136 12400 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 14004 3136 14056 3188
rect 14924 3136 14976 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16764 3136 16816 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18512 3179 18564 3188
rect 18512 3145 18521 3179
rect 18521 3145 18555 3179
rect 18555 3145 18564 3179
rect 18512 3136 18564 3145
rect 19340 3136 19392 3188
rect 21732 3136 21784 3188
rect 22100 3136 22152 3188
rect 23112 3179 23164 3188
rect 23112 3145 23121 3179
rect 23121 3145 23155 3179
rect 23155 3145 23164 3179
rect 23112 3136 23164 3145
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 26424 3136 26476 3188
rect 27252 3179 27304 3188
rect 27252 3145 27261 3179
rect 27261 3145 27295 3179
rect 27295 3145 27304 3179
rect 27252 3136 27304 3145
rect 27988 3136 28040 3188
rect 29552 3136 29604 3188
rect 9680 3068 9732 3120
rect 11796 3111 11848 3120
rect 11796 3077 11805 3111
rect 11805 3077 11839 3111
rect 11839 3077 11848 3111
rect 11796 3068 11848 3077
rect 11980 3068 12032 3120
rect 12164 3111 12216 3120
rect 12164 3077 12173 3111
rect 12173 3077 12207 3111
rect 12207 3077 12216 3111
rect 12164 3068 12216 3077
rect 14372 3068 14424 3120
rect 16580 3068 16632 3120
rect 22468 3111 22520 3120
rect 22468 3077 22477 3111
rect 22477 3077 22511 3111
rect 22511 3077 22520 3111
rect 22468 3068 22520 3077
rect 23848 3068 23900 3120
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 9588 2932 9640 2984
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 17868 3000 17920 3052
rect 26332 3043 26384 3052
rect 26332 3009 26341 3043
rect 26341 3009 26375 3043
rect 26375 3009 26384 3043
rect 26332 3000 26384 3009
rect 26976 3043 27028 3052
rect 26976 3009 26985 3043
rect 26985 3009 27019 3043
rect 27019 3009 27028 3043
rect 26976 3000 27028 3009
rect 29460 3043 29512 3052
rect 29460 3009 29469 3043
rect 29469 3009 29503 3043
rect 29503 3009 29512 3043
rect 29460 3000 29512 3009
rect 30104 3043 30156 3052
rect 30104 3009 30113 3043
rect 30113 3009 30147 3043
rect 30147 3009 30156 3043
rect 30104 3000 30156 3009
rect 15016 2975 15068 2984
rect 15016 2941 15022 2975
rect 15022 2941 15068 2975
rect 15016 2932 15068 2941
rect 16304 2932 16356 2984
rect 16672 2975 16724 2984
rect 16672 2941 16681 2975
rect 16681 2941 16715 2975
rect 16715 2941 16724 2975
rect 16672 2932 16724 2941
rect 18328 2932 18380 2984
rect 20260 2932 20312 2984
rect 20812 2975 20864 2984
rect 20812 2941 20821 2975
rect 20821 2941 20855 2975
rect 20855 2941 20864 2975
rect 20812 2932 20864 2941
rect 21732 2975 21784 2984
rect 8392 2864 8444 2916
rect 14832 2907 14884 2916
rect 14832 2873 14841 2907
rect 14841 2873 14875 2907
rect 14875 2873 14884 2907
rect 14832 2864 14884 2873
rect 21732 2941 21741 2975
rect 21741 2941 21775 2975
rect 21775 2941 21784 2975
rect 21732 2932 21784 2941
rect 22008 2975 22060 2984
rect 22008 2941 22017 2975
rect 22017 2941 22051 2975
rect 22051 2941 22060 2975
rect 22008 2932 22060 2941
rect 22560 2932 22612 2984
rect 23296 2932 23348 2984
rect 24584 2932 24636 2984
rect 27068 2932 27120 2984
rect 21088 2864 21140 2916
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 18420 2796 18472 2848
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 19156 2796 19208 2805
rect 20996 2796 21048 2848
rect 21824 2864 21876 2916
rect 23112 2864 23164 2916
rect 23756 2864 23808 2916
rect 25044 2864 25096 2916
rect 26516 2864 26568 2916
rect 27620 2864 27672 2916
rect 29552 2907 29604 2916
rect 29552 2873 29561 2907
rect 29561 2873 29595 2907
rect 29595 2873 29604 2907
rect 29552 2864 29604 2873
rect 23480 2796 23532 2848
rect 24860 2839 24912 2848
rect 24860 2805 24869 2839
rect 24869 2805 24903 2839
rect 24903 2805 24912 2839
rect 24860 2796 24912 2805
rect 28356 2839 28408 2848
rect 28356 2805 28365 2839
rect 28365 2805 28399 2839
rect 28399 2805 28408 2839
rect 28356 2796 28408 2805
rect 29828 2796 29880 2848
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 2688 2592 2740 2644
rect 8116 2635 8168 2644
rect 8116 2601 8125 2635
rect 8125 2601 8159 2635
rect 8159 2601 8168 2635
rect 8116 2592 8168 2601
rect 8392 2592 8444 2644
rect 8852 2635 8904 2644
rect 8852 2601 8861 2635
rect 8861 2601 8895 2635
rect 8895 2601 8904 2635
rect 8852 2592 8904 2601
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11888 2592 11940 2644
rect 13636 2592 13688 2644
rect 14924 2635 14976 2644
rect 14924 2601 14933 2635
rect 14933 2601 14967 2635
rect 14967 2601 14976 2635
rect 14924 2592 14976 2601
rect 16304 2592 16356 2644
rect 16764 2592 16816 2644
rect 17960 2635 18012 2644
rect 17960 2601 17969 2635
rect 17969 2601 18003 2635
rect 18003 2601 18012 2635
rect 17960 2592 18012 2601
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 7840 2567 7892 2576
rect 7840 2533 7849 2567
rect 7849 2533 7883 2567
rect 7883 2533 7892 2567
rect 7840 2524 7892 2533
rect 2228 2499 2280 2508
rect 2228 2465 2272 2499
rect 2272 2465 2280 2499
rect 2228 2456 2280 2465
rect 6092 2456 6144 2508
rect 7104 2456 7156 2508
rect 8300 2456 8352 2508
rect 14648 2524 14700 2576
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 11520 2499 11572 2508
rect 11520 2465 11564 2499
rect 11564 2465 11572 2499
rect 11520 2456 11572 2465
rect 12900 2499 12952 2508
rect 12900 2465 12902 2499
rect 12902 2465 12952 2499
rect 13360 2499 13412 2508
rect 12900 2456 12952 2465
rect 13360 2465 13369 2499
rect 13369 2465 13403 2499
rect 13403 2465 13412 2499
rect 13360 2456 13412 2465
rect 14740 2456 14792 2508
rect 19248 2592 19300 2644
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 23756 2635 23808 2644
rect 20628 2524 20680 2576
rect 21088 2524 21140 2576
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 25228 2635 25280 2644
rect 23388 2524 23440 2576
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 26240 2592 26292 2644
rect 29092 2635 29144 2644
rect 29092 2601 29101 2635
rect 29101 2601 29135 2635
rect 29135 2601 29144 2635
rect 29092 2592 29144 2601
rect 29460 2635 29512 2644
rect 29460 2601 29469 2635
rect 29469 2601 29503 2635
rect 29503 2601 29512 2635
rect 29460 2592 29512 2601
rect 21272 2499 21324 2508
rect 21272 2465 21290 2499
rect 21290 2465 21324 2499
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16672 2388 16724 2440
rect 21272 2456 21324 2465
rect 26332 2456 26384 2508
rect 27436 2456 27488 2508
rect 27896 2499 27948 2508
rect 27896 2465 27940 2499
rect 27940 2465 27948 2499
rect 27896 2456 27948 2465
rect 29552 2524 29604 2576
rect 29828 2499 29880 2508
rect 29828 2465 29837 2499
rect 29837 2465 29871 2499
rect 29871 2465 29880 2499
rect 29828 2456 29880 2465
rect 30380 2456 30432 2508
rect 22468 2431 22520 2440
rect 8300 2320 8352 2372
rect 20260 2320 20312 2372
rect 22468 2397 22477 2431
rect 22477 2397 22511 2431
rect 22511 2397 22520 2431
rect 22468 2388 22520 2397
rect 21364 2320 21416 2372
rect 24768 2363 24820 2372
rect 24768 2329 24777 2363
rect 24777 2329 24811 2363
rect 24811 2329 24820 2363
rect 24768 2320 24820 2329
rect 26240 2363 26292 2372
rect 26240 2329 26249 2363
rect 26249 2329 26283 2363
rect 26283 2329 26292 2363
rect 26240 2320 26292 2329
rect 26516 2295 26568 2304
rect 26516 2261 26525 2295
rect 26525 2261 26559 2295
rect 26559 2261 26568 2295
rect 26516 2252 26568 2261
rect 27436 2295 27488 2304
rect 27436 2261 27445 2295
rect 27445 2261 27479 2295
rect 27479 2261 27488 2295
rect 27436 2252 27488 2261
rect 28908 2252 28960 2304
rect 31668 2252 31720 2304
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 18052 552 18104 604
rect 18328 552 18380 604
<< metal2 >>
rect 2502 15520 2558 16000
rect 2686 15600 2742 15609
rect 2686 15535 2742 15544
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1490 13832 1546 13841
rect 1490 13767 1546 13776
rect 1504 12986 1532 13767
rect 1596 13530 1624 14583
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1688 12986 1716 13330
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 1582 12064 1638 12073
rect 1582 11999 1638 12008
rect 1596 11898 1624 11999
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 2056 11830 2084 12242
rect 2044 11824 2096 11830
rect 2042 11792 2044 11801
rect 2096 11792 2098 11801
rect 2042 11727 2098 11736
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1582 11112 1638 11121
rect 1582 11047 1584 11056
rect 1636 11047 1638 11056
rect 1584 11018 1636 11024
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10305 1624 10406
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1688 10062 1716 11154
rect 2148 10606 2176 12582
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2044 10464 2096 10470
rect 2042 10432 2044 10441
rect 2096 10432 2098 10441
rect 2042 10367 2098 10376
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1676 10056 1728 10062
rect 1674 10024 1676 10033
rect 1728 10024 1730 10033
rect 1674 9959 1730 9968
rect 1490 9072 1546 9081
rect 1490 9007 1492 9016
rect 1544 9007 1546 9016
rect 1492 8978 1544 8984
rect 1504 8634 1532 8978
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1582 8528 1638 8537
rect 1582 8463 1638 8472
rect 1596 6458 1624 8463
rect 1780 7954 1808 10202
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2148 9382 2176 10066
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1872 8498 1900 8774
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1780 7002 1808 7890
rect 1768 6996 1820 7002
rect 1768 6938 1820 6944
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1688 5574 1716 6122
rect 2044 5840 2096 5846
rect 2044 5782 2096 5788
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1688 5098 1716 5510
rect 2056 5370 2084 5782
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1688 4282 1716 4626
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1780 3738 1808 5102
rect 2056 4826 2084 5306
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1964 4146 1992 4422
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 1964 3738 1992 4082
rect 2056 4010 2084 4762
rect 2044 4004 2096 4010
rect 2044 3946 2096 3952
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3505 1992 3538
rect 1950 3496 2006 3505
rect 1950 3431 2006 3440
rect 1964 2990 1992 3431
rect 2148 2990 2176 9318
rect 2240 7313 2268 11698
rect 2332 9586 2360 12038
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11257 2452 11494
rect 2410 11248 2466 11257
rect 2410 11183 2466 11192
rect 2516 10305 2544 15520
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2502 10296 2558 10305
rect 2502 10231 2558 10240
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9654 2452 10066
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2424 8922 2452 9386
rect 2608 9194 2636 11494
rect 2700 11354 2728 15535
rect 7470 15520 7526 16000
rect 12438 15520 12494 16000
rect 17498 15520 17554 16000
rect 22466 15520 22522 16000
rect 27434 15520 27490 16000
rect 32494 15520 32550 16000
rect 36634 15600 36690 15609
rect 36634 15535 36690 15544
rect 3790 12880 3846 12889
rect 3790 12815 3846 12824
rect 3804 12646 3832 12815
rect 3792 12640 3844 12646
rect 3792 12582 3844 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2700 9489 2728 10406
rect 2686 9480 2742 9489
rect 2686 9415 2742 9424
rect 2332 8894 2452 8922
rect 2516 9166 2636 9194
rect 2332 8838 2360 8894
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8362 2360 8774
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2226 7304 2282 7313
rect 2226 7239 2282 7248
rect 2240 6458 2268 7239
rect 2332 7206 2360 7958
rect 2320 7200 2372 7206
rect 2320 7142 2372 7148
rect 2332 6934 2360 7142
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 6186 2360 6870
rect 2516 6322 2544 9166
rect 2792 9160 2820 12038
rect 2962 11792 3018 11801
rect 2962 11727 3018 11736
rect 2700 9132 2820 9160
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2608 8634 2636 9046
rect 2700 8974 2728 9132
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2700 8498 2728 8910
rect 2884 8566 2912 8910
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 8090 2728 8298
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2608 5574 2636 6734
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 6118 2820 6598
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2608 3058 2636 5510
rect 2688 4752 2740 4758
rect 2792 4706 2820 6054
rect 2976 5658 3004 11727
rect 3160 11558 3188 12242
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3056 10600 3108 10606
rect 3054 10568 3056 10577
rect 3108 10568 3110 10577
rect 3054 10503 3110 10512
rect 3160 10169 3188 11494
rect 4802 11248 4858 11257
rect 4802 11183 4804 11192
rect 4856 11183 4858 11192
rect 4804 11154 4856 11160
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10470 3464 10950
rect 3424 10464 3476 10470
rect 4068 10464 4120 10470
rect 3424 10406 3476 10412
rect 3882 10432 3938 10441
rect 3146 10160 3202 10169
rect 3068 10118 3146 10146
rect 3068 7585 3096 10118
rect 3146 10095 3202 10104
rect 3332 9444 3384 9450
rect 3332 9386 3384 9392
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3054 7576 3110 7585
rect 3160 7546 3188 8570
rect 3344 8362 3372 9386
rect 3436 9081 3464 10406
rect 4068 10406 4120 10412
rect 3882 10367 3938 10376
rect 3422 9072 3478 9081
rect 3422 9007 3478 9016
rect 3896 8945 3924 10367
rect 3974 9344 4030 9353
rect 3974 9279 4030 9288
rect 3882 8936 3938 8945
rect 3882 8871 3938 8880
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3054 7511 3110 7520
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3160 6186 3188 7482
rect 3344 6730 3372 8298
rect 3790 7984 3846 7993
rect 3790 7919 3846 7928
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7342 3556 7686
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 6390 3372 6666
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3436 6322 3464 6598
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 3160 5914 3188 6122
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2740 4700 2820 4706
rect 2688 4694 2820 4700
rect 2700 4678 2820 4694
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 3754 2728 4558
rect 2792 4146 2820 4678
rect 2884 5630 3004 5658
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2884 4049 2912 5630
rect 2962 5536 3018 5545
rect 2962 5471 3018 5480
rect 2976 4622 3004 5471
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2976 4214 3004 4558
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2870 4040 2926 4049
rect 2870 3975 2926 3984
rect 2962 3904 3018 3913
rect 2962 3839 3018 3848
rect 2700 3738 2820 3754
rect 2700 3732 2832 3738
rect 2700 3726 2780 3732
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 1964 2650 1992 2926
rect 2700 2650 2728 3726
rect 2780 3674 2832 3680
rect 2976 2990 3004 3839
rect 3252 3194 3280 4966
rect 3332 4072 3384 4078
rect 3330 4040 3332 4049
rect 3384 4040 3386 4049
rect 3330 3975 3386 3984
rect 3528 3942 3556 7278
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3620 6934 3648 7142
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3620 5030 3648 6870
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3712 4826 3740 5102
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3712 3777 3740 4014
rect 3698 3768 3754 3777
rect 3698 3703 3700 3712
rect 3752 3703 3754 3712
rect 3700 3674 3752 3680
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3712 3126 3740 3674
rect 3700 3120 3752 3126
rect 3804 3097 3832 7919
rect 3700 3062 3752 3068
rect 3790 3088 3846 3097
rect 3896 3058 3924 8871
rect 3988 8634 4016 9279
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4080 6798 4108 10406
rect 4158 10296 4214 10305
rect 4158 10231 4160 10240
rect 4212 10231 4214 10240
rect 4160 10202 4212 10208
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 8090 4200 9318
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4172 7410 4200 8026
rect 4264 7886 4292 11018
rect 4816 10810 4844 11154
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4528 9512 4580 9518
rect 4342 9480 4398 9489
rect 4342 9415 4398 9424
rect 4526 9480 4528 9489
rect 4620 9512 4672 9518
rect 4580 9480 4582 9489
rect 4620 9454 4672 9460
rect 4526 9415 4582 9424
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4172 6458 4200 6802
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4356 6322 4384 9415
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4448 6934 4476 7958
rect 4436 6928 4488 6934
rect 4436 6870 4488 6876
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5914 4384 6258
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4172 5166 4200 5646
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3976 4072 4028 4078
rect 3974 4040 3976 4049
rect 4028 4040 4030 4049
rect 3974 3975 4030 3984
rect 4356 3670 4384 5510
rect 4540 4690 4568 9415
rect 4632 9217 4660 9454
rect 4618 9208 4674 9217
rect 4618 9143 4674 9152
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 4632 6186 4660 6258
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4632 5710 4660 6122
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4436 4616 4488 4622
rect 4436 4558 4488 4564
rect 4448 3942 4476 4558
rect 4540 4282 4568 4626
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 3194 4200 3538
rect 4448 3505 4476 3878
rect 4434 3496 4490 3505
rect 4434 3431 4490 3440
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 3790 3023 3846 3032
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 1674 2408 1730 2417
rect 1674 2343 1730 2352
rect 1688 480 1716 2343
rect 2240 2281 2268 2450
rect 2226 2272 2282 2281
rect 2226 2207 2282 2216
rect 4172 2009 4200 3130
rect 4724 3097 4752 10406
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5184 9722 5212 10066
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8022 4844 8910
rect 5092 8378 5120 9046
rect 5184 8974 5212 9658
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8566 5212 8910
rect 5172 8560 5224 8566
rect 5172 8502 5224 8508
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5170 8392 5226 8401
rect 5092 8350 5170 8378
rect 5368 8362 5396 8434
rect 5170 8327 5226 8336
rect 5356 8356 5408 8362
rect 4896 8288 4948 8294
rect 4896 8230 4948 8236
rect 4804 8016 4856 8022
rect 4804 7958 4856 7964
rect 4802 5808 4858 5817
rect 4802 5743 4858 5752
rect 4816 3602 4844 5743
rect 4908 5273 4936 8230
rect 5184 8090 5212 8327
rect 5356 8298 5408 8304
rect 5368 8265 5396 8298
rect 5540 8288 5592 8294
rect 5354 8256 5410 8265
rect 5540 8230 5592 8236
rect 5354 8191 5410 8200
rect 5552 8090 5580 8230
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5644 7857 5672 9454
rect 5828 8090 5856 12582
rect 7484 11121 7512 15520
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 8942 11520 8998 11529
rect 8942 11455 8998 11464
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 5906 11112 5962 11121
rect 5906 11047 5962 11056
rect 7470 11112 7526 11121
rect 7470 11047 7526 11056
rect 8114 11112 8170 11121
rect 8114 11047 8170 11056
rect 5920 9654 5948 11047
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5630 7848 5686 7857
rect 5630 7783 5686 7792
rect 5736 7546 5764 7890
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 5092 6934 5120 7142
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5276 6458 5304 6734
rect 5552 6458 5580 7210
rect 5736 7041 5764 7482
rect 5722 7032 5778 7041
rect 5722 6967 5778 6976
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5906 6352 5962 6361
rect 5906 6287 5962 6296
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 4894 5264 4950 5273
rect 4894 5199 4950 5208
rect 4908 4554 4936 5199
rect 5552 4690 5580 5646
rect 5828 5370 5856 5782
rect 5920 5370 5948 6287
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6012 5545 6040 5646
rect 5998 5536 6054 5545
rect 5998 5471 6054 5480
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5540 4684 5592 4690
rect 5368 4644 5540 4672
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5276 4282 5304 4490
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4816 3194 4844 3538
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4250 3088 4306 3097
rect 4250 3023 4306 3032
rect 4710 3088 4766 3097
rect 4710 3023 4766 3032
rect 4158 2000 4214 2009
rect 4158 1935 4214 1944
rect 4172 1329 4200 1935
rect 4158 1320 4214 1329
rect 4158 1255 4214 1264
rect 4264 513 4292 3023
rect 4908 2689 4936 4218
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4894 2680 4950 2689
rect 4894 2615 4950 2624
rect 4250 504 4306 513
rect 1674 0 1730 480
rect 5000 480 5028 3946
rect 5368 3738 5396 4644
rect 5540 4626 5592 4632
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5644 4010 5672 4626
rect 5920 4214 5948 4626
rect 5908 4208 5960 4214
rect 5722 4176 5778 4185
rect 5908 4150 5960 4156
rect 5722 4111 5778 4120
rect 5736 4078 5764 4111
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5998 4040 6054 4049
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 3738 5764 4014
rect 5998 3975 6054 3984
rect 5908 3936 5960 3942
rect 5906 3904 5908 3913
rect 5960 3904 5962 3913
rect 5906 3839 5962 3848
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 6012 3126 6040 3975
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6104 2514 6132 8230
rect 6196 3505 6224 9318
rect 6564 9110 6592 10406
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6564 8634 6592 9046
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8090 6684 9046
rect 6748 8537 6776 9998
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6734 8528 6790 8537
rect 6734 8463 6790 8472
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6656 6458 6684 6802
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4758 6408 5102
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6274 4584 6330 4593
rect 6274 4519 6330 4528
rect 6182 3496 6238 3505
rect 6182 3431 6238 3440
rect 6288 3126 6316 4519
rect 6656 4049 6684 5306
rect 6748 4826 6776 7278
rect 6840 6798 6868 9318
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6932 8498 6960 9114
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7208 8022 7236 8298
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7206 6960 7822
rect 7208 7206 7236 7958
rect 7300 7449 7328 9454
rect 7392 9382 7420 10066
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 7380 9376 7432 9382
rect 7840 9376 7892 9382
rect 7380 9318 7432 9324
rect 7838 9344 7840 9353
rect 7892 9344 7894 9353
rect 7392 8294 7420 9318
rect 7838 9279 7894 9288
rect 8128 9042 8156 11047
rect 8588 10810 8616 11154
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9625 8248 9862
rect 8206 9616 8262 9625
rect 8206 9551 8262 9560
rect 8404 9382 8432 10066
rect 8588 9489 8616 10746
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9722 8892 9862
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8574 9480 8630 9489
rect 8574 9415 8630 9424
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8298 9208 8354 9217
rect 8298 9143 8354 9152
rect 8312 9042 8340 9143
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 8128 8634 8156 8978
rect 8206 8800 8262 8809
rect 8206 8735 8262 8744
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7840 8424 7892 8430
rect 7838 8392 7840 8401
rect 7892 8392 7894 8401
rect 7838 8327 7894 8336
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 5914 6868 6734
rect 6932 5914 6960 7142
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 6322 7052 6598
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 6186 7052 6258
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7116 5846 7144 7142
rect 7208 6934 7236 7142
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 5370 6868 5646
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 7208 5302 7236 6870
rect 7300 5370 7328 7375
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 6662 8064 7278
rect 8220 6905 8248 8735
rect 8312 8634 8340 8978
rect 8404 8809 8432 9318
rect 8772 8838 8800 9386
rect 8850 8936 8906 8945
rect 8850 8871 8906 8880
rect 8760 8832 8812 8838
rect 8390 8800 8446 8809
rect 8760 8774 8812 8780
rect 8390 8735 8446 8744
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8206 6896 8262 6905
rect 8206 6831 8262 6840
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8312 6458 8340 8570
rect 8864 8430 8892 8871
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8758 8256 8814 8265
rect 8758 8191 8814 8200
rect 8772 7546 8800 8191
rect 8956 8090 8984 11455
rect 9140 10606 9168 12922
rect 11336 12300 11388 12306
rect 11336 12242 11388 12248
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11762 10180 12038
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 9692 10962 9720 11698
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 11082 10088 11154
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10060 10985 10088 11018
rect 9600 10934 9720 10962
rect 10046 10976 10102 10985
rect 9600 10742 9628 10934
rect 10046 10911 10102 10920
rect 9954 10840 10010 10849
rect 9954 10775 10010 10784
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9968 10606 9996 10775
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9586 9076 9862
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 8634 9076 9522
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 9048 7410 9076 7890
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8758 7168 8814 7177
rect 8758 7103 8814 7112
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8312 6186 8340 6394
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8312 5778 8340 6122
rect 8496 6118 8524 6598
rect 8680 6474 8708 6802
rect 8772 6730 8800 7103
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 9048 6662 9076 7346
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8680 6446 8800 6474
rect 8666 6352 8722 6361
rect 8666 6287 8722 6296
rect 8680 6254 8708 6287
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8680 5914 8708 6190
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8772 5574 8800 6446
rect 9048 6322 9076 6598
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9140 5817 9168 5850
rect 9126 5808 9182 5817
rect 9126 5743 9182 5752
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6840 4978 6868 5034
rect 6840 4950 6960 4978
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6550 3768 6606 3777
rect 6550 3703 6552 3712
rect 6604 3703 6606 3712
rect 6552 3674 6604 3680
rect 6366 3632 6422 3641
rect 6366 3567 6368 3576
rect 6420 3567 6422 3576
rect 6368 3538 6420 3544
rect 6380 3194 6408 3538
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6932 3058 6960 4950
rect 8220 4758 8248 5102
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7472 4684 7524 4690
rect 7472 4626 7524 4632
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 4282 7144 4490
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7208 3670 7236 4626
rect 7484 4214 7512 4626
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7378 4040 7434 4049
rect 7378 3975 7380 3984
rect 7432 3975 7434 3984
rect 7380 3946 7432 3952
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7392 3602 7420 3946
rect 7484 3942 7512 4150
rect 8404 4078 8432 4422
rect 8496 4078 8524 4490
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7840 3936 7892 3942
rect 7840 3878 7892 3884
rect 7852 3602 7880 3878
rect 8128 3738 8156 4014
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7116 2854 7144 3470
rect 7392 2990 7420 3538
rect 8128 3398 8156 3674
rect 8404 3670 8432 4014
rect 8496 3738 8524 4014
rect 8772 3913 8800 5510
rect 9126 5400 9182 5409
rect 9126 5335 9128 5344
rect 9180 5335 9182 5344
rect 9128 5306 9180 5312
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8852 3936 8904 3942
rect 8758 3904 8814 3913
rect 8852 3878 8904 3884
rect 8758 3839 8814 3848
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8392 3664 8444 3670
rect 8864 3641 8892 3878
rect 9048 3641 9076 3946
rect 9232 3777 9260 10406
rect 10060 10266 10088 10911
rect 10048 10260 10100 10266
rect 9678 10194 9734 10203
rect 10048 10202 10100 10208
rect 9678 10129 9734 10138
rect 9310 10024 9366 10033
rect 9692 9994 9720 10129
rect 9310 9959 9366 9968
rect 9680 9988 9732 9994
rect 9324 9586 9352 9959
rect 9680 9930 9732 9936
rect 9678 9888 9734 9897
rect 9678 9823 9734 9832
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9692 9042 9720 9823
rect 10152 9586 10180 11290
rect 10704 11218 10732 11494
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10538 10272 10950
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 8634 9720 8978
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9678 8528 9734 8537
rect 9678 8463 9734 8472
rect 9496 8424 9548 8430
rect 9494 8392 9496 8401
rect 9548 8392 9550 8401
rect 9494 8327 9550 8336
rect 9692 7546 9720 8463
rect 9784 8362 9812 9318
rect 10152 9178 10180 9522
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10244 9110 10272 10474
rect 10336 10266 10364 10474
rect 10704 10470 10732 11154
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10520 9722 10548 9998
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10612 8838 10640 10134
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8634 10640 8774
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9784 7750 9812 8298
rect 10704 7936 10732 10406
rect 10796 9178 10824 11562
rect 10980 10996 11008 11698
rect 11348 11558 11376 12242
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10980 10968 11100 10996
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10980 9636 11008 10202
rect 11072 9738 11100 10968
rect 11164 10538 11192 11018
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11164 10062 11192 10474
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9897 11192 9998
rect 11150 9888 11206 9897
rect 11150 9823 11206 9832
rect 11072 9710 11192 9738
rect 11060 9648 11112 9654
rect 10980 9608 11060 9636
rect 11060 9590 11112 9596
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10796 8498 10824 9114
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10782 8392 10838 8401
rect 10782 8327 10838 8336
rect 10796 8090 10824 8327
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10980 7954 11008 8191
rect 11058 7984 11114 7993
rect 10784 7948 10836 7954
rect 10704 7908 10784 7936
rect 10784 7890 10836 7896
rect 10968 7948 11020 7954
rect 11164 7954 11192 9710
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 11256 8362 11284 9046
rect 11244 8356 11296 8362
rect 11244 8298 11296 8304
rect 11348 7993 11376 11494
rect 11440 10198 11468 12038
rect 12452 11529 12480 15520
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 15474 11656 15530 11665
rect 15474 11591 15530 11600
rect 12438 11520 12494 11529
rect 12438 11455 12494 11464
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10674 11560 11086
rect 11624 10810 11652 11222
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13174 11112 13230 11121
rect 13174 11047 13176 11056
rect 13228 11047 13230 11056
rect 13176 11018 13228 11024
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11624 10266 11652 10746
rect 12728 10606 12756 10950
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11440 9722 11468 10134
rect 11624 9722 11652 10202
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11612 9716 11664 9722
rect 11612 9658 11664 9664
rect 11624 9178 11652 9658
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 12360 9042 12388 10406
rect 12624 9648 12676 9654
rect 12530 9616 12586 9625
rect 12624 9590 12676 9596
rect 12530 9551 12532 9560
rect 12584 9551 12586 9560
rect 12532 9522 12584 9528
rect 12544 9178 12572 9522
rect 12636 9450 12664 9590
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 8634 12388 8978
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 11334 7984 11390 7993
rect 11058 7919 11114 7928
rect 11152 7948 11204 7954
rect 10968 7890 11020 7896
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9784 6934 9812 7686
rect 9968 7478 9996 7822
rect 10796 7546 10824 7890
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 9956 7472 10008 7478
rect 9954 7440 9956 7449
rect 10008 7440 10010 7449
rect 9954 7375 10010 7384
rect 10244 7274 10272 7482
rect 11072 7449 11100 7919
rect 11334 7919 11390 7928
rect 11152 7890 11204 7896
rect 11058 7440 11114 7449
rect 10968 7404 11020 7410
rect 11058 7375 11114 7384
rect 10968 7346 11020 7352
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10506 7032 10562 7041
rect 10612 7002 10640 7142
rect 10506 6967 10562 6976
rect 10600 6996 10652 7002
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9784 6118 9812 6870
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10244 6118 10272 6734
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 9586 5944 9642 5953
rect 9586 5879 9588 5888
rect 9640 5879 9642 5888
rect 9588 5850 9640 5856
rect 9784 5846 9812 6054
rect 9496 5840 9548 5846
rect 9772 5840 9824 5846
rect 9586 5808 9642 5817
rect 9548 5788 9586 5794
rect 9496 5782 9586 5788
rect 9508 5766 9586 5782
rect 9772 5782 9824 5788
rect 9586 5743 9642 5752
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9588 4480 9640 4486
rect 9692 4468 9720 5646
rect 9784 5370 9812 5782
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9784 5098 9812 5306
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9640 4440 9720 4468
rect 9588 4422 9640 4428
rect 9586 3904 9642 3913
rect 9586 3839 9642 3848
rect 9218 3768 9274 3777
rect 9218 3703 9220 3712
rect 9272 3703 9274 3712
rect 9220 3674 9272 3680
rect 8392 3606 8444 3612
rect 8850 3632 8906 3641
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8128 3194 8156 3334
rect 8116 3188 8168 3194
rect 8116 3130 8168 3136
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7840 2984 7892 2990
rect 7840 2926 7892 2932
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2514 7144 2790
rect 7852 2582 7880 2926
rect 8128 2650 8156 3130
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 7104 2508 7156 2514
rect 8220 2496 8248 3470
rect 8404 2922 8432 3606
rect 8850 3567 8906 3576
rect 9034 3632 9090 3641
rect 9034 3567 9090 3576
rect 9232 2990 9260 3674
rect 9600 3618 9628 3839
rect 9692 3738 9720 4440
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9600 3602 9720 3618
rect 9600 3596 9732 3602
rect 9600 3590 9680 3596
rect 9680 3538 9732 3544
rect 9692 3126 9720 3538
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 3058 9812 4694
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9876 3194 9904 4626
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9968 4078 9996 4490
rect 9956 4072 10008 4078
rect 9954 4040 9956 4049
rect 10008 4040 10010 4049
rect 9954 3975 10010 3984
rect 9968 3670 9996 3975
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8404 2650 8432 2858
rect 8850 2680 8906 2689
rect 8392 2644 8444 2650
rect 9600 2650 9628 2926
rect 10060 2650 10088 4966
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10152 4185 10180 4558
rect 10138 4176 10194 4185
rect 10138 4111 10194 4120
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 3738 10180 4014
rect 10244 3942 10272 6054
rect 10520 5545 10548 6967
rect 10600 6938 10652 6944
rect 10690 6488 10746 6497
rect 10690 6423 10746 6432
rect 10704 5817 10732 6423
rect 10980 6304 11008 7346
rect 11060 6316 11112 6322
rect 10980 6276 11060 6304
rect 11060 6258 11112 6264
rect 10874 6216 10930 6225
rect 10784 6180 10836 6186
rect 10874 6151 10876 6160
rect 10784 6122 10836 6128
rect 10928 6151 10930 6160
rect 10876 6122 10928 6128
rect 10690 5808 10746 5817
rect 10690 5743 10746 5752
rect 10506 5536 10562 5545
rect 10506 5471 10562 5480
rect 10704 4826 10732 5743
rect 10796 5658 10824 6122
rect 10874 5672 10930 5681
rect 10796 5630 10874 5658
rect 10874 5607 10876 5616
rect 10928 5607 10930 5616
rect 10876 5578 10928 5584
rect 11518 5536 11574 5545
rect 11518 5471 11574 5480
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10704 4078 10732 4762
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10888 3942 10916 4422
rect 10980 4146 11008 4626
rect 11532 4185 11560 5471
rect 11518 4176 11574 4185
rect 10968 4140 11020 4146
rect 11808 4146 11836 8191
rect 12728 7954 12756 10542
rect 13464 10470 13492 11154
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13096 10033 13124 10202
rect 13082 10024 13138 10033
rect 13082 9959 13138 9968
rect 13096 9654 13124 9959
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12820 8498 12848 8774
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12820 8401 12848 8434
rect 12806 8392 12862 8401
rect 12806 8327 12862 8336
rect 13464 8265 13492 10406
rect 14200 10130 14228 10542
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 14289 10288 14585 10308
rect 14188 10124 14240 10130
rect 14188 10066 14240 10072
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13726 9888 13782 9897
rect 13726 9823 13782 9832
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13450 8256 13506 8265
rect 13450 8191 13506 8200
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12176 7478 12204 7890
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12636 7546 12664 7754
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12624 7336 12676 7342
rect 12622 7304 12624 7313
rect 12676 7304 12678 7313
rect 12622 7239 12678 7248
rect 12728 7177 12756 7890
rect 13556 7478 13584 9454
rect 13740 8974 13768 9823
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8090 13768 8910
rect 13832 8634 13860 9046
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13818 7984 13874 7993
rect 13740 7928 13818 7936
rect 13740 7908 13820 7928
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 12808 7200 12860 7206
rect 12714 7168 12770 7177
rect 12808 7142 12860 7148
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12714 7103 12770 7112
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 5914 12020 6734
rect 12084 6458 12112 6802
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12084 6186 12112 6394
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11888 5704 11940 5710
rect 12176 5681 12204 5782
rect 11888 5646 11940 5652
rect 12162 5672 12218 5681
rect 11900 4486 11928 5646
rect 12162 5607 12218 5616
rect 12176 5370 12204 5607
rect 12254 5536 12310 5545
rect 12360 5522 12388 5850
rect 12820 5846 12848 7142
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 6225 12940 6598
rect 12992 6248 13044 6254
rect 12898 6216 12954 6225
rect 12992 6190 13044 6196
rect 12898 6151 12954 6160
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12360 5494 12480 5522
rect 12254 5471 12310 5480
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 12162 5264 12218 5273
rect 12162 5199 12218 5208
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11518 4111 11574 4120
rect 11796 4140 11848 4146
rect 10968 4082 11020 4088
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10152 3505 10180 3674
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10138 3496 10194 3505
rect 10138 3431 10194 3440
rect 10336 3194 10364 3538
rect 10324 3188 10376 3194
rect 10244 3148 10324 3176
rect 8850 2615 8852 2624
rect 8392 2586 8444 2592
rect 8904 2615 8906 2624
rect 9588 2644 9640 2650
rect 8852 2586 8904 2592
rect 9588 2586 9640 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10244 2514 10272 3148
rect 10324 3130 10376 3136
rect 11532 2514 11560 4111
rect 11796 4082 11848 4088
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 8300 2508 8352 2514
rect 8220 2468 8300 2496
rect 7104 2450 7156 2456
rect 8300 2450 8352 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 8300 2372 8352 2378
rect 8300 2314 8352 2320
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 8312 480 8340 2314
rect 11624 480 11652 3878
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 11808 3126 11836 3538
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11900 2650 11928 4422
rect 12176 3777 12204 5199
rect 12268 4690 12296 5471
rect 12452 4826 12480 5494
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12622 4720 12678 4729
rect 12256 4684 12308 4690
rect 12622 4655 12624 4664
rect 12256 4626 12308 4632
rect 12676 4655 12678 4664
rect 12624 4626 12676 4632
rect 12268 4282 12296 4626
rect 12440 4480 12492 4486
rect 12360 4428 12440 4434
rect 12360 4422 12492 4428
rect 12360 4406 12480 4422
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12162 3768 12218 3777
rect 12162 3703 12218 3712
rect 12176 3126 12204 3703
rect 12256 3664 12308 3670
rect 12254 3632 12256 3641
rect 12308 3632 12310 3641
rect 12254 3567 12310 3576
rect 12360 3194 12388 4406
rect 12636 3738 12664 4626
rect 13004 4146 13032 6190
rect 13096 5273 13124 7142
rect 13176 6180 13228 6186
rect 13176 6122 13228 6128
rect 13188 5914 13216 6122
rect 13176 5908 13228 5914
rect 13176 5850 13228 5856
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13082 5264 13138 5273
rect 13082 5199 13138 5208
rect 13176 5092 13228 5098
rect 13176 5034 13228 5040
rect 13188 4486 13216 5034
rect 13464 4826 13492 5782
rect 13556 4865 13584 7414
rect 13648 7274 13676 7686
rect 13740 7546 13768 7908
rect 13872 7919 13874 7928
rect 13820 7890 13872 7896
rect 13818 7848 13874 7857
rect 13818 7783 13874 7792
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13832 7410 13860 7783
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13648 6236 13676 7210
rect 13740 6458 13768 7210
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13648 6208 13768 6236
rect 13924 6225 13952 9318
rect 14108 8945 14136 9998
rect 14200 9722 14228 10066
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14094 8936 14150 8945
rect 14094 8871 14150 8880
rect 14108 8838 14136 8871
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 7750 14044 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7002 14044 7686
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6458 14044 6598
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13740 5642 13768 6208
rect 13910 6216 13966 6225
rect 13910 6151 13966 6160
rect 13924 5914 13952 6151
rect 14108 6100 14136 8774
rect 14200 6730 14228 9658
rect 14384 9586 14412 9998
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 14660 8022 14688 8366
rect 14738 8256 14794 8265
rect 14738 8191 14794 8200
rect 14752 8090 14780 8191
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14648 8016 14700 8022
rect 14648 7958 14700 7964
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14568 7546 14596 7822
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14844 6798 14872 10406
rect 14936 9110 14964 10610
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 15120 10266 15148 10474
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15212 9654 15240 10474
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9178 15056 9522
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 15290 7576 15346 7585
rect 15290 7511 15292 7520
rect 15344 7511 15346 7520
rect 15292 7482 15344 7488
rect 14924 7200 14976 7206
rect 14924 7142 14976 7148
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14188 6724 14240 6730
rect 14188 6666 14240 6672
rect 14936 6497 14964 7142
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14922 6488 14978 6497
rect 14922 6423 14978 6432
rect 14186 6352 14242 6361
rect 14186 6287 14242 6296
rect 14200 6254 14228 6287
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 15028 6118 15056 6802
rect 15384 6248 15436 6254
rect 15198 6216 15254 6225
rect 15384 6190 15436 6196
rect 15198 6151 15254 6160
rect 14188 6112 14240 6118
rect 14108 6072 14188 6100
rect 14188 6054 14240 6060
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13740 5302 13768 5578
rect 14108 5409 14136 5782
rect 14200 5545 14228 6054
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14924 5704 14976 5710
rect 14830 5672 14886 5681
rect 14924 5646 14976 5652
rect 14830 5607 14886 5616
rect 14740 5568 14792 5574
rect 14186 5536 14242 5545
rect 14740 5510 14792 5516
rect 14186 5471 14242 5480
rect 14094 5400 14150 5409
rect 14094 5335 14096 5344
rect 14148 5335 14150 5344
rect 14096 5306 14148 5312
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 14752 5234 14780 5510
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 13832 5114 13860 5170
rect 13648 5086 13860 5114
rect 14844 5098 14872 5607
rect 14936 5234 14964 5646
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 5092 14884 5098
rect 13542 4856 13598 4865
rect 13452 4820 13504 4826
rect 13542 4791 13598 4800
rect 13452 4762 13504 4768
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12728 3602 12756 4014
rect 12716 3596 12768 3602
rect 12716 3538 12768 3544
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 3194 13216 3470
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 11980 3120 12032 3126
rect 11980 3062 12032 3068
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11992 1873 12020 3062
rect 13648 2650 13676 5086
rect 14832 5034 14884 5040
rect 13728 5024 13780 5030
rect 14738 4992 14794 5001
rect 13780 4972 13860 4978
rect 13728 4966 13860 4972
rect 13740 4950 13860 4966
rect 13832 4758 13860 4950
rect 14289 4924 14585 4944
rect 14738 4927 14794 4936
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 3942 13768 4558
rect 13832 4282 13860 4694
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 3194 14044 3878
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14384 3505 14412 3538
rect 14648 3528 14700 3534
rect 14370 3496 14426 3505
rect 14648 3470 14700 3476
rect 14370 3431 14426 3440
rect 14004 3188 14056 3194
rect 14004 3130 14056 3136
rect 14384 3126 14412 3431
rect 14372 3120 14424 3126
rect 14186 3088 14242 3097
rect 14372 3062 14424 3068
rect 14186 3023 14188 3032
rect 14240 3023 14242 3032
rect 14188 2994 14240 3000
rect 14660 2961 14688 3470
rect 14646 2952 14702 2961
rect 14646 2887 14702 2896
rect 14289 2748 14585 2768
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 14660 2582 14688 2887
rect 14648 2576 14700 2582
rect 13358 2544 13414 2553
rect 12900 2508 12952 2514
rect 14648 2518 14700 2524
rect 14752 2514 14780 4927
rect 14844 4826 14872 5034
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14936 4758 14964 5170
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15028 4457 15056 6054
rect 15212 5710 15240 6151
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15396 5574 15424 6190
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 15014 4448 15070 4457
rect 15014 4383 15070 4392
rect 15120 4146 15148 5034
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 2922 14872 3606
rect 14936 3194 14964 4014
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15212 3398 15240 3878
rect 15304 3738 15332 4626
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 14936 2650 14964 3130
rect 15212 3058 15240 3334
rect 15488 3194 15516 11591
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15842 11520 15898 11529
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10266 15608 11154
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15672 10198 15700 11494
rect 15842 11455 15898 11464
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15672 9722 15700 10134
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15764 9042 15792 11290
rect 15752 9036 15804 9042
rect 15752 8978 15804 8984
rect 15764 8634 15792 8978
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15764 8022 15792 8230
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15764 7274 15792 7958
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15764 6186 15792 7210
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15580 4146 15608 4966
rect 15856 4690 15884 11455
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15948 9110 15976 9386
rect 15936 9104 15988 9110
rect 15936 9046 15988 9052
rect 15948 8294 15976 9046
rect 16040 8566 16068 10911
rect 16132 10538 16160 11086
rect 17512 10810 17540 15520
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 19432 12300 19484 12306
rect 19432 12242 19484 12248
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18604 11688 18656 11694
rect 18602 11656 18604 11665
rect 18656 11656 18658 11665
rect 18602 11591 18658 11600
rect 18234 11384 18290 11393
rect 19352 11370 19380 12038
rect 19444 11558 19472 12242
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 22480 11898 22508 15520
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 22468 11892 22520 11898
rect 22468 11834 22520 11840
rect 19524 11824 19576 11830
rect 19524 11766 19576 11772
rect 19432 11552 19484 11558
rect 19430 11520 19432 11529
rect 19484 11520 19486 11529
rect 19430 11455 19486 11464
rect 18234 11319 18290 11328
rect 19260 11342 19380 11370
rect 18248 11218 18276 11319
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10532 16172 10538
rect 16120 10474 16172 10480
rect 16224 10062 16252 10610
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16592 9654 16620 10134
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 16592 9178 16620 9590
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16960 8809 16988 9454
rect 16946 8800 17002 8809
rect 16946 8735 17002 8744
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 16040 8430 16068 8502
rect 16028 8424 16080 8430
rect 16026 8392 16028 8401
rect 16948 8424 17000 8430
rect 16080 8392 16082 8401
rect 16948 8366 17000 8372
rect 16026 8327 16082 8336
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 16670 7848 16726 7857
rect 16670 7783 16726 7792
rect 16580 7268 16632 7274
rect 16580 7210 16632 7216
rect 16592 7041 16620 7210
rect 16578 7032 16634 7041
rect 16578 6967 16634 6976
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16210 6488 16266 6497
rect 16316 6458 16344 6870
rect 16684 6866 16712 7783
rect 16960 7750 16988 8366
rect 17040 8356 17092 8362
rect 17040 8298 17092 8304
rect 17052 8090 17080 8298
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7290 16988 7686
rect 17052 7410 17080 8026
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16960 7262 17080 7290
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16578 6488 16634 6497
rect 16210 6423 16266 6432
rect 16304 6452 16356 6458
rect 16224 5166 16252 6423
rect 16578 6423 16580 6432
rect 16304 6394 16356 6400
rect 16632 6423 16634 6432
rect 16580 6394 16632 6400
rect 16684 6066 16712 6802
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 6458 16896 6734
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16684 6038 16804 6066
rect 16672 5908 16724 5914
rect 16672 5850 16724 5856
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16408 5234 16436 5782
rect 16488 5568 16540 5574
rect 16540 5528 16620 5556
rect 16488 5510 16540 5516
rect 16592 5234 16620 5528
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16684 4758 16712 5850
rect 16776 5710 16804 6038
rect 16960 5846 16988 6598
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 17052 4826 17080 7262
rect 17144 5166 17172 9590
rect 17408 9512 17460 9518
rect 17406 9480 17408 9489
rect 17460 9480 17462 9489
rect 17406 9415 17462 9424
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17328 8498 17356 9318
rect 17604 9178 17632 10066
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17604 8106 17632 9114
rect 17512 8078 17632 8106
rect 17512 6361 17540 8078
rect 17592 8016 17644 8022
rect 17592 7958 17644 7964
rect 17604 7546 17632 7958
rect 17696 7585 17724 10542
rect 17868 10124 17920 10130
rect 17868 10066 17920 10072
rect 17880 9654 17908 10066
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17866 9072 17922 9081
rect 17866 9007 17868 9016
rect 17920 9007 17922 9016
rect 17868 8978 17920 8984
rect 17880 8634 17908 8978
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17972 7886 18000 11018
rect 18248 10470 18276 11154
rect 18786 10704 18842 10713
rect 18786 10639 18842 10648
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 9761 18276 10406
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18234 9752 18290 9761
rect 18234 9687 18290 9696
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 8095 18092 8230
rect 18050 8086 18106 8095
rect 18050 8021 18106 8030
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17682 7576 17738 7585
rect 17592 7540 17644 7546
rect 17682 7511 17738 7520
rect 17592 7482 17644 7488
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17040 4820 17092 4826
rect 17040 4762 17092 4768
rect 17512 4758 17540 6287
rect 17696 5953 17724 7511
rect 17972 7002 18000 7822
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17788 6458 17816 6802
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17682 5944 17738 5953
rect 17788 5914 17816 6394
rect 17866 6216 17922 6225
rect 17866 6151 17922 6160
rect 17682 5879 17738 5888
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17788 5370 17816 5850
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17776 5024 17828 5030
rect 17774 4992 17776 5001
rect 17828 4992 17830 5001
rect 17774 4927 17830 4936
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 17500 4752 17552 4758
rect 17552 4700 17632 4706
rect 17500 4694 17632 4700
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16316 4010 16344 4626
rect 16408 4078 16436 4694
rect 17512 4678 17632 4694
rect 17132 4616 17184 4622
rect 17130 4584 17132 4593
rect 17184 4584 17186 4593
rect 17130 4519 17186 4528
rect 16672 4480 16724 4486
rect 16948 4480 17000 4486
rect 16724 4440 16804 4468
rect 16672 4422 16724 4428
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16304 4004 16356 4010
rect 16304 3946 16356 3952
rect 15842 3768 15898 3777
rect 15842 3703 15844 3712
rect 15896 3703 15898 3712
rect 15844 3674 15896 3680
rect 16316 3602 16344 3946
rect 16500 3738 16528 4014
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 16316 2990 16344 3538
rect 16592 3466 16620 4150
rect 16776 4146 16804 4440
rect 16948 4422 17000 4428
rect 17038 4448 17094 4457
rect 16960 4282 16988 4422
rect 17038 4383 17094 4392
rect 16948 4276 17000 4282
rect 16948 4218 17000 4224
rect 17052 4146 17080 4383
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 16776 3942 16804 4082
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16592 3126 16620 3402
rect 16776 3194 16804 3878
rect 17604 3738 17632 4678
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17788 3534 17816 3946
rect 17880 3738 17908 6151
rect 18156 5574 18184 6734
rect 18340 5778 18368 9998
rect 18800 9994 18828 10639
rect 19156 10532 19208 10538
rect 19156 10474 19208 10480
rect 18878 10432 18934 10441
rect 18878 10367 18934 10376
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18800 9722 18828 9930
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18800 9518 18828 9658
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18708 9178 18736 9318
rect 18696 9172 18748 9178
rect 18696 9114 18748 9120
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 8362 18460 8774
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18420 8356 18472 8362
rect 18420 8298 18472 8304
rect 18432 7750 18460 8298
rect 18524 8090 18552 8434
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7886 18644 8434
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18708 7954 18736 8298
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18616 7290 18644 7822
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18800 7478 18828 7511
rect 18788 7472 18840 7478
rect 18788 7414 18840 7420
rect 18616 7262 18736 7290
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18420 6724 18472 6730
rect 18420 6666 18472 6672
rect 18432 6118 18460 6666
rect 18524 6322 18552 6802
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18616 6186 18644 7142
rect 18708 6769 18736 7262
rect 18694 6760 18750 6769
rect 18694 6695 18750 6704
rect 18708 6322 18736 6695
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18432 4865 18460 6054
rect 18616 5914 18644 6122
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18418 4856 18474 4865
rect 18418 4791 18474 4800
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 18064 4282 18092 4422
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18064 4128 18092 4218
rect 18144 4140 18196 4146
rect 18064 4100 18144 4128
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 3194 17816 3470
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 15016 2984 15068 2990
rect 15016 2926 15068 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 13358 2479 13360 2488
rect 12900 2450 12952 2456
rect 13412 2479 13414 2488
rect 14740 2508 14792 2514
rect 13360 2450 13412 2456
rect 14740 2450 14792 2456
rect 12912 2009 12940 2450
rect 12898 2000 12954 2009
rect 12898 1935 12954 1944
rect 11978 1864 12034 1873
rect 11978 1799 12034 1808
rect 15028 480 15056 2926
rect 16316 2650 16344 2926
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16684 2446 16712 2926
rect 16776 2650 16804 3130
rect 17880 3058 17908 3674
rect 17972 3602 18000 4014
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17972 2650 18000 3402
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 15200 2440 15252 2446
rect 15198 2408 15200 2417
rect 16672 2440 16724 2446
rect 15252 2408 15254 2417
rect 16672 2382 16724 2388
rect 15198 2343 15254 2352
rect 18064 610 18092 4100
rect 18144 4082 18196 4088
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18340 2990 18368 3402
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18432 2854 18460 4791
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18524 3194 18552 3538
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 18708 2650 18736 4626
rect 18788 4004 18840 4010
rect 18788 3946 18840 3952
rect 18800 3097 18828 3946
rect 18892 3738 18920 10367
rect 19168 10266 19196 10474
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19168 9586 19196 10202
rect 19260 10062 19288 11342
rect 19536 11218 19564 11766
rect 20718 11656 20774 11665
rect 20718 11591 20774 11600
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19352 11121 19380 11154
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19352 10810 19380 11047
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19536 10470 19564 11154
rect 19720 10674 19748 11494
rect 20168 11008 20220 11014
rect 20168 10950 20220 10956
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19352 9382 19380 10066
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18984 8072 19012 8842
rect 19076 8362 19104 9046
rect 19168 8430 19196 9318
rect 19444 8634 19472 10202
rect 19536 10130 19564 10406
rect 20088 10266 20116 10610
rect 20180 10538 20208 10950
rect 20732 10849 20760 11591
rect 24136 11558 24164 12242
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24306 11792 24362 11801
rect 24306 11727 24362 11736
rect 24320 11694 24348 11727
rect 24308 11688 24360 11694
rect 24308 11630 24360 11636
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20718 10840 20774 10849
rect 20718 10775 20774 10784
rect 20168 10532 20220 10538
rect 20168 10474 20220 10480
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19812 8945 19840 9318
rect 19996 8974 20024 10066
rect 20180 9722 20208 10474
rect 20732 10146 20760 10775
rect 20824 10470 20852 11222
rect 21652 11150 21680 11494
rect 23386 11384 23442 11393
rect 23386 11319 23442 11328
rect 23400 11218 23428 11319
rect 24136 11257 24164 11494
rect 24412 11286 24440 12038
rect 24400 11280 24452 11286
rect 24122 11248 24178 11257
rect 23388 11212 23440 11218
rect 23440 11172 23520 11200
rect 24400 11222 24452 11228
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24122 11183 24178 11192
rect 23388 11154 23440 11160
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21640 11144 21692 11150
rect 21640 11086 21692 11092
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20640 10118 20760 10146
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20640 9058 20668 10118
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20732 9178 20760 9998
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20640 9042 20760 9058
rect 20640 9036 20772 9042
rect 20640 9030 20720 9036
rect 20720 8978 20772 8984
rect 19984 8968 20036 8974
rect 19798 8936 19854 8945
rect 19524 8900 19576 8906
rect 19798 8871 19854 8880
rect 19982 8936 19984 8945
rect 20036 8936 20038 8945
rect 19982 8871 20038 8880
rect 19524 8842 19576 8848
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 19432 8288 19484 8294
rect 19430 8256 19432 8265
rect 19484 8256 19486 8265
rect 19430 8191 19486 8200
rect 19064 8084 19116 8090
rect 18984 8044 19064 8072
rect 18984 7886 19012 8044
rect 19064 8026 19116 8032
rect 19156 8016 19208 8022
rect 19076 7964 19156 7970
rect 19076 7958 19208 7964
rect 19076 7942 19196 7958
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 19076 7818 19104 7942
rect 19536 7886 19564 8842
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19524 7880 19576 7886
rect 19430 7848 19486 7857
rect 19064 7812 19116 7818
rect 19524 7822 19576 7828
rect 19430 7783 19486 7792
rect 19064 7754 19116 7760
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19168 6866 19196 7346
rect 19260 7206 19288 7686
rect 19444 7585 19472 7783
rect 19430 7576 19486 7585
rect 19430 7511 19486 7520
rect 19536 7478 19564 7822
rect 19524 7472 19576 7478
rect 19524 7414 19576 7420
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19246 7032 19302 7041
rect 19246 6967 19302 6976
rect 19260 6866 19288 6967
rect 19628 6866 19656 8230
rect 20166 7440 20222 7449
rect 20166 7375 20222 7384
rect 20180 7342 20208 7375
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19156 6860 19208 6866
rect 19156 6802 19208 6808
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 4758 19012 6598
rect 19628 6186 19656 6802
rect 20168 6248 20220 6254
rect 20168 6190 20220 6196
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19628 5846 19656 6122
rect 19890 5944 19946 5953
rect 19812 5888 19890 5896
rect 19812 5868 19892 5888
rect 19616 5840 19668 5846
rect 19616 5782 19668 5788
rect 19248 5772 19300 5778
rect 19248 5714 19300 5720
rect 19064 5092 19116 5098
rect 19064 5034 19116 5040
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 19076 4690 19104 5034
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19064 4684 19116 4690
rect 19064 4626 19116 4632
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19168 3505 19196 4966
rect 19260 4826 19288 5714
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19352 4690 19380 5510
rect 19628 5370 19656 5782
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19812 5166 19840 5868
rect 19944 5879 19946 5888
rect 19892 5850 19944 5856
rect 20180 5574 20208 6190
rect 20168 5568 20220 5574
rect 20168 5510 20220 5516
rect 20180 5234 20208 5510
rect 20548 5370 20576 8298
rect 20732 7562 20760 8774
rect 20824 8634 20852 10406
rect 20996 10056 21048 10062
rect 20994 10024 20996 10033
rect 21048 10024 21050 10033
rect 20994 9959 21050 9968
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 21284 9586 21312 11018
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 21376 9897 21404 10746
rect 21468 10470 21496 11086
rect 21652 10674 21680 11086
rect 23204 11008 23256 11014
rect 21730 10976 21786 10985
rect 23204 10950 23256 10956
rect 21730 10911 21786 10920
rect 21744 10810 21772 10911
rect 23110 10840 23166 10849
rect 21732 10804 21784 10810
rect 23110 10775 23112 10784
rect 21732 10746 21784 10752
rect 23164 10775 23166 10784
rect 23112 10746 23164 10752
rect 21640 10668 21692 10674
rect 21640 10610 21692 10616
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21456 10464 21508 10470
rect 21560 10441 21588 10542
rect 21456 10406 21508 10412
rect 21546 10432 21602 10441
rect 21468 10305 21496 10406
rect 21546 10367 21602 10376
rect 21454 10296 21510 10305
rect 21454 10231 21510 10240
rect 21652 10130 21680 10610
rect 23124 10606 23152 10746
rect 22192 10600 22244 10606
rect 22192 10542 22244 10548
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21362 9888 21418 9897
rect 21362 9823 21418 9832
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 9178 21312 9522
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21272 9036 21324 9042
rect 21272 8978 21324 8984
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 21284 8566 21312 8978
rect 21376 8634 21404 9823
rect 21928 9722 21956 10134
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21272 8560 21324 8566
rect 21272 8502 21324 8508
rect 21376 8430 21404 8570
rect 21364 8424 21416 8430
rect 21270 8392 21326 8401
rect 21468 8401 21496 9318
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21560 8430 21588 8774
rect 21548 8424 21600 8430
rect 21364 8366 21416 8372
rect 21454 8392 21510 8401
rect 21270 8327 21326 8336
rect 21548 8366 21600 8372
rect 21454 8327 21510 8336
rect 20812 7744 20864 7750
rect 20810 7712 20812 7721
rect 20864 7712 20866 7721
rect 20810 7647 20866 7656
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20640 7546 20760 7562
rect 20628 7540 20760 7546
rect 20680 7534 20760 7540
rect 20628 7482 20680 7488
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20720 6792 20772 6798
rect 20718 6760 20720 6769
rect 20772 6760 20774 6769
rect 20718 6695 20774 6704
rect 20824 6458 20852 6802
rect 21284 6730 21312 8327
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21560 7410 21588 8230
rect 22008 8016 22060 8022
rect 22008 7958 22060 7964
rect 22020 7546 22048 7958
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 21272 6724 21324 6730
rect 21272 6666 21324 6672
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 21376 6186 21404 7210
rect 21560 6662 21588 7346
rect 22020 7002 22048 7482
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22112 6798 22140 7754
rect 22204 7342 22232 10542
rect 22928 10464 22980 10470
rect 22926 10432 22928 10441
rect 22980 10432 22982 10441
rect 22926 10367 22982 10376
rect 23216 10198 23244 10950
rect 23492 10452 23520 11172
rect 24412 10810 24440 11222
rect 24400 10804 24452 10810
rect 24400 10746 24452 10752
rect 23572 10464 23624 10470
rect 23492 10424 23572 10452
rect 23572 10406 23624 10412
rect 24400 10464 24452 10470
rect 24504 10452 24532 11222
rect 24596 10674 24624 12582
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24676 11552 24728 11558
rect 24676 11494 24728 11500
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24452 10424 24532 10452
rect 24400 10406 24452 10412
rect 23478 10296 23534 10305
rect 23478 10231 23534 10240
rect 23204 10192 23256 10198
rect 23204 10134 23256 10140
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 23216 9722 23244 10134
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23308 9654 23336 10134
rect 23492 10062 23520 10231
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9722 23520 9998
rect 23480 9716 23532 9722
rect 23480 9658 23532 9664
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23020 9512 23072 9518
rect 23020 9454 23072 9460
rect 23032 9110 23060 9454
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 22560 9036 22612 9042
rect 22560 8978 22612 8984
rect 22744 9036 22796 9042
rect 22744 8978 22796 8984
rect 22572 8362 22600 8978
rect 22756 8945 22784 8978
rect 22742 8936 22798 8945
rect 22742 8871 22798 8880
rect 22756 8634 22784 8871
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 22560 8356 22612 8362
rect 22560 8298 22612 8304
rect 22572 7750 22600 8298
rect 23492 8090 23520 8570
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22664 7206 22692 7890
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7313 23336 7686
rect 23400 7342 23428 7890
rect 23388 7336 23440 7342
rect 23294 7304 23350 7313
rect 23388 7278 23440 7284
rect 23294 7239 23350 7248
rect 22652 7200 22704 7206
rect 22652 7142 22704 7148
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 22100 6792 22152 6798
rect 22100 6734 22152 6740
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5846 20760 6054
rect 21652 5846 21680 6734
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21836 6458 21864 6666
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21836 6254 21864 6394
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 21640 5840 21692 5846
rect 21640 5782 21692 5788
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20548 5166 20576 5306
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19996 4729 20024 4762
rect 19982 4720 20038 4729
rect 19340 4684 19392 4690
rect 19982 4655 20038 4664
rect 19340 4626 19392 4632
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19904 4282 19932 4422
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 19248 4072 19300 4078
rect 19248 4014 19300 4020
rect 19154 3496 19210 3505
rect 19154 3431 19210 3440
rect 18786 3088 18842 3097
rect 18786 3023 18842 3032
rect 19168 2854 19196 3431
rect 19156 2848 19208 2854
rect 19154 2816 19156 2825
rect 19208 2816 19210 2825
rect 19154 2751 19210 2760
rect 19260 2650 19288 4014
rect 19890 3904 19946 3913
rect 19890 3839 19946 3848
rect 19904 3670 19932 3839
rect 19892 3664 19944 3670
rect 19892 3606 19944 3612
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19352 3194 19380 3538
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19352 2961 19380 3130
rect 19338 2952 19394 2961
rect 19338 2887 19394 2896
rect 19536 2825 19564 3538
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 19522 2816 19578 2825
rect 19522 2751 19578 2760
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 20272 2553 20300 2926
rect 20640 2582 20668 5034
rect 20732 4826 20760 5782
rect 22296 5710 22324 6054
rect 22572 5914 22600 6190
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 20824 5370 20852 5646
rect 21732 5568 21784 5574
rect 21732 5510 21784 5516
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 20824 4826 20852 5306
rect 21270 5264 21326 5273
rect 21270 5199 21326 5208
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20812 4820 20864 4826
rect 20812 4762 20864 4768
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20720 4004 20772 4010
rect 20720 3946 20772 3952
rect 20732 3738 20760 3946
rect 20916 3777 20944 4014
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 20902 3768 20958 3777
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20812 3732 20864 3738
rect 20902 3703 20958 3712
rect 20812 3674 20864 3680
rect 20732 3534 20760 3674
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20824 2990 20852 3674
rect 20916 3602 20944 3703
rect 21100 3641 21128 3878
rect 21086 3632 21142 3641
rect 20904 3596 20956 3602
rect 21086 3567 21142 3576
rect 20904 3538 20956 3544
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 20628 2576 20680 2582
rect 20258 2544 20314 2553
rect 20628 2518 20680 2524
rect 20258 2479 20314 2488
rect 20272 2378 20300 2479
rect 21008 2394 21036 2790
rect 21100 2582 21128 2858
rect 21088 2576 21140 2582
rect 21088 2518 21140 2524
rect 21284 2514 21312 5199
rect 21744 5166 21772 5510
rect 22296 5370 22324 5646
rect 22284 5364 22336 5370
rect 22284 5306 22336 5312
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21652 3942 21680 4014
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21744 3194 21772 5102
rect 22572 5098 22600 5850
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22296 4078 22324 4422
rect 22284 4072 22336 4078
rect 22284 4014 22336 4020
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 21744 2990 21772 3130
rect 21732 2984 21784 2990
rect 21732 2926 21784 2932
rect 21836 2922 21864 3538
rect 22020 2990 22048 3878
rect 22296 3534 22324 4014
rect 22664 3942 22692 7142
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23124 5953 23152 6394
rect 23110 5944 23166 5953
rect 23110 5879 23166 5888
rect 23308 5166 23336 7239
rect 23400 6882 23428 7278
rect 23400 6854 23520 6882
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23400 6497 23428 6598
rect 23386 6488 23442 6497
rect 23386 6423 23442 6432
rect 23492 6225 23520 6854
rect 23478 6216 23534 6225
rect 23478 6151 23534 6160
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23400 5846 23428 6054
rect 23388 5840 23440 5846
rect 23388 5782 23440 5788
rect 23296 5160 23348 5166
rect 23296 5102 23348 5108
rect 22742 4856 22798 4865
rect 23308 4826 23336 5102
rect 23400 5030 23428 5782
rect 23492 5370 23520 6151
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 22742 4791 22798 4800
rect 23296 4820 23348 4826
rect 22756 4690 22784 4791
rect 23296 4762 23348 4768
rect 22744 4684 22796 4690
rect 22744 4626 22796 4632
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22756 4570 22784 4626
rect 22756 4542 22876 4570
rect 22848 4146 22876 4542
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 22664 3641 22692 3878
rect 22650 3632 22706 3641
rect 22848 3602 22876 4082
rect 22940 4078 22968 4626
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23216 4185 23244 4422
rect 23202 4176 23258 4185
rect 23202 4111 23258 4120
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 23400 4010 23428 4966
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 22650 3567 22706 3576
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22468 3392 22520 3398
rect 22468 3334 22520 3340
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 21638 2816 21694 2825
rect 21638 2751 21694 2760
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20824 2366 21036 2394
rect 21362 2408 21418 2417
rect 20824 1873 20852 2366
rect 21362 2343 21364 2352
rect 21416 2343 21418 2352
rect 21364 2314 21416 2320
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20810 1864 20866 1873
rect 20810 1799 20866 1808
rect 18052 604 18104 610
rect 18052 546 18104 552
rect 18328 604 18380 610
rect 18328 546 18380 552
rect 18340 480 18368 546
rect 21652 480 21680 2751
rect 22112 2650 22140 3130
rect 22480 3126 22508 3334
rect 23124 3194 23152 3538
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 22468 3120 22520 3126
rect 22468 3062 22520 3068
rect 22560 2984 22612 2990
rect 22558 2952 22560 2961
rect 22612 2952 22614 2961
rect 23124 2922 23152 3130
rect 23308 2990 23336 3878
rect 23492 3194 23520 5063
rect 23584 4457 23612 10406
rect 24124 9920 24176 9926
rect 24124 9862 24176 9868
rect 24136 9518 24164 9862
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 23664 9376 23716 9382
rect 24412 9353 24440 10406
rect 24596 10198 24624 10474
rect 24584 10192 24636 10198
rect 24584 10134 24636 10140
rect 24688 9586 24716 11494
rect 24768 10192 24820 10198
rect 24872 10180 24900 12038
rect 24964 10713 24992 12582
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25240 11558 25268 12242
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25412 11552 25464 11558
rect 25412 11494 25464 11500
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24950 10704 25006 10713
rect 24950 10639 25006 10648
rect 25056 10538 25084 11086
rect 25044 10532 25096 10538
rect 25044 10474 25096 10480
rect 24820 10152 24900 10180
rect 24768 10134 24820 10140
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 23664 9318 23716 9324
rect 24398 9344 24454 9353
rect 23676 9110 23704 9318
rect 24398 9279 24454 9288
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23676 8838 23704 9046
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23676 8294 23704 8774
rect 24412 8634 24440 9279
rect 24872 9178 24900 10152
rect 24952 10192 25004 10198
rect 24952 10134 25004 10140
rect 24964 9722 24992 10134
rect 25056 10062 25084 10474
rect 25044 10056 25096 10062
rect 25042 10024 25044 10033
rect 25096 10024 25098 10033
rect 25042 9959 25098 9968
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24964 9382 24992 9658
rect 24952 9376 25004 9382
rect 24952 9318 25004 9324
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24964 9042 24992 9318
rect 25136 9172 25188 9178
rect 25136 9114 25188 9120
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 25148 8974 25176 9114
rect 25240 9081 25268 11494
rect 25226 9072 25282 9081
rect 25226 9007 25282 9016
rect 25136 8968 25188 8974
rect 25136 8910 25188 8916
rect 25148 8634 25176 8910
rect 25424 8634 25452 11494
rect 27448 11354 27476 15520
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 29552 12232 29604 12238
rect 29552 12174 29604 12180
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 29564 11286 29592 12174
rect 29734 11792 29790 11801
rect 29734 11727 29790 11736
rect 29552 11280 29604 11286
rect 29552 11222 29604 11228
rect 27068 11212 27120 11218
rect 27068 11154 27120 11160
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 27080 10810 27108 11154
rect 27620 11008 27672 11014
rect 27618 10976 27620 10985
rect 27672 10976 27674 10985
rect 27674 10934 27752 10962
rect 27618 10911 27674 10920
rect 27068 10804 27120 10810
rect 27068 10746 27120 10752
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 25976 9897 26004 10542
rect 26160 10266 26188 10542
rect 26240 10464 26292 10470
rect 26240 10406 26292 10412
rect 26606 10432 26662 10441
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 25962 9888 26018 9897
rect 25962 9823 26018 9832
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25516 9110 25544 9522
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 24400 8628 24452 8634
rect 24400 8570 24452 8576
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 24216 8424 24268 8430
rect 24216 8366 24268 8372
rect 25778 8392 25834 8401
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 24124 8084 24176 8090
rect 24124 8026 24176 8032
rect 23938 7440 23994 7449
rect 23938 7375 23994 7384
rect 23952 7342 23980 7375
rect 24136 7342 24164 8026
rect 24228 7750 24256 8366
rect 25778 8327 25834 8336
rect 25872 8356 25924 8362
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 25226 8256 25282 8265
rect 24688 8022 24716 8230
rect 25226 8191 25282 8200
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24228 7410 24256 7686
rect 24216 7404 24268 7410
rect 24216 7346 24268 7352
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 23952 6934 23980 7278
rect 24688 7206 24716 7958
rect 25044 7880 25096 7886
rect 25044 7822 25096 7828
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24676 7200 24728 7206
rect 24676 7142 24728 7148
rect 23940 6928 23992 6934
rect 23940 6870 23992 6876
rect 24030 6896 24086 6905
rect 24030 6831 24032 6840
rect 24084 6831 24086 6840
rect 24032 6802 24084 6808
rect 24044 6458 24072 6802
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 24584 6384 24636 6390
rect 24582 6352 24584 6361
rect 24636 6352 24638 6361
rect 24582 6287 24638 6296
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23676 5914 23704 6190
rect 24688 6118 24716 7142
rect 24872 6866 24900 7754
rect 25056 7206 25084 7822
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25056 6934 25084 7142
rect 25044 6928 25096 6934
rect 25044 6870 25096 6876
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24952 6724 25004 6730
rect 24952 6666 25004 6672
rect 24964 6458 24992 6666
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24676 6112 24728 6118
rect 24676 6054 24728 6060
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23676 5030 23704 5850
rect 24860 5772 24912 5778
rect 24860 5714 24912 5720
rect 25136 5772 25188 5778
rect 25136 5714 25188 5720
rect 24122 5672 24178 5681
rect 24872 5658 24900 5714
rect 24122 5607 24124 5616
rect 24176 5607 24178 5616
rect 24780 5630 24900 5658
rect 24124 5578 24176 5584
rect 24780 5370 24808 5630
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 24032 5092 24084 5098
rect 24032 5034 24084 5040
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23570 4448 23626 4457
rect 23570 4383 23626 4392
rect 24044 4282 24072 5034
rect 24950 4992 25006 5001
rect 24950 4927 25006 4936
rect 24492 4480 24544 4486
rect 24492 4422 24544 4428
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 24504 4078 24532 4422
rect 23940 4072 23992 4078
rect 23940 4014 23992 4020
rect 24492 4072 24544 4078
rect 24492 4014 24544 4020
rect 23952 3738 23980 4014
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 23848 3596 23900 3602
rect 23848 3538 23900 3544
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 23860 3233 23888 3538
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 23846 3224 23902 3233
rect 23480 3188 23532 3194
rect 23846 3159 23902 3168
rect 23480 3130 23532 3136
rect 23860 3126 23888 3159
rect 23848 3120 23900 3126
rect 23848 3062 23900 3068
rect 24596 2990 24624 3334
rect 23296 2984 23348 2990
rect 23296 2926 23348 2932
rect 24584 2984 24636 2990
rect 24584 2926 24636 2932
rect 22558 2887 22614 2896
rect 23112 2916 23164 2922
rect 23112 2858 23164 2864
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23480 2848 23532 2854
rect 23400 2796 23480 2802
rect 23400 2790 23532 2796
rect 23400 2774 23520 2790
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 23400 2582 23428 2774
rect 23768 2650 23796 2858
rect 24872 2854 24900 3538
rect 24860 2848 24912 2854
rect 24860 2790 24912 2796
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23388 2576 23440 2582
rect 22466 2544 22522 2553
rect 23388 2518 23440 2524
rect 24766 2544 24822 2553
rect 22466 2479 22522 2488
rect 24766 2479 24822 2488
rect 22480 2446 22508 2479
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22480 2281 22508 2382
rect 24780 2378 24808 2479
rect 24768 2372 24820 2378
rect 24768 2314 24820 2320
rect 22466 2272 22522 2281
rect 22466 2207 22522 2216
rect 24964 480 24992 4927
rect 25148 4826 25176 5714
rect 25240 5370 25268 8191
rect 25320 6860 25372 6866
rect 25320 6802 25372 6808
rect 25332 6458 25360 6802
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25504 5704 25556 5710
rect 25504 5646 25556 5652
rect 25228 5364 25280 5370
rect 25228 5306 25280 5312
rect 25240 5166 25268 5306
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 25320 5092 25372 5098
rect 25320 5034 25372 5040
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 25148 4214 25176 4762
rect 25332 4690 25360 5034
rect 25320 4684 25372 4690
rect 25320 4626 25372 4632
rect 25136 4208 25188 4214
rect 25136 4150 25188 4156
rect 25516 4049 25544 5646
rect 25792 4622 25820 8327
rect 25872 8298 25924 8304
rect 26056 8356 26108 8362
rect 26056 8298 26108 8304
rect 25884 8090 25912 8298
rect 26068 8265 26096 8298
rect 26054 8256 26110 8265
rect 26054 8191 26110 8200
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 26160 7528 26188 10202
rect 26068 7500 26188 7528
rect 26068 6730 26096 7500
rect 26252 7426 26280 10406
rect 26606 10367 26662 10376
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 26528 9382 26556 10202
rect 26620 10198 26648 10367
rect 26608 10192 26660 10198
rect 26608 10134 26660 10140
rect 26516 9376 26568 9382
rect 26514 9344 26516 9353
rect 26568 9344 26570 9353
rect 26514 9279 26570 9288
rect 26330 9072 26386 9081
rect 26330 9007 26386 9016
rect 26516 9036 26568 9042
rect 26344 7585 26372 9007
rect 26516 8978 26568 8984
rect 26528 8566 26556 8978
rect 26620 8974 26648 10134
rect 26884 10056 26936 10062
rect 26884 9998 26936 10004
rect 26896 9722 26924 9998
rect 26884 9716 26936 9722
rect 26884 9658 26936 9664
rect 26976 9036 27028 9042
rect 26976 8978 27028 8984
rect 26608 8968 26660 8974
rect 26988 8945 27016 8978
rect 26608 8910 26660 8916
rect 26974 8936 27030 8945
rect 26974 8871 27030 8880
rect 26988 8634 27016 8871
rect 26976 8628 27028 8634
rect 26976 8570 27028 8576
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26528 8362 26556 8502
rect 27080 8498 27108 10746
rect 27724 10606 27752 10934
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27988 10600 28040 10606
rect 27988 10542 28040 10548
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 28000 10266 28028 10542
rect 28092 10470 28120 11154
rect 28908 11144 28960 11150
rect 28908 11086 28960 11092
rect 28356 10532 28408 10538
rect 28356 10474 28408 10480
rect 28080 10464 28132 10470
rect 28080 10406 28132 10412
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28000 9897 28028 10202
rect 27986 9888 28042 9897
rect 27986 9823 28042 9832
rect 28000 9654 28028 9823
rect 27988 9648 28040 9654
rect 27988 9590 28040 9596
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27724 8430 27752 8774
rect 28092 8566 28120 10406
rect 28172 9444 28224 9450
rect 28172 9386 28224 9392
rect 28080 8560 28132 8566
rect 28080 8502 28132 8508
rect 27712 8424 27764 8430
rect 27712 8366 27764 8372
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 26884 8016 26936 8022
rect 26884 7958 26936 7964
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26330 7576 26386 7585
rect 26330 7511 26386 7520
rect 26160 7410 26280 7426
rect 26148 7404 26280 7410
rect 26200 7398 26280 7404
rect 26148 7346 26200 7352
rect 26160 7002 26188 7346
rect 26148 6996 26200 7002
rect 26148 6938 26200 6944
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 25872 6248 25924 6254
rect 25872 6190 25924 6196
rect 25884 5574 25912 6190
rect 25872 5568 25924 5574
rect 25872 5510 25924 5516
rect 25884 5234 25912 5510
rect 26068 5370 26096 6666
rect 26240 6656 26292 6662
rect 26160 6604 26240 6610
rect 26160 6598 26292 6604
rect 26160 6582 26280 6598
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 25872 5228 25924 5234
rect 25872 5170 25924 5176
rect 26068 5166 26096 5306
rect 26056 5160 26108 5166
rect 26056 5102 26108 5108
rect 26160 4758 26188 6582
rect 26344 5914 26372 6734
rect 26528 6662 26556 7822
rect 26896 7546 26924 7958
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 27712 7744 27764 7750
rect 27712 7686 27764 7692
rect 26884 7540 26936 7546
rect 26884 7482 26936 7488
rect 26896 7274 26924 7482
rect 26884 7268 26936 7274
rect 26884 7210 26936 7216
rect 27448 6934 27476 7686
rect 27724 7410 27752 7686
rect 28092 7410 28120 8230
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28080 7404 28132 7410
rect 28080 7346 28132 7352
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 27436 6928 27488 6934
rect 27436 6870 27488 6876
rect 26516 6656 26568 6662
rect 26516 6598 26568 6604
rect 27342 6488 27398 6497
rect 27448 6458 27476 6870
rect 27342 6423 27398 6432
rect 27436 6452 27488 6458
rect 27158 6352 27214 6361
rect 27158 6287 27214 6296
rect 26332 5908 26384 5914
rect 26332 5850 26384 5856
rect 26344 5817 26372 5850
rect 27172 5846 27200 6287
rect 27160 5840 27212 5846
rect 26330 5808 26386 5817
rect 27160 5782 27212 5788
rect 26330 5743 26386 5752
rect 27068 5704 27120 5710
rect 26882 5672 26938 5681
rect 27068 5646 27120 5652
rect 26882 5607 26938 5616
rect 26896 5370 26924 5607
rect 27080 5545 27108 5646
rect 27066 5536 27122 5545
rect 27066 5471 27122 5480
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 27172 4826 27200 5782
rect 27252 5364 27304 5370
rect 27252 5306 27304 5312
rect 27264 5098 27292 5306
rect 27252 5092 27304 5098
rect 27252 5034 27304 5040
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 26148 4752 26200 4758
rect 27356 4729 27384 6423
rect 27436 6394 27488 6400
rect 28000 6322 28028 7346
rect 28092 6934 28120 7346
rect 28184 7041 28212 9386
rect 28368 9042 28396 10474
rect 28816 10192 28868 10198
rect 28920 10180 28948 11086
rect 29564 10810 29592 11222
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 29460 10736 29512 10742
rect 29460 10678 29512 10684
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 29000 10192 29052 10198
rect 28920 10152 29000 10180
rect 28816 10134 28868 10140
rect 29000 10134 29052 10140
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 28552 9586 28580 9998
rect 28828 9654 28856 10134
rect 28816 9648 28868 9654
rect 28816 9590 28868 9596
rect 29012 9586 29040 10134
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28552 9178 28580 9522
rect 29184 9444 29236 9450
rect 29184 9386 29236 9392
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 29196 9110 29224 9386
rect 29184 9104 29236 9110
rect 29184 9046 29236 9052
rect 28356 9036 28408 9042
rect 28356 8978 28408 8984
rect 28368 8634 28396 8978
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 29196 8514 29224 9046
rect 28920 8486 29224 8514
rect 28920 8362 28948 8486
rect 29000 8424 29052 8430
rect 29000 8366 29052 8372
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 29012 7954 29040 8366
rect 29196 8022 29224 8486
rect 29184 8016 29236 8022
rect 29184 7958 29236 7964
rect 29000 7948 29052 7954
rect 29000 7890 29052 7896
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 28736 7274 28764 7822
rect 28724 7268 28776 7274
rect 28724 7210 28776 7216
rect 28170 7032 28226 7041
rect 28170 6967 28226 6976
rect 28080 6928 28132 6934
rect 28080 6870 28132 6876
rect 28080 6384 28132 6390
rect 28080 6326 28132 6332
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 28000 5846 28028 6258
rect 27988 5840 28040 5846
rect 27988 5782 28040 5788
rect 28000 5234 28028 5782
rect 28092 5574 28120 6326
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 28184 5386 28212 6967
rect 28632 5840 28684 5846
rect 28092 5358 28212 5386
rect 28552 5800 28632 5828
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 26148 4694 26200 4700
rect 27342 4720 27398 4729
rect 27160 4684 27212 4690
rect 28092 4690 28120 5358
rect 28552 5030 28580 5800
rect 28632 5782 28684 5788
rect 28172 5024 28224 5030
rect 28172 4966 28224 4972
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 27342 4655 27398 4664
rect 28080 4684 28132 4690
rect 27160 4626 27212 4632
rect 28080 4626 28132 4632
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 25792 4282 25820 4558
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 26424 4140 26476 4146
rect 26424 4082 26476 4088
rect 25502 4040 25558 4049
rect 25044 4004 25096 4010
rect 26436 4010 26464 4082
rect 25502 3975 25558 3984
rect 26424 4004 26476 4010
rect 25044 3946 25096 3952
rect 26424 3946 26476 3952
rect 25056 3670 25084 3946
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 25044 3664 25096 3670
rect 25044 3606 25096 3612
rect 25056 2922 25084 3606
rect 26252 3398 26280 3878
rect 26422 3768 26478 3777
rect 26422 3703 26478 3712
rect 26436 3602 26464 3703
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 25228 3392 25280 3398
rect 25228 3334 25280 3340
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 25240 2650 25268 3334
rect 26252 2650 26280 3334
rect 26344 3058 26372 3334
rect 26436 3194 26464 3538
rect 26424 3188 26476 3194
rect 26424 3130 26476 3136
rect 26332 3052 26384 3058
rect 26332 2994 26384 3000
rect 26528 2922 26556 4558
rect 27172 4282 27200 4626
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 26976 4004 27028 4010
rect 26976 3946 27028 3952
rect 26988 3505 27016 3946
rect 27172 3942 27200 4218
rect 27986 4176 28042 4185
rect 28092 4146 28120 4626
rect 28184 4214 28212 4966
rect 28552 4826 28580 4966
rect 28540 4820 28592 4826
rect 28540 4762 28592 4768
rect 28736 4758 28764 7210
rect 28816 6928 28868 6934
rect 28816 6870 28868 6876
rect 28828 6458 28856 6870
rect 28908 6792 28960 6798
rect 29092 6792 29144 6798
rect 28960 6752 29040 6780
rect 28908 6734 28960 6740
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 28828 6186 28856 6394
rect 28816 6180 28868 6186
rect 28816 6122 28868 6128
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 28920 5234 28948 5646
rect 29012 5370 29040 6752
rect 29092 6734 29144 6740
rect 29104 6322 29132 6734
rect 29092 6316 29144 6322
rect 29092 6258 29144 6264
rect 29104 5817 29132 6258
rect 29184 6112 29236 6118
rect 29184 6054 29236 6060
rect 29090 5808 29146 5817
rect 29090 5743 29146 5752
rect 29104 5710 29132 5743
rect 29092 5704 29144 5710
rect 29196 5681 29224 6054
rect 29288 5778 29316 10610
rect 29472 10266 29500 10678
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 29368 6180 29420 6186
rect 29368 6122 29420 6128
rect 29276 5772 29328 5778
rect 29276 5714 29328 5720
rect 29092 5646 29144 5652
rect 29182 5672 29238 5681
rect 29380 5642 29408 6122
rect 29182 5607 29238 5616
rect 29368 5636 29420 5642
rect 29368 5578 29420 5584
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29000 5364 29052 5370
rect 29000 5306 29052 5312
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 29104 4826 29132 5510
rect 29748 5370 29776 11727
rect 30104 11688 30156 11694
rect 30010 11656 30066 11665
rect 30066 11636 30104 11642
rect 30066 11630 30156 11636
rect 30066 11614 30144 11630
rect 32036 11620 32088 11626
rect 30010 11591 30066 11600
rect 32036 11562 32088 11568
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 29920 11280 29972 11286
rect 29826 11248 29882 11257
rect 29920 11222 29972 11228
rect 29826 11183 29882 11192
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29748 5166 29776 5306
rect 29736 5160 29788 5166
rect 29736 5102 29788 5108
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 28724 4752 28776 4758
rect 28724 4694 28776 4700
rect 28264 4684 28316 4690
rect 28264 4626 28316 4632
rect 28276 4282 28304 4626
rect 28264 4276 28316 4282
rect 28264 4218 28316 4224
rect 28172 4208 28224 4214
rect 28172 4150 28224 4156
rect 27986 4111 28042 4120
rect 28080 4140 28132 4146
rect 27804 4072 27856 4078
rect 27802 4040 27804 4049
rect 27856 4040 27858 4049
rect 27802 3975 27858 3984
rect 27160 3936 27212 3942
rect 27066 3904 27122 3913
rect 27160 3878 27212 3884
rect 27066 3839 27122 3848
rect 26974 3496 27030 3505
rect 26974 3431 27030 3440
rect 26988 3058 27016 3431
rect 26976 3052 27028 3058
rect 26976 2994 27028 3000
rect 27080 2990 27108 3839
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 28000 3534 28028 4111
rect 28080 4082 28132 4088
rect 29840 4078 29868 11183
rect 29932 10742 29960 11222
rect 29920 10736 29972 10742
rect 29920 10678 29972 10684
rect 30104 10532 30156 10538
rect 30104 10474 30156 10480
rect 30116 9926 30144 10474
rect 30300 10282 30328 11494
rect 30470 11384 30526 11393
rect 31496 11354 31524 11494
rect 30470 11319 30526 11328
rect 31484 11348 31536 11354
rect 30484 11286 30512 11319
rect 31484 11290 31536 11296
rect 30472 11280 30524 11286
rect 30472 11222 30524 11228
rect 30484 10674 30512 11222
rect 31496 10742 31524 11290
rect 31760 11212 31812 11218
rect 31760 11154 31812 11160
rect 31666 11112 31722 11121
rect 31666 11047 31722 11056
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 30472 10668 30524 10674
rect 30472 10610 30524 10616
rect 30472 10532 30524 10538
rect 30472 10474 30524 10480
rect 31576 10532 31628 10538
rect 31576 10474 31628 10480
rect 30300 10266 30420 10282
rect 30300 10260 30432 10266
rect 30300 10254 30380 10260
rect 30380 10202 30432 10208
rect 30104 9920 30156 9926
rect 30104 9862 30156 9868
rect 30116 9178 30144 9862
rect 30392 9722 30420 10202
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 30484 9042 30512 10474
rect 31116 10464 31168 10470
rect 31116 10406 31168 10412
rect 30564 10192 30616 10198
rect 30564 10134 30616 10140
rect 30576 9654 30604 10134
rect 31128 10062 31156 10406
rect 31588 10266 31616 10474
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 31482 10160 31538 10169
rect 31482 10095 31538 10104
rect 31116 10056 31168 10062
rect 31114 10024 31116 10033
rect 31168 10024 31170 10033
rect 31114 9959 31170 9968
rect 31496 9654 31524 10095
rect 30564 9648 30616 9654
rect 31484 9648 31536 9654
rect 30564 9590 30616 9596
rect 30746 9616 30802 9625
rect 31484 9590 31536 9596
rect 30746 9551 30802 9560
rect 30760 9518 30788 9551
rect 30748 9512 30800 9518
rect 30748 9454 30800 9460
rect 30472 9036 30524 9042
rect 30472 8978 30524 8984
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30196 8832 30248 8838
rect 30196 8774 30248 8780
rect 30208 8362 30236 8774
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 30196 8356 30248 8362
rect 30196 8298 30248 8304
rect 30208 8090 30236 8298
rect 30196 8084 30248 8090
rect 30196 8026 30248 8032
rect 30104 7948 30156 7954
rect 30104 7890 30156 7896
rect 30116 7410 30144 7890
rect 30104 7404 30156 7410
rect 30104 7346 30156 7352
rect 30392 6866 30420 8434
rect 30484 8401 30512 8978
rect 30944 8498 30972 8978
rect 31680 8634 31708 11047
rect 31772 10470 31800 11154
rect 31760 10464 31812 10470
rect 31760 10406 31812 10412
rect 32048 9761 32076 11562
rect 32404 11212 32456 11218
rect 32404 11154 32456 11160
rect 32416 10674 32444 11154
rect 32508 11121 32536 15520
rect 36358 14648 36414 14657
rect 36358 14583 36414 14592
rect 35622 13832 35678 13841
rect 35622 13767 35678 13776
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 35636 12442 35664 13767
rect 35714 12880 35770 12889
rect 35714 12815 35770 12824
rect 35624 12436 35676 12442
rect 35624 12378 35676 12384
rect 34612 12300 34664 12306
rect 34612 12242 34664 12248
rect 35440 12300 35492 12306
rect 35440 12242 35492 12248
rect 34152 12096 34204 12102
rect 34152 12038 34204 12044
rect 33416 11824 33468 11830
rect 33416 11766 33468 11772
rect 32680 11144 32732 11150
rect 32494 11112 32550 11121
rect 32680 11086 32732 11092
rect 32494 11047 32550 11056
rect 32404 10668 32456 10674
rect 32404 10610 32456 10616
rect 32220 10532 32272 10538
rect 32220 10474 32272 10480
rect 32232 10062 32260 10474
rect 32416 10470 32444 10610
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32220 10056 32272 10062
rect 32220 9998 32272 10004
rect 32416 9926 32444 10406
rect 32692 10266 32720 11086
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 32864 10464 32916 10470
rect 32864 10406 32916 10412
rect 32680 10260 32732 10266
rect 32680 10202 32732 10208
rect 32404 9920 32456 9926
rect 32402 9888 32404 9897
rect 32456 9888 32458 9897
rect 32402 9823 32458 9832
rect 32034 9752 32090 9761
rect 32034 9687 32090 9696
rect 31668 8628 31720 8634
rect 31852 8628 31904 8634
rect 31668 8570 31720 8576
rect 31772 8588 31852 8616
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31576 8424 31628 8430
rect 30470 8392 30526 8401
rect 30470 8327 30526 8336
rect 31574 8392 31576 8401
rect 31628 8392 31630 8401
rect 31772 8378 31800 8588
rect 31852 8570 31904 8576
rect 31574 8327 31630 8336
rect 31680 8350 31800 8378
rect 30484 8090 30512 8327
rect 30656 8288 30708 8294
rect 30656 8230 30708 8236
rect 30668 8090 30696 8230
rect 30472 8084 30524 8090
rect 30472 8026 30524 8032
rect 30656 8084 30708 8090
rect 30656 8026 30708 8032
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30576 7857 30604 7890
rect 30562 7848 30618 7857
rect 30562 7783 30618 7792
rect 31024 7812 31076 7818
rect 31024 7754 31076 7760
rect 31036 7546 31064 7754
rect 31024 7540 31076 7546
rect 31024 7482 31076 7488
rect 31390 7440 31446 7449
rect 31390 7375 31446 7384
rect 30562 7304 30618 7313
rect 30562 7239 30618 7248
rect 30576 6866 30604 7239
rect 30380 6860 30432 6866
rect 30380 6802 30432 6808
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30576 6458 30604 6802
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 30838 6488 30894 6497
rect 30564 6452 30616 6458
rect 30838 6423 30894 6432
rect 30564 6394 30616 6400
rect 30852 5846 30880 6423
rect 31128 6322 31156 6734
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 31128 5914 31156 6258
rect 31404 6254 31432 7375
rect 31680 6882 31708 8350
rect 32048 7342 32076 9687
rect 32416 9042 32444 9823
rect 32692 9586 32720 10202
rect 32680 9580 32732 9586
rect 32680 9522 32732 9528
rect 32680 9444 32732 9450
rect 32680 9386 32732 9392
rect 32128 9036 32180 9042
rect 32128 8978 32180 8984
rect 32404 9036 32456 9042
rect 32404 8978 32456 8984
rect 32140 8634 32168 8978
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 32416 8090 32444 8978
rect 32692 8362 32720 9386
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 32784 8498 32812 9046
rect 32772 8492 32824 8498
rect 32772 8434 32824 8440
rect 32680 8356 32732 8362
rect 32680 8298 32732 8304
rect 32404 8084 32456 8090
rect 32404 8026 32456 8032
rect 32692 7410 32720 8298
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32784 7546 32812 7890
rect 32772 7540 32824 7546
rect 32772 7482 32824 7488
rect 32680 7404 32732 7410
rect 32680 7346 32732 7352
rect 32036 7336 32088 7342
rect 32036 7278 32088 7284
rect 32692 6934 32720 7346
rect 31588 6866 31708 6882
rect 32680 6928 32732 6934
rect 32680 6870 32732 6876
rect 31576 6860 31708 6866
rect 31628 6854 31708 6860
rect 31576 6802 31628 6808
rect 32218 6760 32274 6769
rect 32218 6695 32274 6704
rect 31392 6248 31444 6254
rect 31392 6190 31444 6196
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 30840 5840 30892 5846
rect 30840 5782 30892 5788
rect 32232 5778 32260 6695
rect 32692 6458 32720 6870
rect 32680 6452 32732 6458
rect 32680 6394 32732 6400
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 32692 5914 32720 6190
rect 32680 5908 32732 5914
rect 32680 5850 32732 5856
rect 30104 5772 30156 5778
rect 30104 5714 30156 5720
rect 30380 5772 30432 5778
rect 30380 5714 30432 5720
rect 32220 5772 32272 5778
rect 32220 5714 32272 5720
rect 30116 5370 30144 5714
rect 30392 5658 30420 5714
rect 30300 5630 30420 5658
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 30300 4826 30328 5630
rect 30378 5536 30434 5545
rect 30378 5471 30434 5480
rect 30392 5370 30420 5471
rect 32232 5370 32260 5714
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 32220 5364 32272 5370
rect 32220 5306 32272 5312
rect 31298 5264 31354 5273
rect 31298 5199 31354 5208
rect 31312 5166 31340 5199
rect 31300 5160 31352 5166
rect 32232 5137 32260 5306
rect 32784 5302 32812 7482
rect 32876 7449 32904 10406
rect 33140 10192 33192 10198
rect 33140 10134 33192 10140
rect 33152 9722 33180 10134
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 33048 9512 33100 9518
rect 33244 9500 33272 10746
rect 33100 9472 33272 9500
rect 33048 9454 33100 9460
rect 33140 7744 33192 7750
rect 33140 7686 33192 7692
rect 32862 7440 32918 7449
rect 33152 7410 33180 7686
rect 32862 7375 32918 7384
rect 33140 7404 33192 7410
rect 33140 7346 33192 7352
rect 33152 7002 33180 7346
rect 33232 7200 33284 7206
rect 33230 7168 33232 7177
rect 33284 7168 33286 7177
rect 33230 7103 33286 7112
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 33048 6656 33100 6662
rect 33048 6598 33100 6604
rect 33060 6390 33088 6598
rect 33048 6384 33100 6390
rect 33048 6326 33100 6332
rect 33428 6225 33456 11766
rect 33876 11688 33928 11694
rect 33876 11630 33928 11636
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 33690 11384 33746 11393
rect 33690 11319 33746 11328
rect 33508 11280 33560 11286
rect 33508 11222 33560 11228
rect 33520 10849 33548 11222
rect 33506 10840 33562 10849
rect 33506 10775 33562 10784
rect 33704 10198 33732 11319
rect 33692 10192 33744 10198
rect 33692 10134 33744 10140
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 33520 6662 33548 7822
rect 33600 7812 33652 7818
rect 33600 7754 33652 7760
rect 33612 7274 33640 7754
rect 33600 7268 33652 7274
rect 33600 7210 33652 7216
rect 33796 6905 33824 11494
rect 33888 8514 33916 11630
rect 34060 11552 34112 11558
rect 34060 11494 34112 11500
rect 33968 11212 34020 11218
rect 33968 11154 34020 11160
rect 33980 10810 34008 11154
rect 34072 11121 34100 11494
rect 34058 11112 34114 11121
rect 34058 11047 34114 11056
rect 34058 10976 34114 10985
rect 34058 10911 34114 10920
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 34072 10742 34100 10911
rect 34060 10736 34112 10742
rect 34060 10678 34112 10684
rect 34060 10532 34112 10538
rect 34060 10474 34112 10480
rect 34072 8974 34100 10474
rect 34164 9586 34192 12038
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 34624 11626 34652 12242
rect 35452 11898 35480 12242
rect 35622 12064 35678 12073
rect 35622 11999 35678 12008
rect 35440 11892 35492 11898
rect 35440 11834 35492 11840
rect 35438 11792 35494 11801
rect 35438 11727 35494 11736
rect 35348 11688 35400 11694
rect 35348 11630 35400 11636
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 35072 11144 35124 11150
rect 35072 11086 35124 11092
rect 34796 11008 34848 11014
rect 34796 10950 34848 10956
rect 34980 11008 35032 11014
rect 34980 10950 35032 10956
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 34610 10432 34666 10441
rect 34610 10367 34666 10376
rect 34624 10062 34652 10367
rect 34808 10305 34836 10950
rect 34992 10538 35020 10950
rect 35084 10538 35112 11086
rect 34980 10532 35032 10538
rect 34980 10474 35032 10480
rect 35072 10532 35124 10538
rect 35072 10474 35124 10480
rect 34794 10296 34850 10305
rect 34794 10231 34850 10240
rect 34704 10192 34756 10198
rect 34992 10169 35020 10474
rect 34704 10134 34756 10140
rect 34978 10160 35034 10169
rect 34612 10056 34664 10062
rect 34612 9998 34664 10004
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 34624 9722 34652 9998
rect 34612 9716 34664 9722
rect 34612 9658 34664 9664
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 34336 9376 34388 9382
rect 34336 9318 34388 9324
rect 34152 9104 34204 9110
rect 34152 9046 34204 9052
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 34164 8634 34192 9046
rect 34348 9042 34376 9318
rect 34716 9042 34744 10134
rect 34978 10095 35034 10104
rect 34888 10056 34940 10062
rect 34886 10024 34888 10033
rect 34940 10024 34942 10033
rect 34886 9959 34942 9968
rect 34900 9654 34928 9959
rect 34888 9648 34940 9654
rect 34888 9590 34940 9596
rect 35084 9450 35112 10474
rect 35164 9580 35216 9586
rect 35164 9522 35216 9528
rect 35072 9444 35124 9450
rect 35072 9386 35124 9392
rect 35176 9178 35204 9522
rect 35164 9172 35216 9178
rect 35164 9114 35216 9120
rect 34336 9036 34388 9042
rect 34336 8978 34388 8984
rect 34704 9036 34756 9042
rect 34704 8978 34756 8984
rect 34704 8832 34756 8838
rect 34704 8774 34756 8780
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 33966 8528 34022 8537
rect 33888 8486 33966 8514
rect 33966 8463 34022 8472
rect 33782 6896 33838 6905
rect 33782 6831 33838 6840
rect 33876 6792 33928 6798
rect 33876 6734 33928 6740
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 33520 6497 33548 6598
rect 33506 6488 33562 6497
rect 33888 6458 33916 6734
rect 33506 6423 33562 6432
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 33414 6216 33470 6225
rect 33414 6151 33470 6160
rect 33428 5778 33456 6151
rect 33416 5772 33468 5778
rect 33416 5714 33468 5720
rect 33428 5370 33456 5714
rect 33416 5364 33468 5370
rect 33416 5306 33468 5312
rect 32772 5296 32824 5302
rect 32772 5238 32824 5244
rect 31300 5102 31352 5108
rect 32218 5128 32274 5137
rect 32218 5063 32274 5072
rect 31760 5024 31812 5030
rect 31758 4992 31760 5001
rect 31812 4992 31814 5001
rect 31758 4927 31814 4936
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 31574 4720 31630 4729
rect 30196 4684 30248 4690
rect 31574 4655 31630 4664
rect 30196 4626 30248 4632
rect 30208 4321 30236 4626
rect 30194 4312 30250 4321
rect 30194 4247 30196 4256
rect 30248 4247 30250 4256
rect 30196 4218 30248 4224
rect 30208 4187 30236 4218
rect 29828 4072 29880 4078
rect 29826 4040 29828 4049
rect 30288 4072 30340 4078
rect 29880 4040 29882 4049
rect 30288 4014 30340 4020
rect 29826 3975 29882 3984
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 28356 3664 28408 3670
rect 28356 3606 28408 3612
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27618 3224 27674 3233
rect 27252 3188 27304 3194
rect 28000 3194 28028 3470
rect 27618 3159 27674 3168
rect 27988 3188 28040 3194
rect 27252 3130 27304 3136
rect 27068 2984 27120 2990
rect 27264 2961 27292 3130
rect 27068 2926 27120 2932
rect 27250 2952 27306 2961
rect 26516 2916 26568 2922
rect 27632 2922 27660 3159
rect 27988 3130 28040 3136
rect 27250 2887 27306 2896
rect 27620 2916 27672 2922
rect 26516 2858 26568 2864
rect 27620 2858 27672 2864
rect 28368 2854 28396 3606
rect 28356 2848 28408 2854
rect 28356 2790 28408 2796
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 26330 2680 26386 2689
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 26240 2644 26292 2650
rect 27622 2672 27918 2692
rect 26330 2615 26386 2624
rect 26240 2586 26292 2592
rect 26344 2514 26372 2615
rect 27894 2544 27950 2553
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 27436 2508 27488 2514
rect 27894 2479 27896 2488
rect 27436 2450 27488 2456
rect 27948 2479 27950 2488
rect 27896 2450 27948 2456
rect 26238 2408 26294 2417
rect 26238 2343 26240 2352
rect 26292 2343 26294 2352
rect 26240 2314 26292 2320
rect 27448 2310 27476 2450
rect 26516 2304 26568 2310
rect 26514 2272 26516 2281
rect 27436 2304 27488 2310
rect 26568 2272 26570 2281
rect 26514 2207 26570 2216
rect 27434 2272 27436 2281
rect 27488 2272 27490 2281
rect 27434 2207 27490 2216
rect 28368 480 28396 2790
rect 29104 2650 29132 3674
rect 29552 3528 29604 3534
rect 29550 3496 29552 3505
rect 29604 3496 29606 3505
rect 29550 3431 29606 3440
rect 30104 3460 30156 3466
rect 29564 3194 29592 3431
rect 30104 3402 30156 3408
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 30116 3058 30144 3402
rect 30300 3097 30328 4014
rect 30472 3936 30524 3942
rect 30472 3878 30524 3884
rect 30484 3641 30512 3878
rect 30470 3632 30526 3641
rect 30470 3567 30526 3576
rect 30286 3088 30342 3097
rect 29460 3052 29512 3058
rect 29460 2994 29512 3000
rect 30104 3052 30156 3058
rect 30286 3023 30342 3032
rect 30104 2994 30156 3000
rect 29472 2650 29500 2994
rect 29552 2916 29604 2922
rect 29552 2858 29604 2864
rect 29092 2644 29144 2650
rect 29092 2586 29144 2592
rect 29460 2644 29512 2650
rect 29460 2586 29512 2592
rect 29564 2582 29592 2858
rect 29828 2848 29880 2854
rect 29828 2790 29880 2796
rect 29552 2576 29604 2582
rect 29552 2518 29604 2524
rect 29840 2514 29868 2790
rect 30116 2530 30144 2994
rect 30116 2514 30420 2530
rect 29828 2508 29880 2514
rect 30116 2508 30432 2514
rect 30116 2502 30380 2508
rect 29828 2450 29880 2456
rect 30380 2450 30432 2456
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 28920 1601 28948 2246
rect 28906 1592 28962 1601
rect 28906 1527 28962 1536
rect 31588 1306 31616 4655
rect 33980 2689 34008 8463
rect 34164 8362 34192 8570
rect 34716 8498 34744 8774
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34152 8356 34204 8362
rect 34152 8298 34204 8304
rect 34164 8022 34192 8298
rect 34152 8016 34204 8022
rect 34152 7958 34204 7964
rect 34164 7546 34192 7958
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 34152 7540 34204 7546
rect 34152 7482 34204 7488
rect 34428 7336 34480 7342
rect 34716 7290 34744 8434
rect 35268 8401 35296 8434
rect 35254 8392 35310 8401
rect 35254 8327 35310 8336
rect 35360 7970 35388 11630
rect 35452 11218 35480 11727
rect 35636 11354 35664 11999
rect 35728 11898 35756 12815
rect 35716 11892 35768 11898
rect 35716 11834 35768 11840
rect 35624 11348 35676 11354
rect 35624 11290 35676 11296
rect 35440 11212 35492 11218
rect 35440 11154 35492 11160
rect 35900 11212 35952 11218
rect 35900 11154 35952 11160
rect 35912 10810 35940 11154
rect 35900 10804 35952 10810
rect 35900 10746 35952 10752
rect 35808 10532 35860 10538
rect 35860 10492 35940 10520
rect 35808 10474 35860 10480
rect 35820 10266 35848 10474
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 35912 9586 35940 10492
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 36096 10130 36124 10406
rect 36372 10266 36400 14583
rect 36544 11688 36596 11694
rect 36544 11630 36596 11636
rect 36556 11393 36584 11630
rect 36542 11384 36598 11393
rect 36542 11319 36598 11328
rect 36450 11112 36506 11121
rect 36450 11047 36506 11056
rect 36464 10266 36492 11047
rect 36648 10810 36676 15535
rect 37462 15520 37518 16000
rect 37476 11914 37504 15520
rect 37200 11898 37504 11914
rect 37188 11892 37504 11898
rect 37240 11886 37504 11892
rect 37188 11834 37240 11840
rect 37004 11212 37056 11218
rect 37004 11154 37056 11160
rect 36726 11112 36782 11121
rect 36726 11047 36728 11056
rect 36780 11047 36782 11056
rect 36728 11018 36780 11024
rect 37016 10810 37044 11154
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 37004 10804 37056 10810
rect 37004 10746 37056 10752
rect 37280 10464 37332 10470
rect 37278 10432 37280 10441
rect 37332 10432 37334 10441
rect 37278 10367 37334 10376
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 36452 10260 36504 10266
rect 36452 10202 36504 10208
rect 36084 10124 36136 10130
rect 36084 10066 36136 10072
rect 35900 9580 35952 9586
rect 35900 9522 35952 9528
rect 36096 9518 36124 10066
rect 36084 9512 36136 9518
rect 36082 9480 36084 9489
rect 36136 9480 36138 9489
rect 36464 9466 36492 10202
rect 36464 9450 36584 9466
rect 36082 9415 36138 9424
rect 36360 9444 36412 9450
rect 36464 9444 36596 9450
rect 36464 9438 36544 9444
rect 36360 9386 36412 9392
rect 36544 9386 36596 9392
rect 36728 9444 36780 9450
rect 36728 9386 36780 9392
rect 36372 9178 36400 9386
rect 36634 9344 36690 9353
rect 36634 9279 36690 9288
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 35900 9104 35952 9110
rect 35900 9046 35952 9052
rect 35912 8634 35940 9046
rect 36268 8968 36320 8974
rect 36268 8910 36320 8916
rect 36280 8634 36308 8910
rect 36648 8634 36676 9279
rect 36740 9178 36768 9386
rect 36728 9172 36780 9178
rect 36728 9114 36780 9120
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 36268 8628 36320 8634
rect 36268 8570 36320 8576
rect 36636 8628 36688 8634
rect 36636 8570 36688 8576
rect 36634 8528 36690 8537
rect 36634 8463 36690 8472
rect 36084 8424 36136 8430
rect 35990 8392 36046 8401
rect 36084 8366 36136 8372
rect 35990 8327 36046 8336
rect 36004 8022 36032 8327
rect 35176 7954 35388 7970
rect 35440 8016 35492 8022
rect 35440 7958 35492 7964
rect 35992 8016 36044 8022
rect 35992 7958 36044 7964
rect 35164 7948 35388 7954
rect 35216 7942 35388 7948
rect 35164 7890 35216 7896
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 34900 7478 34928 7686
rect 34888 7472 34940 7478
rect 34888 7414 34940 7420
rect 35360 7410 35388 7822
rect 35452 7546 35480 7958
rect 36096 7834 36124 8366
rect 36004 7806 36124 7834
rect 35440 7540 35492 7546
rect 35440 7482 35492 7488
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 34480 7284 34744 7290
rect 34428 7278 34744 7284
rect 34440 7262 34744 7278
rect 34612 6928 34664 6934
rect 34612 6870 34664 6876
rect 34152 6792 34204 6798
rect 34152 6734 34204 6740
rect 34164 5914 34192 6734
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 34624 6390 34652 6870
rect 34612 6384 34664 6390
rect 34612 6326 34664 6332
rect 34612 6248 34664 6254
rect 34612 6190 34664 6196
rect 34624 6118 34652 6190
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 34152 5908 34204 5914
rect 34152 5850 34204 5856
rect 34624 5846 34652 6054
rect 34716 5846 34744 7262
rect 34794 7168 34850 7177
rect 34794 7103 34850 7112
rect 34612 5840 34664 5846
rect 34612 5782 34664 5788
rect 34704 5840 34756 5846
rect 34808 5817 34836 7103
rect 35360 7002 35388 7346
rect 35348 6996 35400 7002
rect 35348 6938 35400 6944
rect 35360 6322 35388 6938
rect 35348 6316 35400 6322
rect 35348 6258 35400 6264
rect 35900 6248 35952 6254
rect 35900 6190 35952 6196
rect 34980 6180 35032 6186
rect 34980 6122 35032 6128
rect 34992 5914 35020 6122
rect 34980 5908 35032 5914
rect 34980 5850 35032 5856
rect 34704 5782 34756 5788
rect 34794 5808 34850 5817
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 34164 5370 34192 5646
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 34624 5370 34652 5782
rect 34794 5743 34850 5752
rect 34992 5370 35020 5850
rect 34152 5364 34204 5370
rect 34152 5306 34204 5312
rect 34612 5364 34664 5370
rect 34612 5306 34664 5312
rect 34980 5364 35032 5370
rect 34980 5306 35032 5312
rect 35440 5024 35492 5030
rect 34702 4992 34758 5001
rect 35440 4966 35492 4972
rect 34702 4927 34758 4936
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 34289 3216 34585 3236
rect 33966 2680 34022 2689
rect 33966 2615 34022 2624
rect 31668 2304 31720 2310
rect 31668 2246 31720 2252
rect 31680 1465 31708 2246
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 31666 1456 31722 1465
rect 31666 1391 31722 1400
rect 31588 1278 31708 1306
rect 31680 480 31708 1278
rect 34716 513 34744 4927
rect 35452 4865 35480 4966
rect 35438 4856 35494 4865
rect 35438 4791 35494 4800
rect 35452 4282 35480 4791
rect 35440 4276 35492 4282
rect 35440 4218 35492 4224
rect 35806 2952 35862 2961
rect 35912 2938 35940 6190
rect 36004 5778 36032 7806
rect 36648 7546 36676 8463
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36452 7336 36504 7342
rect 36452 7278 36504 7284
rect 36176 6928 36228 6934
rect 36176 6870 36228 6876
rect 36084 6792 36136 6798
rect 36084 6734 36136 6740
rect 36096 6458 36124 6734
rect 36084 6452 36136 6458
rect 36084 6394 36136 6400
rect 36188 6390 36216 6870
rect 36360 6792 36412 6798
rect 36464 6769 36492 7278
rect 36360 6734 36412 6740
rect 36450 6760 36506 6769
rect 36176 6384 36228 6390
rect 36176 6326 36228 6332
rect 36372 5846 36400 6734
rect 36450 6695 36506 6704
rect 36452 6452 36504 6458
rect 36452 6394 36504 6400
rect 36464 5914 36492 6394
rect 36452 5908 36504 5914
rect 36452 5850 36504 5856
rect 36360 5840 36412 5846
rect 36360 5782 36412 5788
rect 35992 5772 36044 5778
rect 35992 5714 36044 5720
rect 36004 5030 36032 5714
rect 35992 5024 36044 5030
rect 35992 4966 36044 4972
rect 35862 2910 35940 2938
rect 35806 2887 35862 2896
rect 34978 1592 35034 1601
rect 34978 1527 35034 1536
rect 34702 504 34758 513
rect 4250 439 4306 448
rect 4986 0 5042 480
rect 8298 0 8354 480
rect 11610 0 11666 480
rect 15014 0 15070 480
rect 18326 0 18382 480
rect 21638 0 21694 480
rect 24950 0 25006 480
rect 28354 0 28410 480
rect 31666 0 31722 480
rect 34992 480 35020 1527
rect 35820 1329 35848 2887
rect 36004 2553 36032 4966
rect 35990 2544 36046 2553
rect 35990 2479 36046 2488
rect 38290 1456 38346 1465
rect 38290 1391 38346 1400
rect 35806 1320 35862 1329
rect 35806 1255 35862 1264
rect 38304 480 38332 1391
rect 34702 439 34758 448
rect 34978 0 35034 480
rect 38290 0 38346 480
<< via2 >>
rect 2686 15544 2742 15600
rect 1582 14592 1638 14648
rect 1490 13776 1546 13832
rect 1582 12008 1638 12064
rect 2042 11772 2044 11792
rect 2044 11772 2096 11792
rect 2096 11772 2098 11792
rect 2042 11736 2098 11772
rect 1582 11076 1638 11112
rect 1582 11056 1584 11076
rect 1584 11056 1636 11076
rect 1636 11056 1638 11076
rect 1582 10240 1638 10296
rect 2042 10412 2044 10432
rect 2044 10412 2096 10432
rect 2096 10412 2098 10432
rect 2042 10376 2098 10412
rect 1674 10004 1676 10024
rect 1676 10004 1728 10024
rect 1728 10004 1730 10024
rect 1674 9968 1730 10004
rect 1490 9036 1546 9072
rect 1490 9016 1492 9036
rect 1492 9016 1544 9036
rect 1544 9016 1546 9036
rect 1582 8472 1638 8528
rect 1950 3440 2006 3496
rect 2410 11192 2466 11248
rect 2502 10240 2558 10296
rect 36634 15544 36690 15600
rect 3790 12824 3846 12880
rect 2686 9424 2742 9480
rect 2226 7248 2282 7304
rect 2962 11736 3018 11792
rect 3054 10548 3056 10568
rect 3056 10548 3108 10568
rect 3108 10548 3110 10568
rect 3054 10512 3110 10548
rect 4802 11212 4858 11248
rect 4802 11192 4804 11212
rect 4804 11192 4856 11212
rect 4856 11192 4858 11212
rect 3146 10104 3202 10160
rect 3054 7520 3110 7576
rect 3882 10376 3938 10432
rect 3422 9016 3478 9072
rect 3974 9288 4030 9344
rect 3882 8880 3938 8936
rect 3790 7928 3846 7984
rect 2962 5480 3018 5536
rect 2870 3984 2926 4040
rect 2962 3848 3018 3904
rect 3330 4020 3332 4040
rect 3332 4020 3384 4040
rect 3384 4020 3386 4040
rect 3330 3984 3386 4020
rect 3698 3732 3754 3768
rect 3698 3712 3700 3732
rect 3700 3712 3752 3732
rect 3752 3712 3754 3732
rect 3790 3032 3846 3088
rect 4158 10260 4214 10296
rect 4158 10240 4160 10260
rect 4160 10240 4212 10260
rect 4212 10240 4214 10260
rect 4342 9424 4398 9480
rect 4526 9460 4528 9480
rect 4528 9460 4580 9480
rect 4580 9460 4582 9480
rect 4526 9424 4582 9460
rect 3974 4020 3976 4040
rect 3976 4020 4028 4040
rect 4028 4020 4030 4040
rect 3974 3984 4030 4020
rect 4618 9152 4674 9208
rect 4434 3440 4490 3496
rect 1674 2352 1730 2408
rect 2226 2216 2282 2272
rect 5170 8336 5226 8392
rect 4802 5752 4858 5808
rect 5354 8200 5410 8256
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 8942 11464 8998 11520
rect 5906 11056 5962 11112
rect 7470 11056 7526 11112
rect 8114 11056 8170 11112
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 5630 7792 5686 7848
rect 5722 6976 5778 7032
rect 5906 6296 5962 6352
rect 4894 5208 4950 5264
rect 5998 5480 6054 5536
rect 4250 3032 4306 3088
rect 4710 3032 4766 3088
rect 4158 1944 4214 2000
rect 4158 1264 4214 1320
rect 4894 2624 4950 2680
rect 4250 448 4306 504
rect 5722 4120 5778 4176
rect 5998 3984 6054 4040
rect 5906 3884 5908 3904
rect 5908 3884 5960 3904
rect 5960 3884 5962 3904
rect 5906 3848 5962 3884
rect 6734 8472 6790 8528
rect 6274 4528 6330 4584
rect 6182 3440 6238 3496
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 7838 9324 7840 9344
rect 7840 9324 7892 9344
rect 7892 9324 7894 9344
rect 7838 9288 7894 9324
rect 8206 9560 8262 9616
rect 8574 9424 8630 9480
rect 8298 9152 8354 9208
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 8206 8744 8262 8800
rect 7838 8372 7840 8392
rect 7840 8372 7892 8392
rect 7892 8372 7894 8392
rect 7838 8336 7894 8372
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 7286 7384 7342 7440
rect 8850 8880 8906 8936
rect 8390 8744 8446 8800
rect 8206 6840 8262 6896
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 8758 8200 8814 8256
rect 10046 10920 10102 10976
rect 9954 10784 10010 10840
rect 8758 7112 8814 7168
rect 8666 6296 8722 6352
rect 9126 5752 9182 5808
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 6642 3984 6698 4040
rect 6550 3732 6606 3768
rect 6550 3712 6552 3732
rect 6552 3712 6604 3732
rect 6604 3712 6606 3732
rect 6366 3596 6422 3632
rect 6366 3576 6368 3596
rect 6368 3576 6420 3596
rect 6420 3576 6422 3596
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7378 4004 7434 4040
rect 7378 3984 7380 4004
rect 7380 3984 7432 4004
rect 7432 3984 7434 4004
rect 9126 5364 9182 5400
rect 9126 5344 9128 5364
rect 9128 5344 9180 5364
rect 9180 5344 9182 5364
rect 8758 3848 8814 3904
rect 9678 10138 9734 10194
rect 9310 9968 9366 10024
rect 9678 9832 9734 9888
rect 9678 8472 9734 8528
rect 9494 8372 9496 8392
rect 9496 8372 9548 8392
rect 9548 8372 9550 8392
rect 9494 8336 9550 8372
rect 11150 9832 11206 9888
rect 10782 8336 10838 8392
rect 10966 8200 11022 8256
rect 11058 7928 11114 7984
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 15474 11600 15530 11656
rect 12438 11464 12494 11520
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 13174 11076 13230 11112
rect 13174 11056 13176 11076
rect 13176 11056 13228 11076
rect 13228 11056 13230 11076
rect 12530 9580 12586 9616
rect 12530 9560 12532 9580
rect 12532 9560 12584 9580
rect 12584 9560 12586 9580
rect 11794 8200 11850 8256
rect 9954 7420 9956 7440
rect 9956 7420 10008 7440
rect 10008 7420 10010 7440
rect 9954 7384 10010 7420
rect 11334 7928 11390 7984
rect 11058 7384 11114 7440
rect 10506 6976 10562 7032
rect 9586 5908 9642 5944
rect 9586 5888 9588 5908
rect 9588 5888 9640 5908
rect 9640 5888 9642 5908
rect 9586 5752 9642 5808
rect 9586 3848 9642 3904
rect 9218 3732 9274 3768
rect 9218 3712 9220 3732
rect 9220 3712 9272 3732
rect 9272 3712 9274 3732
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 8850 3576 8906 3632
rect 9034 3576 9090 3632
rect 9954 4020 9956 4040
rect 9956 4020 10008 4040
rect 10008 4020 10010 4040
rect 9954 3984 10010 4020
rect 8850 2644 8906 2680
rect 10138 4120 10194 4176
rect 10690 6432 10746 6488
rect 10874 6180 10930 6216
rect 10874 6160 10876 6180
rect 10876 6160 10928 6180
rect 10928 6160 10930 6180
rect 10690 5752 10746 5808
rect 10506 5480 10562 5536
rect 10874 5636 10930 5672
rect 10874 5616 10876 5636
rect 10876 5616 10928 5636
rect 10928 5616 10930 5636
rect 11518 5480 11574 5536
rect 11518 4120 11574 4176
rect 13082 9968 13138 10024
rect 12806 8336 12862 8392
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 13726 9832 13782 9888
rect 13450 8200 13506 8256
rect 12622 7284 12624 7304
rect 12624 7284 12676 7304
rect 12676 7284 12678 7304
rect 12622 7248 12678 7284
rect 13818 7948 13874 7984
rect 13818 7928 13820 7948
rect 13820 7928 13872 7948
rect 13872 7928 13874 7948
rect 12714 7112 12770 7168
rect 12162 5616 12218 5672
rect 12254 5480 12310 5536
rect 12898 6160 12954 6216
rect 12162 5208 12218 5264
rect 10138 3440 10194 3496
rect 8850 2624 8852 2644
rect 8852 2624 8904 2644
rect 8904 2624 8906 2644
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 12622 4684 12678 4720
rect 12622 4664 12624 4684
rect 12624 4664 12676 4684
rect 12676 4664 12678 4684
rect 12162 3712 12218 3768
rect 12254 3612 12256 3632
rect 12256 3612 12308 3632
rect 12308 3612 12310 3632
rect 12254 3576 12310 3612
rect 13082 5208 13138 5264
rect 13818 7792 13874 7848
rect 14094 8880 14150 8936
rect 13910 6160 13966 6216
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 14738 8200 14794 8256
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 15290 7540 15346 7576
rect 15290 7520 15292 7540
rect 15292 7520 15344 7540
rect 15344 7520 15346 7540
rect 14922 6432 14978 6488
rect 14186 6296 14242 6352
rect 15198 6160 15254 6216
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 14830 5616 14886 5672
rect 14186 5480 14242 5536
rect 14094 5364 14150 5400
rect 14094 5344 14096 5364
rect 14096 5344 14148 5364
rect 14148 5344 14150 5364
rect 13542 4800 13598 4856
rect 14738 4936 14794 4992
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14370 3440 14426 3496
rect 14186 3052 14242 3088
rect 14186 3032 14188 3052
rect 14188 3032 14240 3052
rect 14240 3032 14242 3052
rect 14646 2896 14702 2952
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 13358 2508 13414 2544
rect 15014 4392 15070 4448
rect 15842 11464 15898 11520
rect 16026 10920 16082 10976
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 18602 11636 18604 11656
rect 18604 11636 18656 11656
rect 18656 11636 18658 11656
rect 18602 11600 18658 11636
rect 18234 11328 18290 11384
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 19430 11500 19432 11520
rect 19432 11500 19484 11520
rect 19484 11500 19486 11520
rect 19430 11464 19486 11500
rect 16946 8744 17002 8800
rect 16026 8372 16028 8392
rect 16028 8372 16080 8392
rect 16080 8372 16082 8392
rect 16026 8336 16082 8372
rect 16670 7792 16726 7848
rect 16578 6976 16634 7032
rect 16210 6432 16266 6488
rect 16578 6452 16634 6488
rect 16578 6432 16580 6452
rect 16580 6432 16632 6452
rect 16632 6432 16634 6452
rect 17406 9460 17408 9480
rect 17408 9460 17460 9480
rect 17460 9460 17462 9480
rect 17406 9424 17462 9460
rect 17866 9036 17922 9072
rect 17866 9016 17868 9036
rect 17868 9016 17920 9036
rect 17920 9016 17922 9036
rect 18786 10648 18842 10704
rect 18234 9696 18290 9752
rect 18050 8030 18106 8086
rect 17682 7520 17738 7576
rect 17498 6296 17554 6352
rect 17682 5888 17738 5944
rect 17866 6160 17922 6216
rect 17774 4972 17776 4992
rect 17776 4972 17828 4992
rect 17828 4972 17830 4992
rect 17774 4936 17830 4972
rect 17130 4564 17132 4584
rect 17132 4564 17184 4584
rect 17184 4564 17186 4584
rect 17130 4528 17186 4564
rect 15842 3732 15898 3768
rect 15842 3712 15844 3732
rect 15844 3712 15896 3732
rect 15896 3712 15898 3732
rect 17038 4392 17094 4448
rect 18878 10376 18934 10432
rect 18786 7520 18842 7576
rect 18694 6704 18750 6760
rect 18418 4800 18474 4856
rect 13358 2488 13360 2508
rect 13360 2488 13412 2508
rect 13412 2488 13414 2508
rect 12898 1944 12954 2000
rect 11978 1808 12034 1864
rect 15198 2388 15200 2408
rect 15200 2388 15252 2408
rect 15252 2388 15254 2408
rect 15198 2352 15254 2388
rect 20718 11600 20774 11656
rect 19338 11056 19394 11112
rect 24306 11736 24362 11792
rect 20718 10784 20774 10840
rect 23386 11328 23442 11384
rect 24122 11192 24178 11248
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 19798 8880 19854 8936
rect 19982 8916 19984 8936
rect 19984 8916 20036 8936
rect 20036 8916 20038 8936
rect 19982 8880 20038 8916
rect 19430 8236 19432 8256
rect 19432 8236 19484 8256
rect 19484 8236 19486 8256
rect 19430 8200 19486 8236
rect 19430 7792 19486 7848
rect 19430 7520 19486 7576
rect 19246 6976 19302 7032
rect 20166 7384 20222 7440
rect 19890 5908 19946 5944
rect 19890 5888 19892 5908
rect 19892 5888 19944 5908
rect 19944 5888 19946 5908
rect 20994 10004 20996 10024
rect 20996 10004 21048 10024
rect 21048 10004 21050 10024
rect 20994 9968 21050 10004
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 21730 10920 21786 10976
rect 23110 10804 23166 10840
rect 23110 10784 23112 10804
rect 23112 10784 23164 10804
rect 23164 10784 23166 10804
rect 21546 10376 21602 10432
rect 21454 10240 21510 10296
rect 21362 9832 21418 9888
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 21270 8336 21326 8392
rect 21454 8336 21510 8392
rect 20810 7692 20812 7712
rect 20812 7692 20864 7712
rect 20864 7692 20866 7712
rect 20810 7656 20866 7692
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20718 6740 20720 6760
rect 20720 6740 20772 6760
rect 20772 6740 20774 6760
rect 20718 6704 20774 6740
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 22926 10412 22928 10432
rect 22928 10412 22980 10432
rect 22980 10412 22982 10432
rect 22926 10376 22982 10412
rect 23478 10240 23534 10296
rect 22742 8880 22798 8936
rect 23294 7248 23350 7304
rect 19982 4664 20038 4720
rect 19154 3440 19210 3496
rect 18786 3032 18842 3088
rect 19154 2796 19156 2816
rect 19156 2796 19208 2816
rect 19208 2796 19210 2816
rect 19154 2760 19210 2796
rect 19890 3848 19946 3904
rect 19338 2896 19394 2952
rect 19522 2760 19578 2816
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21270 5208 21326 5264
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20902 3712 20958 3768
rect 21086 3576 21142 3632
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20258 2488 20314 2544
rect 23110 5888 23166 5944
rect 23386 6432 23442 6488
rect 23478 6160 23534 6216
rect 22742 4800 22798 4856
rect 23478 5072 23534 5128
rect 22650 3576 22706 3632
rect 23202 4120 23258 4176
rect 21638 2760 21694 2816
rect 21362 2372 21418 2408
rect 21362 2352 21364 2372
rect 21364 2352 21416 2372
rect 21416 2352 21418 2372
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 20810 1808 20866 1864
rect 22558 2932 22560 2952
rect 22560 2932 22612 2952
rect 22612 2932 22614 2952
rect 22558 2896 22614 2932
rect 24950 10648 25006 10704
rect 24398 9288 24454 9344
rect 25042 10004 25044 10024
rect 25044 10004 25096 10024
rect 25096 10004 25098 10024
rect 25042 9968 25098 10004
rect 25226 9016 25282 9072
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 29734 11736 29790 11792
rect 27618 10956 27620 10976
rect 27620 10956 27672 10976
rect 27672 10956 27674 10976
rect 27618 10920 27674 10956
rect 25962 9832 26018 9888
rect 23938 7384 23994 7440
rect 25778 8336 25834 8392
rect 25226 8200 25282 8256
rect 24030 6860 24086 6896
rect 24030 6840 24032 6860
rect 24032 6840 24084 6860
rect 24084 6840 24086 6860
rect 24582 6332 24584 6352
rect 24584 6332 24636 6352
rect 24636 6332 24638 6352
rect 24582 6296 24638 6332
rect 24122 5636 24178 5672
rect 24122 5616 24124 5636
rect 24124 5616 24176 5636
rect 24176 5616 24178 5636
rect 23570 4392 23626 4448
rect 24950 4936 25006 4992
rect 23846 3168 23902 3224
rect 22466 2488 22522 2544
rect 24766 2488 24822 2544
rect 22466 2216 22522 2272
rect 26054 8200 26110 8256
rect 26606 10376 26662 10432
rect 26514 9324 26516 9344
rect 26516 9324 26568 9344
rect 26568 9324 26570 9344
rect 26514 9288 26570 9324
rect 26330 9016 26386 9072
rect 26974 8880 27030 8936
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 27986 9832 28042 9888
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 26330 7520 26386 7576
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 27342 6432 27398 6488
rect 27158 6296 27214 6352
rect 26330 5752 26386 5808
rect 26882 5616 26938 5672
rect 27066 5480 27122 5536
rect 28170 6976 28226 7032
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 27342 4664 27398 4720
rect 25502 3984 25558 4040
rect 26422 3712 26478 3768
rect 27986 4120 28042 4176
rect 29090 5752 29146 5808
rect 29182 5616 29238 5672
rect 30010 11600 30066 11656
rect 29826 11192 29882 11248
rect 27802 4020 27804 4040
rect 27804 4020 27856 4040
rect 27856 4020 27858 4040
rect 27802 3984 27858 4020
rect 27066 3848 27122 3904
rect 26974 3440 27030 3496
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 30470 11328 30526 11384
rect 31666 11056 31722 11112
rect 31482 10104 31538 10160
rect 31114 10004 31116 10024
rect 31116 10004 31168 10024
rect 31168 10004 31170 10024
rect 31114 9968 31170 10004
rect 30746 9560 30802 9616
rect 36358 14592 36414 14648
rect 35622 13776 35678 13832
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 35714 12824 35770 12880
rect 32494 11056 32550 11112
rect 32402 9868 32404 9888
rect 32404 9868 32456 9888
rect 32456 9868 32458 9888
rect 32402 9832 32458 9868
rect 32034 9696 32090 9752
rect 30470 8336 30526 8392
rect 31574 8372 31576 8392
rect 31576 8372 31628 8392
rect 31628 8372 31630 8392
rect 31574 8336 31630 8372
rect 30562 7792 30618 7848
rect 31390 7384 31446 7440
rect 30562 7248 30618 7304
rect 30838 6432 30894 6488
rect 32218 6704 32274 6760
rect 30378 5480 30434 5536
rect 31298 5208 31354 5264
rect 32862 7384 32918 7440
rect 33230 7148 33232 7168
rect 33232 7148 33284 7168
rect 33284 7148 33286 7168
rect 33230 7112 33286 7148
rect 33690 11328 33746 11384
rect 33506 10784 33562 10840
rect 34058 11056 34114 11112
rect 34058 10920 34114 10976
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 35622 12008 35678 12064
rect 35438 11736 35494 11792
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 34610 10376 34666 10432
rect 34794 10240 34850 10296
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 34978 10104 35034 10160
rect 34886 10004 34888 10024
rect 34888 10004 34940 10024
rect 34940 10004 34942 10024
rect 34886 9968 34942 10004
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 33966 8472 34022 8528
rect 33782 6840 33838 6896
rect 33506 6432 33562 6488
rect 33414 6160 33470 6216
rect 32218 5072 32274 5128
rect 31758 4972 31760 4992
rect 31760 4972 31812 4992
rect 31812 4972 31814 4992
rect 31758 4936 31814 4972
rect 31574 4664 31630 4720
rect 30194 4276 30250 4312
rect 30194 4256 30196 4276
rect 30196 4256 30248 4276
rect 30248 4256 30250 4276
rect 29826 4020 29828 4040
rect 29828 4020 29880 4040
rect 29880 4020 29882 4040
rect 29826 3984 29882 4020
rect 27618 3168 27674 3224
rect 27250 2896 27306 2952
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 26330 2624 26386 2680
rect 27894 2508 27950 2544
rect 27894 2488 27896 2508
rect 27896 2488 27948 2508
rect 27948 2488 27950 2508
rect 26238 2372 26294 2408
rect 26238 2352 26240 2372
rect 26240 2352 26292 2372
rect 26292 2352 26294 2372
rect 26514 2252 26516 2272
rect 26516 2252 26568 2272
rect 26568 2252 26570 2272
rect 26514 2216 26570 2252
rect 27434 2252 27436 2272
rect 27436 2252 27488 2272
rect 27488 2252 27490 2272
rect 27434 2216 27490 2252
rect 29550 3476 29552 3496
rect 29552 3476 29604 3496
rect 29604 3476 29606 3496
rect 29550 3440 29606 3476
rect 30470 3576 30526 3632
rect 30286 3032 30342 3088
rect 28906 1536 28962 1592
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 35254 8336 35310 8392
rect 36542 11328 36598 11384
rect 36450 11056 36506 11112
rect 36726 11076 36782 11112
rect 36726 11056 36728 11076
rect 36728 11056 36780 11076
rect 36780 11056 36782 11076
rect 37278 10412 37280 10432
rect 37280 10412 37332 10432
rect 37332 10412 37334 10432
rect 37278 10376 37334 10412
rect 36082 9460 36084 9480
rect 36084 9460 36136 9480
rect 36136 9460 36138 9480
rect 36082 9424 36138 9460
rect 36634 9288 36690 9344
rect 36634 8472 36690 8528
rect 35990 8336 36046 8392
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 34794 7112 34850 7168
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 34794 5752 34850 5808
rect 34702 4936 34758 4992
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 33966 2624 34022 2680
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 31666 1400 31722 1456
rect 35438 4800 35494 4856
rect 35806 2896 35862 2952
rect 36450 6704 36506 6760
rect 34978 1536 35034 1592
rect 34702 448 34758 504
rect 35990 2488 36046 2544
rect 38290 1400 38346 1456
rect 35806 1264 35862 1320
<< metal3 >>
rect 0 15602 480 15632
rect 2681 15602 2747 15605
rect 0 15600 2747 15602
rect 0 15544 2686 15600
rect 2742 15544 2747 15600
rect 0 15542 2747 15544
rect 0 15512 480 15542
rect 2681 15539 2747 15542
rect 36629 15602 36695 15605
rect 39520 15602 40000 15632
rect 36629 15600 40000 15602
rect 36629 15544 36634 15600
rect 36690 15544 40000 15600
rect 36629 15542 40000 15544
rect 36629 15539 36695 15542
rect 39520 15512 40000 15542
rect 0 14650 480 14680
rect 1577 14650 1643 14653
rect 0 14648 1643 14650
rect 0 14592 1582 14648
rect 1638 14592 1643 14648
rect 0 14590 1643 14592
rect 0 14560 480 14590
rect 1577 14587 1643 14590
rect 36353 14650 36419 14653
rect 39520 14650 40000 14680
rect 36353 14648 40000 14650
rect 36353 14592 36358 14648
rect 36414 14592 40000 14648
rect 36353 14590 40000 14592
rect 36353 14587 36419 14590
rect 39520 14560 40000 14590
rect 0 13834 480 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 480 13774
rect 1485 13771 1551 13774
rect 35617 13834 35683 13837
rect 39520 13834 40000 13864
rect 35617 13832 40000 13834
rect 35617 13776 35622 13832
rect 35678 13776 40000 13832
rect 35617 13774 40000 13776
rect 35617 13771 35683 13774
rect 39520 13744 40000 13774
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 0 12882 480 12912
rect 3785 12882 3851 12885
rect 0 12880 3851 12882
rect 0 12824 3790 12880
rect 3846 12824 3851 12880
rect 0 12822 3851 12824
rect 0 12792 480 12822
rect 3785 12819 3851 12822
rect 35709 12882 35775 12885
rect 39520 12882 40000 12912
rect 35709 12880 40000 12882
rect 35709 12824 35714 12880
rect 35770 12824 40000 12880
rect 35709 12822 40000 12824
rect 35709 12819 35775 12822
rect 39520 12792 40000 12822
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 0 12066 480 12096
rect 1577 12066 1643 12069
rect 0 12064 1643 12066
rect 0 12008 1582 12064
rect 1638 12008 1643 12064
rect 0 12006 1643 12008
rect 0 11976 480 12006
rect 1577 12003 1643 12006
rect 35617 12066 35683 12069
rect 39520 12066 40000 12096
rect 35617 12064 40000 12066
rect 35617 12008 35622 12064
rect 35678 12008 40000 12064
rect 35617 12006 40000 12008
rect 35617 12003 35683 12006
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 39520 11976 40000 12006
rect 34277 11935 34597 11936
rect 2037 11794 2103 11797
rect 2957 11794 3023 11797
rect 24301 11794 24367 11797
rect 29729 11794 29795 11797
rect 35433 11794 35499 11797
rect 2037 11792 35499 11794
rect 2037 11736 2042 11792
rect 2098 11736 2962 11792
rect 3018 11736 24306 11792
rect 24362 11736 29734 11792
rect 29790 11736 35438 11792
rect 35494 11736 35499 11792
rect 2037 11734 35499 11736
rect 2037 11731 2103 11734
rect 2957 11731 3023 11734
rect 24301 11731 24367 11734
rect 29729 11731 29795 11734
rect 35433 11731 35499 11734
rect 15469 11658 15535 11661
rect 18597 11658 18663 11661
rect 15469 11656 18663 11658
rect 15469 11600 15474 11656
rect 15530 11600 18602 11656
rect 18658 11600 18663 11656
rect 15469 11598 18663 11600
rect 15469 11595 15535 11598
rect 18597 11595 18663 11598
rect 20713 11658 20779 11661
rect 30005 11658 30071 11661
rect 20713 11656 30071 11658
rect 20713 11600 20718 11656
rect 20774 11600 30010 11656
rect 30066 11600 30071 11656
rect 20713 11598 30071 11600
rect 20713 11595 20779 11598
rect 30005 11595 30071 11598
rect 8937 11522 9003 11525
rect 12433 11522 12499 11525
rect 8937 11520 12499 11522
rect 8937 11464 8942 11520
rect 8998 11464 12438 11520
rect 12494 11464 12499 11520
rect 8937 11462 12499 11464
rect 8937 11459 9003 11462
rect 12433 11459 12499 11462
rect 15837 11522 15903 11525
rect 19425 11522 19491 11525
rect 15837 11520 19491 11522
rect 15837 11464 15842 11520
rect 15898 11464 19430 11520
rect 19486 11464 19491 11520
rect 15837 11462 19491 11464
rect 15837 11459 15903 11462
rect 19425 11459 19491 11462
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 18229 11386 18295 11389
rect 23381 11386 23447 11389
rect 18229 11384 23447 11386
rect 18229 11328 18234 11384
rect 18290 11328 23386 11384
rect 23442 11328 23447 11384
rect 18229 11326 23447 11328
rect 18229 11323 18295 11326
rect 23381 11323 23447 11326
rect 30465 11386 30531 11389
rect 33685 11386 33751 11389
rect 36537 11386 36603 11389
rect 30465 11384 36603 11386
rect 30465 11328 30470 11384
rect 30526 11328 33690 11384
rect 33746 11328 36542 11384
rect 36598 11328 36603 11384
rect 30465 11326 36603 11328
rect 30465 11323 30531 11326
rect 33685 11323 33751 11326
rect 36537 11323 36603 11326
rect 2405 11250 2471 11253
rect 4797 11250 4863 11253
rect 24117 11250 24183 11253
rect 29821 11250 29887 11253
rect 2405 11248 29887 11250
rect 2405 11192 2410 11248
rect 2466 11192 4802 11248
rect 4858 11192 24122 11248
rect 24178 11192 29826 11248
rect 29882 11192 29887 11248
rect 2405 11190 29887 11192
rect 2405 11187 2471 11190
rect 4797 11187 4863 11190
rect 24117 11187 24183 11190
rect 29821 11187 29887 11190
rect 0 11114 480 11144
rect 1577 11114 1643 11117
rect 0 11112 1643 11114
rect 0 11056 1582 11112
rect 1638 11056 1643 11112
rect 0 11054 1643 11056
rect 0 11024 480 11054
rect 1577 11051 1643 11054
rect 5901 11114 5967 11117
rect 7465 11114 7531 11117
rect 5901 11112 7531 11114
rect 5901 11056 5906 11112
rect 5962 11056 7470 11112
rect 7526 11056 7531 11112
rect 5901 11054 7531 11056
rect 5901 11051 5967 11054
rect 7465 11051 7531 11054
rect 8109 11114 8175 11117
rect 13169 11114 13235 11117
rect 19333 11114 19399 11117
rect 8109 11112 19399 11114
rect 8109 11056 8114 11112
rect 8170 11056 13174 11112
rect 13230 11056 19338 11112
rect 19394 11056 19399 11112
rect 8109 11054 19399 11056
rect 8109 11051 8175 11054
rect 13169 11051 13235 11054
rect 19333 11051 19399 11054
rect 31661 11114 31727 11117
rect 32489 11114 32555 11117
rect 31661 11112 32555 11114
rect 31661 11056 31666 11112
rect 31722 11056 32494 11112
rect 32550 11056 32555 11112
rect 31661 11054 32555 11056
rect 31661 11051 31727 11054
rect 32489 11051 32555 11054
rect 34053 11114 34119 11117
rect 36445 11114 36511 11117
rect 34053 11112 36511 11114
rect 34053 11056 34058 11112
rect 34114 11056 36450 11112
rect 36506 11056 36511 11112
rect 34053 11054 36511 11056
rect 34053 11051 34119 11054
rect 36445 11051 36511 11054
rect 36721 11114 36787 11117
rect 39520 11114 40000 11144
rect 36721 11112 40000 11114
rect 36721 11056 36726 11112
rect 36782 11056 40000 11112
rect 36721 11054 40000 11056
rect 36721 11051 36787 11054
rect 39520 11024 40000 11054
rect 10041 10978 10107 10981
rect 16021 10978 16087 10981
rect 10041 10976 16087 10978
rect 10041 10920 10046 10976
rect 10102 10920 16026 10976
rect 16082 10920 16087 10976
rect 10041 10918 16087 10920
rect 10041 10915 10107 10918
rect 16021 10915 16087 10918
rect 21725 10978 21791 10981
rect 27613 10978 27679 10981
rect 21725 10976 27679 10978
rect 21725 10920 21730 10976
rect 21786 10920 27618 10976
rect 27674 10920 27679 10976
rect 21725 10918 27679 10920
rect 21725 10915 21791 10918
rect 27613 10915 27679 10918
rect 28942 10916 28948 10980
rect 29012 10978 29018 10980
rect 34053 10978 34119 10981
rect 29012 10976 34119 10978
rect 29012 10920 34058 10976
rect 34114 10920 34119 10976
rect 29012 10918 34119 10920
rect 29012 10916 29018 10918
rect 34053 10915 34119 10918
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 9949 10842 10015 10845
rect 20713 10842 20779 10845
rect 9949 10840 20779 10842
rect 9949 10784 9954 10840
rect 10010 10784 20718 10840
rect 20774 10784 20779 10840
rect 9949 10782 20779 10784
rect 9949 10779 10015 10782
rect 20713 10779 20779 10782
rect 23105 10842 23171 10845
rect 33501 10842 33567 10845
rect 23105 10840 33567 10842
rect 23105 10784 23110 10840
rect 23166 10784 33506 10840
rect 33562 10784 33567 10840
rect 23105 10782 33567 10784
rect 23105 10779 23171 10782
rect 33501 10779 33567 10782
rect 18781 10706 18847 10709
rect 24945 10706 25011 10709
rect 28942 10706 28948 10708
rect 18781 10704 28948 10706
rect 18781 10648 18786 10704
rect 18842 10648 24950 10704
rect 25006 10648 28948 10704
rect 18781 10646 28948 10648
rect 18781 10643 18847 10646
rect 24945 10643 25011 10646
rect 28942 10644 28948 10646
rect 29012 10644 29018 10708
rect 3049 10570 3115 10573
rect 3049 10568 28090 10570
rect 3049 10512 3054 10568
rect 3110 10512 28090 10568
rect 3049 10510 28090 10512
rect 3049 10507 3115 10510
rect 2037 10434 2103 10437
rect 3877 10434 3943 10437
rect 2037 10432 3943 10434
rect 2037 10376 2042 10432
rect 2098 10376 3882 10432
rect 3938 10376 3943 10432
rect 2037 10374 3943 10376
rect 2037 10371 2103 10374
rect 3877 10371 3943 10374
rect 18873 10434 18939 10437
rect 21541 10434 21607 10437
rect 18873 10432 21607 10434
rect 18873 10376 18878 10432
rect 18934 10376 21546 10432
rect 21602 10376 21607 10432
rect 18873 10374 21607 10376
rect 18873 10371 18939 10374
rect 21541 10371 21607 10374
rect 22921 10434 22987 10437
rect 26601 10434 26667 10437
rect 22921 10432 26667 10434
rect 22921 10376 22926 10432
rect 22982 10376 26606 10432
rect 26662 10376 26667 10432
rect 22921 10374 26667 10376
rect 28030 10434 28090 10510
rect 28942 10434 28948 10436
rect 28030 10374 28948 10434
rect 22921 10371 22987 10374
rect 26601 10371 26667 10374
rect 28942 10372 28948 10374
rect 29012 10372 29018 10436
rect 34605 10434 34671 10437
rect 37273 10434 37339 10437
rect 34605 10432 37339 10434
rect 34605 10376 34610 10432
rect 34666 10376 37278 10432
rect 37334 10376 37339 10432
rect 34605 10374 37339 10376
rect 34605 10371 34671 10374
rect 37273 10371 37339 10374
rect 14277 10368 14597 10369
rect 0 10298 480 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 480 10238
rect 1577 10235 1643 10238
rect 2497 10298 2563 10301
rect 4153 10298 4219 10301
rect 2497 10296 4219 10298
rect 2497 10240 2502 10296
rect 2558 10240 4158 10296
rect 4214 10240 4219 10296
rect 2497 10238 4219 10240
rect 2497 10235 2563 10238
rect 4153 10235 4219 10238
rect 21449 10298 21515 10301
rect 23473 10298 23539 10301
rect 21449 10296 23539 10298
rect 21449 10240 21454 10296
rect 21510 10240 23478 10296
rect 23534 10240 23539 10296
rect 21449 10238 23539 10240
rect 21449 10235 21515 10238
rect 23473 10235 23539 10238
rect 34789 10298 34855 10301
rect 39520 10298 40000 10328
rect 34789 10296 40000 10298
rect 34789 10240 34794 10296
rect 34850 10240 40000 10296
rect 34789 10238 40000 10240
rect 34789 10235 34855 10238
rect 39520 10208 40000 10238
rect 9673 10196 9739 10199
rect 9630 10194 9739 10196
rect 3141 10162 3207 10165
rect 9630 10162 9678 10194
rect 3141 10160 9678 10162
rect 3141 10104 3146 10160
rect 3202 10138 9678 10160
rect 9734 10138 9739 10194
rect 3202 10133 9739 10138
rect 31477 10162 31543 10165
rect 34973 10162 35039 10165
rect 31477 10160 35039 10162
rect 3202 10104 9690 10133
rect 3141 10102 9690 10104
rect 31477 10104 31482 10160
rect 31538 10104 34978 10160
rect 35034 10104 35039 10160
rect 31477 10102 35039 10104
rect 3141 10099 3207 10102
rect 31477 10099 31543 10102
rect 34973 10099 35039 10102
rect 1669 10026 1735 10029
rect 9305 10026 9371 10029
rect 13077 10026 13143 10029
rect 1669 10024 9138 10026
rect 1669 9968 1674 10024
rect 1730 9968 9138 10024
rect 1669 9966 9138 9968
rect 1669 9963 1735 9966
rect 9078 9890 9138 9966
rect 9305 10024 13143 10026
rect 9305 9968 9310 10024
rect 9366 9968 13082 10024
rect 13138 9968 13143 10024
rect 9305 9966 13143 9968
rect 9305 9963 9371 9966
rect 13077 9963 13143 9966
rect 20989 10026 21055 10029
rect 25037 10026 25103 10029
rect 20989 10024 25103 10026
rect 20989 9968 20994 10024
rect 21050 9968 25042 10024
rect 25098 9968 25103 10024
rect 20989 9966 25103 9968
rect 20989 9963 21055 9966
rect 25037 9963 25103 9966
rect 31109 10026 31175 10029
rect 34881 10026 34947 10029
rect 31109 10024 34947 10026
rect 31109 9968 31114 10024
rect 31170 9968 34886 10024
rect 34942 9968 34947 10024
rect 31109 9966 34947 9968
rect 31109 9963 31175 9966
rect 34881 9963 34947 9966
rect 9673 9890 9739 9893
rect 11145 9890 11211 9893
rect 13721 9890 13787 9893
rect 9078 9888 9874 9890
rect 9078 9832 9678 9888
rect 9734 9832 9874 9888
rect 9078 9830 9874 9832
rect 9673 9827 9739 9830
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 9814 9754 9874 9830
rect 11145 9888 13787 9890
rect 11145 9832 11150 9888
rect 11206 9832 13726 9888
rect 13782 9832 13787 9888
rect 11145 9830 13787 9832
rect 11145 9827 11211 9830
rect 13721 9827 13787 9830
rect 21357 9890 21423 9893
rect 25957 9890 26023 9893
rect 21357 9888 26023 9890
rect 21357 9832 21362 9888
rect 21418 9832 25962 9888
rect 26018 9832 26023 9888
rect 21357 9830 26023 9832
rect 21357 9827 21423 9830
rect 25957 9827 26023 9830
rect 27981 9890 28047 9893
rect 32397 9890 32463 9893
rect 27981 9888 32463 9890
rect 27981 9832 27986 9888
rect 28042 9832 32402 9888
rect 32458 9832 32463 9888
rect 27981 9830 32463 9832
rect 27981 9827 28047 9830
rect 32397 9827 32463 9830
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 18229 9754 18295 9757
rect 9814 9752 18295 9754
rect 9814 9696 18234 9752
rect 18290 9696 18295 9752
rect 9814 9694 18295 9696
rect 18229 9691 18295 9694
rect 28942 9692 28948 9756
rect 29012 9754 29018 9756
rect 32029 9754 32095 9757
rect 29012 9752 32095 9754
rect 29012 9696 32034 9752
rect 32090 9696 32095 9752
rect 29012 9694 32095 9696
rect 29012 9692 29018 9694
rect 32029 9691 32095 9694
rect 8201 9618 8267 9621
rect 12525 9618 12591 9621
rect 30741 9618 30807 9621
rect 8201 9616 12591 9618
rect 8201 9560 8206 9616
rect 8262 9560 12530 9616
rect 12586 9560 12591 9616
rect 8201 9558 12591 9560
rect 8201 9555 8267 9558
rect 12525 9555 12591 9558
rect 14046 9616 30807 9618
rect 14046 9560 30746 9616
rect 30802 9560 30807 9616
rect 14046 9558 30807 9560
rect 2681 9482 2747 9485
rect 4337 9482 4403 9485
rect 2681 9480 4403 9482
rect 2681 9424 2686 9480
rect 2742 9424 4342 9480
rect 4398 9424 4403 9480
rect 2681 9422 4403 9424
rect 2681 9419 2747 9422
rect 4337 9419 4403 9422
rect 4521 9482 4587 9485
rect 8569 9482 8635 9485
rect 4521 9480 8635 9482
rect 4521 9424 4526 9480
rect 4582 9424 8574 9480
rect 8630 9424 8635 9480
rect 4521 9422 8635 9424
rect 4521 9419 4587 9422
rect 8569 9419 8635 9422
rect 0 9346 480 9376
rect 3969 9346 4035 9349
rect 0 9344 4035 9346
rect 0 9288 3974 9344
rect 4030 9288 4035 9344
rect 0 9286 4035 9288
rect 0 9256 480 9286
rect 3969 9283 4035 9286
rect 7833 9346 7899 9349
rect 14046 9346 14106 9558
rect 30741 9555 30807 9558
rect 17401 9482 17467 9485
rect 36077 9482 36143 9485
rect 17401 9480 36143 9482
rect 17401 9424 17406 9480
rect 17462 9424 36082 9480
rect 36138 9424 36143 9480
rect 17401 9422 36143 9424
rect 17401 9419 17467 9422
rect 36077 9419 36143 9422
rect 7833 9344 14106 9346
rect 7833 9288 7838 9344
rect 7894 9288 14106 9344
rect 7833 9286 14106 9288
rect 24393 9346 24459 9349
rect 26509 9346 26575 9349
rect 24393 9344 26575 9346
rect 24393 9288 24398 9344
rect 24454 9288 26514 9344
rect 26570 9288 26575 9344
rect 24393 9286 26575 9288
rect 7833 9283 7899 9286
rect 24393 9283 24459 9286
rect 26509 9283 26575 9286
rect 36629 9346 36695 9349
rect 39520 9346 40000 9376
rect 36629 9344 40000 9346
rect 36629 9288 36634 9344
rect 36690 9288 40000 9344
rect 36629 9286 40000 9288
rect 36629 9283 36695 9286
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 39520 9256 40000 9286
rect 27610 9215 27930 9216
rect 4613 9210 4679 9213
rect 8293 9210 8359 9213
rect 4613 9208 8359 9210
rect 4613 9152 4618 9208
rect 4674 9152 8298 9208
rect 8354 9152 8359 9208
rect 4613 9150 8359 9152
rect 4613 9147 4679 9150
rect 8293 9147 8359 9150
rect 1485 9074 1551 9077
rect 3417 9074 3483 9077
rect 17861 9074 17927 9077
rect 25221 9074 25287 9077
rect 26325 9074 26391 9077
rect 1485 9072 26391 9074
rect 1485 9016 1490 9072
rect 1546 9016 3422 9072
rect 3478 9016 17866 9072
rect 17922 9016 25226 9072
rect 25282 9016 26330 9072
rect 26386 9016 26391 9072
rect 1485 9014 26391 9016
rect 1485 9011 1551 9014
rect 3417 9011 3483 9014
rect 17861 9011 17927 9014
rect 25221 9011 25287 9014
rect 26325 9011 26391 9014
rect 3877 8938 3943 8941
rect 8845 8938 8911 8941
rect 3877 8936 8911 8938
rect 3877 8880 3882 8936
rect 3938 8880 8850 8936
rect 8906 8880 8911 8936
rect 3877 8878 8911 8880
rect 3877 8875 3943 8878
rect 8845 8875 8911 8878
rect 14089 8938 14155 8941
rect 19793 8938 19859 8941
rect 14089 8936 19859 8938
rect 14089 8880 14094 8936
rect 14150 8880 19798 8936
rect 19854 8880 19859 8936
rect 14089 8878 19859 8880
rect 14089 8875 14155 8878
rect 19793 8875 19859 8878
rect 19977 8938 20043 8941
rect 22737 8938 22803 8941
rect 26969 8938 27035 8941
rect 19977 8936 27035 8938
rect 19977 8880 19982 8936
rect 20038 8880 22742 8936
rect 22798 8880 26974 8936
rect 27030 8880 27035 8936
rect 19977 8878 27035 8880
rect 19977 8875 20043 8878
rect 22737 8875 22803 8878
rect 26969 8875 27035 8878
rect 8201 8802 8267 8805
rect 8385 8802 8451 8805
rect 16941 8802 17007 8805
rect 8201 8800 17007 8802
rect 8201 8744 8206 8800
rect 8262 8744 8390 8800
rect 8446 8744 16946 8800
rect 17002 8744 17007 8800
rect 8201 8742 17007 8744
rect 8201 8739 8267 8742
rect 8385 8739 8451 8742
rect 16941 8739 17007 8742
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 0 8530 480 8560
rect 1577 8530 1643 8533
rect 0 8528 1643 8530
rect 0 8472 1582 8528
rect 1638 8472 1643 8528
rect 0 8470 1643 8472
rect 0 8440 480 8470
rect 1577 8467 1643 8470
rect 6729 8530 6795 8533
rect 9673 8530 9739 8533
rect 33961 8530 34027 8533
rect 6729 8528 9739 8530
rect 6729 8472 6734 8528
rect 6790 8472 9678 8528
rect 9734 8472 9739 8528
rect 6729 8470 9739 8472
rect 6729 8467 6795 8470
rect 9673 8467 9739 8470
rect 9814 8528 34027 8530
rect 9814 8472 33966 8528
rect 34022 8472 34027 8528
rect 9814 8470 34027 8472
rect 5165 8394 5231 8397
rect 7833 8394 7899 8397
rect 5165 8392 7899 8394
rect 5165 8336 5170 8392
rect 5226 8336 7838 8392
rect 7894 8336 7899 8392
rect 5165 8334 7899 8336
rect 5165 8331 5231 8334
rect 7833 8331 7899 8334
rect 9489 8394 9555 8397
rect 9814 8394 9874 8470
rect 33961 8467 34027 8470
rect 36629 8530 36695 8533
rect 39520 8530 40000 8560
rect 36629 8528 40000 8530
rect 36629 8472 36634 8528
rect 36690 8472 40000 8528
rect 36629 8470 40000 8472
rect 36629 8467 36695 8470
rect 39520 8440 40000 8470
rect 9489 8392 9874 8394
rect 9489 8336 9494 8392
rect 9550 8336 9874 8392
rect 9489 8334 9874 8336
rect 10777 8394 10843 8397
rect 12801 8394 12867 8397
rect 10777 8392 12867 8394
rect 10777 8336 10782 8392
rect 10838 8336 12806 8392
rect 12862 8336 12867 8392
rect 10777 8334 12867 8336
rect 9489 8331 9555 8334
rect 10777 8331 10843 8334
rect 12801 8331 12867 8334
rect 16021 8394 16087 8397
rect 21265 8394 21331 8397
rect 16021 8392 21331 8394
rect 16021 8336 16026 8392
rect 16082 8336 21270 8392
rect 21326 8336 21331 8392
rect 16021 8334 21331 8336
rect 16021 8331 16087 8334
rect 21265 8331 21331 8334
rect 21449 8394 21515 8397
rect 25773 8394 25839 8397
rect 30465 8394 30531 8397
rect 21449 8392 30531 8394
rect 21449 8336 21454 8392
rect 21510 8336 25778 8392
rect 25834 8336 30470 8392
rect 30526 8336 30531 8392
rect 21449 8334 30531 8336
rect 21449 8331 21515 8334
rect 25773 8331 25839 8334
rect 30465 8331 30531 8334
rect 31569 8394 31635 8397
rect 35249 8394 35315 8397
rect 35985 8394 36051 8397
rect 31569 8392 36051 8394
rect 31569 8336 31574 8392
rect 31630 8336 35254 8392
rect 35310 8336 35990 8392
rect 36046 8336 36051 8392
rect 31569 8334 36051 8336
rect 31569 8331 31635 8334
rect 35249 8331 35315 8334
rect 35985 8331 36051 8334
rect 5349 8258 5415 8261
rect 8753 8258 8819 8261
rect 5349 8256 8819 8258
rect 5349 8200 5354 8256
rect 5410 8200 8758 8256
rect 8814 8200 8819 8256
rect 5349 8198 8819 8200
rect 5349 8195 5415 8198
rect 8753 8195 8819 8198
rect 10961 8258 11027 8261
rect 11789 8258 11855 8261
rect 13445 8258 13511 8261
rect 10961 8256 13511 8258
rect 10961 8200 10966 8256
rect 11022 8200 11794 8256
rect 11850 8200 13450 8256
rect 13506 8200 13511 8256
rect 10961 8198 13511 8200
rect 10961 8195 11027 8198
rect 11789 8195 11855 8198
rect 13445 8195 13511 8198
rect 14733 8258 14799 8261
rect 17902 8258 17908 8260
rect 14733 8256 17908 8258
rect 14733 8200 14738 8256
rect 14794 8200 17908 8256
rect 14733 8198 17908 8200
rect 14733 8195 14799 8198
rect 17902 8196 17908 8198
rect 17972 8196 17978 8260
rect 19425 8258 19491 8261
rect 25221 8258 25287 8261
rect 26049 8258 26115 8261
rect 19425 8256 26115 8258
rect 19425 8200 19430 8256
rect 19486 8200 25226 8256
rect 25282 8200 26054 8256
rect 26110 8200 26115 8256
rect 19425 8198 26115 8200
rect 19425 8195 19491 8198
rect 25221 8195 25287 8198
rect 26049 8195 26115 8198
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 14736 8088 17970 8122
rect 18045 8088 18111 8091
rect 14736 8086 18111 8088
rect 14736 8062 18050 8086
rect 3785 7986 3851 7989
rect 11053 7986 11119 7989
rect 11329 7986 11395 7989
rect 3785 7984 11395 7986
rect 3785 7928 3790 7984
rect 3846 7928 11058 7984
rect 11114 7928 11334 7984
rect 11390 7928 11395 7984
rect 3785 7926 11395 7928
rect 3785 7923 3851 7926
rect 11053 7923 11119 7926
rect 11329 7923 11395 7926
rect 13813 7986 13879 7989
rect 14736 7986 14796 8062
rect 17910 8030 18050 8062
rect 18106 8030 18111 8086
rect 17910 8028 18111 8030
rect 18045 8025 18111 8028
rect 13813 7984 14796 7986
rect 13813 7928 13818 7984
rect 13874 7928 14796 7984
rect 13813 7926 14796 7928
rect 13813 7923 13879 7926
rect 5625 7850 5691 7853
rect 13813 7850 13879 7853
rect 16665 7850 16731 7853
rect 5625 7848 16731 7850
rect 5625 7792 5630 7848
rect 5686 7792 13818 7848
rect 13874 7792 16670 7848
rect 16726 7792 16731 7848
rect 5625 7790 16731 7792
rect 5625 7787 5691 7790
rect 13813 7787 13879 7790
rect 16665 7787 16731 7790
rect 19425 7850 19491 7853
rect 30557 7850 30623 7853
rect 19425 7848 30623 7850
rect 19425 7792 19430 7848
rect 19486 7792 30562 7848
rect 30618 7792 30623 7848
rect 19425 7790 30623 7792
rect 19425 7787 19491 7790
rect 30557 7787 30623 7790
rect 17902 7652 17908 7716
rect 17972 7714 17978 7716
rect 20805 7714 20871 7717
rect 17972 7712 20871 7714
rect 17972 7656 20810 7712
rect 20866 7656 20871 7712
rect 17972 7654 20871 7656
rect 17972 7652 17978 7654
rect 20805 7651 20871 7654
rect 7610 7648 7930 7649
rect 0 7578 480 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 3049 7578 3115 7581
rect 0 7576 3115 7578
rect 0 7520 3054 7576
rect 3110 7520 3115 7576
rect 0 7518 3115 7520
rect 0 7488 480 7518
rect 3049 7515 3115 7518
rect 15285 7578 15351 7581
rect 17677 7578 17743 7581
rect 15285 7576 17743 7578
rect 15285 7520 15290 7576
rect 15346 7520 17682 7576
rect 17738 7520 17743 7576
rect 15285 7518 17743 7520
rect 15285 7515 15351 7518
rect 17677 7515 17743 7518
rect 18781 7578 18847 7581
rect 19425 7578 19491 7581
rect 18781 7576 19491 7578
rect 18781 7520 18786 7576
rect 18842 7520 19430 7576
rect 19486 7520 19491 7576
rect 18781 7518 19491 7520
rect 18781 7515 18847 7518
rect 19425 7515 19491 7518
rect 26325 7578 26391 7581
rect 39520 7578 40000 7608
rect 26325 7576 34162 7578
rect 26325 7520 26330 7576
rect 26386 7520 34162 7576
rect 26325 7518 34162 7520
rect 26325 7515 26391 7518
rect 7281 7442 7347 7445
rect 9949 7442 10015 7445
rect 7281 7440 10015 7442
rect 7281 7384 7286 7440
rect 7342 7384 9954 7440
rect 10010 7384 10015 7440
rect 7281 7382 10015 7384
rect 7281 7379 7347 7382
rect 9949 7379 10015 7382
rect 11053 7442 11119 7445
rect 20161 7442 20227 7445
rect 11053 7440 20227 7442
rect 11053 7384 11058 7440
rect 11114 7384 20166 7440
rect 20222 7384 20227 7440
rect 11053 7382 20227 7384
rect 11053 7379 11119 7382
rect 20161 7379 20227 7382
rect 23933 7442 23999 7445
rect 31385 7442 31451 7445
rect 32857 7442 32923 7445
rect 23933 7440 32923 7442
rect 23933 7384 23938 7440
rect 23994 7384 31390 7440
rect 31446 7384 32862 7440
rect 32918 7384 32923 7440
rect 23933 7382 32923 7384
rect 34102 7442 34162 7518
rect 34838 7518 40000 7578
rect 34838 7442 34898 7518
rect 39520 7488 40000 7518
rect 34102 7382 34898 7442
rect 23933 7379 23999 7382
rect 31385 7379 31451 7382
rect 32857 7379 32923 7382
rect 2221 7306 2287 7309
rect 12617 7306 12683 7309
rect 2221 7304 12683 7306
rect 2221 7248 2226 7304
rect 2282 7248 12622 7304
rect 12678 7248 12683 7304
rect 2221 7246 12683 7248
rect 2221 7243 2287 7246
rect 12617 7243 12683 7246
rect 23289 7306 23355 7309
rect 30557 7306 30623 7309
rect 23289 7304 30623 7306
rect 23289 7248 23294 7304
rect 23350 7248 30562 7304
rect 30618 7248 30623 7304
rect 23289 7246 30623 7248
rect 23289 7243 23355 7246
rect 30557 7243 30623 7246
rect 8753 7170 8819 7173
rect 12709 7170 12775 7173
rect 8753 7168 12775 7170
rect 8753 7112 8758 7168
rect 8814 7112 12714 7168
rect 12770 7112 12775 7168
rect 8753 7110 12775 7112
rect 8753 7107 8819 7110
rect 12709 7107 12775 7110
rect 33225 7170 33291 7173
rect 34789 7170 34855 7173
rect 33225 7168 34855 7170
rect 33225 7112 33230 7168
rect 33286 7112 34794 7168
rect 34850 7112 34855 7168
rect 33225 7110 34855 7112
rect 33225 7107 33291 7110
rect 34789 7107 34855 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 5717 7034 5783 7037
rect 10501 7034 10567 7037
rect 5717 7032 10567 7034
rect 5717 6976 5722 7032
rect 5778 6976 10506 7032
rect 10562 6976 10567 7032
rect 5717 6974 10567 6976
rect 5717 6971 5783 6974
rect 10501 6971 10567 6974
rect 16573 7034 16639 7037
rect 19241 7034 19307 7037
rect 28165 7034 28231 7037
rect 16573 7032 19307 7034
rect 16573 6976 16578 7032
rect 16634 6976 19246 7032
rect 19302 6976 19307 7032
rect 16573 6974 19307 6976
rect 16573 6971 16639 6974
rect 19241 6971 19307 6974
rect 28030 7032 28231 7034
rect 28030 6976 28170 7032
rect 28226 6976 28231 7032
rect 28030 6974 28231 6976
rect 8201 6898 8267 6901
rect 2684 6896 8267 6898
rect 2684 6840 8206 6896
rect 8262 6840 8267 6896
rect 2684 6838 8267 6840
rect 0 6626 480 6656
rect 2684 6626 2744 6838
rect 8201 6835 8267 6838
rect 24025 6898 24091 6901
rect 28030 6898 28090 6974
rect 28165 6971 28231 6974
rect 24025 6896 28090 6898
rect 24025 6840 24030 6896
rect 24086 6840 28090 6896
rect 24025 6838 28090 6840
rect 33777 6898 33843 6901
rect 33777 6896 36738 6898
rect 33777 6840 33782 6896
rect 33838 6840 36738 6896
rect 33777 6838 36738 6840
rect 24025 6835 24091 6838
rect 33777 6835 33843 6838
rect 18689 6762 18755 6765
rect 20713 6762 20779 6765
rect 18689 6760 20779 6762
rect 18689 6704 18694 6760
rect 18750 6704 20718 6760
rect 20774 6704 20779 6760
rect 18689 6702 20779 6704
rect 18689 6699 18755 6702
rect 20713 6699 20779 6702
rect 32213 6762 32279 6765
rect 36445 6762 36511 6765
rect 32213 6760 36511 6762
rect 32213 6704 32218 6760
rect 32274 6704 36450 6760
rect 36506 6704 36511 6760
rect 32213 6702 36511 6704
rect 32213 6699 32279 6702
rect 36445 6699 36511 6702
rect 0 6566 2744 6626
rect 36678 6626 36738 6838
rect 39520 6626 40000 6656
rect 36678 6566 40000 6626
rect 0 6536 480 6566
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 39520 6536 40000 6566
rect 34277 6495 34597 6496
rect 10685 6490 10751 6493
rect 14917 6490 14983 6493
rect 16205 6490 16271 6493
rect 16573 6490 16639 6493
rect 10685 6488 16639 6490
rect 10685 6432 10690 6488
rect 10746 6432 14922 6488
rect 14978 6432 16210 6488
rect 16266 6432 16578 6488
rect 16634 6432 16639 6488
rect 10685 6430 16639 6432
rect 10685 6427 10751 6430
rect 14917 6427 14983 6430
rect 16205 6427 16271 6430
rect 16573 6427 16639 6430
rect 23381 6490 23447 6493
rect 27337 6490 27403 6493
rect 23381 6488 27403 6490
rect 23381 6432 23386 6488
rect 23442 6432 27342 6488
rect 27398 6432 27403 6488
rect 23381 6430 27403 6432
rect 23381 6427 23447 6430
rect 27337 6427 27403 6430
rect 30833 6490 30899 6493
rect 33501 6490 33567 6493
rect 30833 6488 33567 6490
rect 30833 6432 30838 6488
rect 30894 6432 33506 6488
rect 33562 6432 33567 6488
rect 30833 6430 33567 6432
rect 30833 6427 30899 6430
rect 33501 6427 33567 6430
rect 5901 6354 5967 6357
rect 8661 6354 8727 6357
rect 14181 6354 14247 6357
rect 17493 6354 17559 6357
rect 5901 6352 17559 6354
rect 5901 6296 5906 6352
rect 5962 6296 8666 6352
rect 8722 6296 14186 6352
rect 14242 6296 17498 6352
rect 17554 6296 17559 6352
rect 5901 6294 17559 6296
rect 5901 6291 5967 6294
rect 8661 6291 8727 6294
rect 14181 6291 14247 6294
rect 17493 6291 17559 6294
rect 24577 6354 24643 6357
rect 27153 6354 27219 6357
rect 24577 6352 27219 6354
rect 24577 6296 24582 6352
rect 24638 6296 27158 6352
rect 27214 6296 27219 6352
rect 24577 6294 27219 6296
rect 24577 6291 24643 6294
rect 27153 6291 27219 6294
rect 10869 6218 10935 6221
rect 12893 6218 12959 6221
rect 10869 6216 12959 6218
rect 10869 6160 10874 6216
rect 10930 6160 12898 6216
rect 12954 6160 12959 6216
rect 10869 6158 12959 6160
rect 10869 6155 10935 6158
rect 12893 6155 12959 6158
rect 13905 6218 13971 6221
rect 15193 6218 15259 6221
rect 13905 6216 15259 6218
rect 13905 6160 13910 6216
rect 13966 6160 15198 6216
rect 15254 6160 15259 6216
rect 13905 6158 15259 6160
rect 13905 6155 13971 6158
rect 15193 6155 15259 6158
rect 17861 6218 17927 6221
rect 23473 6218 23539 6221
rect 33409 6218 33475 6221
rect 17861 6216 23539 6218
rect 17861 6160 17866 6216
rect 17922 6160 23478 6216
rect 23534 6160 23539 6216
rect 17861 6158 23539 6160
rect 17861 6155 17927 6158
rect 23473 6155 23539 6158
rect 26190 6216 33475 6218
rect 26190 6160 33414 6216
rect 33470 6160 33475 6216
rect 26190 6158 33475 6160
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 9581 5946 9647 5949
rect 17677 5946 17743 5949
rect 19885 5946 19951 5949
rect 23105 5946 23171 5949
rect 9581 5944 12312 5946
rect 9581 5888 9586 5944
rect 9642 5912 12312 5944
rect 12390 5912 13140 5946
rect 9642 5888 13140 5912
rect 9581 5886 13140 5888
rect 9581 5883 9647 5886
rect 12252 5852 12450 5886
rect 0 5810 480 5840
rect 4797 5810 4863 5813
rect 9121 5810 9187 5813
rect 0 5808 9187 5810
rect 0 5752 4802 5808
rect 4858 5752 9126 5808
rect 9182 5752 9187 5808
rect 0 5750 9187 5752
rect 0 5720 480 5750
rect 4797 5747 4863 5750
rect 9121 5747 9187 5750
rect 9581 5810 9647 5813
rect 10685 5810 10751 5813
rect 9581 5808 10751 5810
rect 9581 5752 9586 5808
rect 9642 5752 10690 5808
rect 10746 5752 10751 5808
rect 9581 5750 10751 5752
rect 13080 5810 13140 5886
rect 17677 5944 23171 5946
rect 17677 5888 17682 5944
rect 17738 5888 19890 5944
rect 19946 5888 23110 5944
rect 23166 5888 23171 5944
rect 17677 5886 23171 5888
rect 17677 5883 17743 5886
rect 19885 5883 19951 5886
rect 23105 5883 23171 5886
rect 26190 5810 26250 6158
rect 33409 6155 33475 6158
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 13080 5750 26250 5810
rect 26325 5810 26391 5813
rect 29085 5810 29151 5813
rect 26325 5808 29151 5810
rect 26325 5752 26330 5808
rect 26386 5752 29090 5808
rect 29146 5752 29151 5808
rect 26325 5750 29151 5752
rect 9581 5747 9647 5750
rect 10685 5747 10751 5750
rect 26325 5747 26391 5750
rect 29085 5747 29151 5750
rect 34789 5810 34855 5813
rect 39520 5810 40000 5840
rect 34789 5808 40000 5810
rect 34789 5752 34794 5808
rect 34850 5752 40000 5808
rect 34789 5750 40000 5752
rect 34789 5747 34855 5750
rect 39520 5720 40000 5750
rect 10869 5674 10935 5677
rect 6686 5672 10935 5674
rect 6686 5616 10874 5672
rect 10930 5616 10935 5672
rect 6686 5614 10935 5616
rect 2957 5538 3023 5541
rect 5993 5538 6059 5541
rect 6686 5538 6746 5614
rect 10869 5611 10935 5614
rect 12157 5674 12223 5677
rect 14825 5674 14891 5677
rect 12157 5672 14891 5674
rect 12157 5616 12162 5672
rect 12218 5616 14830 5672
rect 14886 5616 14891 5672
rect 12157 5614 14891 5616
rect 12157 5611 12223 5614
rect 14825 5611 14891 5614
rect 24117 5674 24183 5677
rect 26877 5674 26943 5677
rect 29177 5674 29243 5677
rect 24117 5672 29243 5674
rect 24117 5616 24122 5672
rect 24178 5616 26882 5672
rect 26938 5616 29182 5672
rect 29238 5616 29243 5672
rect 24117 5614 29243 5616
rect 24117 5611 24183 5614
rect 26877 5611 26943 5614
rect 29177 5611 29243 5614
rect 2957 5536 6746 5538
rect 2957 5480 2962 5536
rect 3018 5480 5998 5536
rect 6054 5480 6746 5536
rect 2957 5478 6746 5480
rect 10501 5538 10567 5541
rect 11513 5538 11579 5541
rect 10501 5536 11579 5538
rect 10501 5480 10506 5536
rect 10562 5480 11518 5536
rect 11574 5480 11579 5536
rect 10501 5478 11579 5480
rect 2957 5475 3023 5478
rect 5993 5475 6059 5478
rect 10501 5475 10567 5478
rect 11513 5475 11579 5478
rect 12249 5538 12315 5541
rect 14181 5538 14247 5541
rect 12249 5536 14247 5538
rect 12249 5480 12254 5536
rect 12310 5480 14186 5536
rect 14242 5480 14247 5536
rect 12249 5478 14247 5480
rect 12249 5475 12315 5478
rect 14181 5475 14247 5478
rect 27061 5538 27127 5541
rect 30373 5538 30439 5541
rect 27061 5536 30439 5538
rect 27061 5480 27066 5536
rect 27122 5480 30378 5536
rect 30434 5480 30439 5536
rect 27061 5478 30439 5480
rect 27061 5475 27127 5478
rect 30373 5475 30439 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 9121 5402 9187 5405
rect 14089 5402 14155 5405
rect 9121 5400 14155 5402
rect 9121 5344 9126 5400
rect 9182 5344 14094 5400
rect 14150 5344 14155 5400
rect 9121 5342 14155 5344
rect 9121 5339 9187 5342
rect 14089 5339 14155 5342
rect 4889 5266 4955 5269
rect 12157 5266 12223 5269
rect 4889 5264 12223 5266
rect 4889 5208 4894 5264
rect 4950 5208 12162 5264
rect 12218 5208 12223 5264
rect 4889 5206 12223 5208
rect 4889 5203 4955 5206
rect 12157 5203 12223 5206
rect 13077 5266 13143 5269
rect 21265 5266 21331 5269
rect 31293 5266 31359 5269
rect 13077 5264 31359 5266
rect 13077 5208 13082 5264
rect 13138 5208 21270 5264
rect 21326 5208 31298 5264
rect 31354 5208 31359 5264
rect 13077 5206 31359 5208
rect 13077 5203 13143 5206
rect 21265 5203 21331 5206
rect 31293 5203 31359 5206
rect 23473 5130 23539 5133
rect 32213 5130 32279 5133
rect 23473 5128 32279 5130
rect 23473 5072 23478 5128
rect 23534 5072 32218 5128
rect 32274 5072 32279 5128
rect 23473 5070 32279 5072
rect 23473 5067 23539 5070
rect 32213 5067 32279 5070
rect 14733 4994 14799 4997
rect 17769 4994 17835 4997
rect 24945 4994 25011 4997
rect 14733 4992 25011 4994
rect 14733 4936 14738 4992
rect 14794 4936 17774 4992
rect 17830 4936 24950 4992
rect 25006 4936 25011 4992
rect 14733 4934 25011 4936
rect 14733 4931 14799 4934
rect 17769 4931 17835 4934
rect 24945 4931 25011 4934
rect 31753 4994 31819 4997
rect 34697 4994 34763 4997
rect 31753 4992 34763 4994
rect 31753 4936 31758 4992
rect 31814 4936 34702 4992
rect 34758 4936 34763 4992
rect 31753 4934 34763 4936
rect 31753 4931 31819 4934
rect 34697 4931 34763 4934
rect 14277 4928 14597 4929
rect 0 4858 480 4888
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 13537 4858 13603 4861
rect 0 4856 13603 4858
rect 0 4800 13542 4856
rect 13598 4800 13603 4856
rect 0 4798 13603 4800
rect 0 4768 480 4798
rect 13537 4795 13603 4798
rect 18413 4858 18479 4861
rect 22737 4858 22803 4861
rect 18413 4856 22803 4858
rect 18413 4800 18418 4856
rect 18474 4800 22742 4856
rect 22798 4800 22803 4856
rect 18413 4798 22803 4800
rect 18413 4795 18479 4798
rect 22737 4795 22803 4798
rect 35433 4858 35499 4861
rect 39520 4858 40000 4888
rect 35433 4856 40000 4858
rect 35433 4800 35438 4856
rect 35494 4800 40000 4856
rect 35433 4798 40000 4800
rect 35433 4795 35499 4798
rect 39520 4768 40000 4798
rect 12617 4722 12683 4725
rect 19977 4722 20043 4725
rect 12617 4720 20043 4722
rect 12617 4664 12622 4720
rect 12678 4664 19982 4720
rect 20038 4664 20043 4720
rect 12617 4662 20043 4664
rect 12617 4659 12683 4662
rect 19977 4659 20043 4662
rect 27337 4722 27403 4725
rect 31569 4722 31635 4725
rect 27337 4720 31635 4722
rect 27337 4664 27342 4720
rect 27398 4664 31574 4720
rect 31630 4664 31635 4720
rect 27337 4662 31635 4664
rect 27337 4659 27403 4662
rect 31569 4659 31635 4662
rect 6269 4586 6335 4589
rect 17125 4586 17191 4589
rect 6269 4584 17191 4586
rect 6269 4528 6274 4584
rect 6330 4528 17130 4584
rect 17186 4528 17191 4584
rect 6269 4526 17191 4528
rect 6269 4523 6335 4526
rect 17125 4523 17191 4526
rect 15009 4450 15075 4453
rect 17033 4450 17099 4453
rect 15009 4448 17099 4450
rect 15009 4392 15014 4448
rect 15070 4392 17038 4448
rect 17094 4392 17099 4448
rect 15009 4390 17099 4392
rect 15009 4387 15075 4390
rect 17033 4387 17099 4390
rect 23565 4450 23631 4453
rect 28942 4450 28948 4452
rect 23565 4448 28948 4450
rect 23565 4392 23570 4448
rect 23626 4392 28948 4448
rect 23565 4390 28948 4392
rect 23565 4387 23631 4390
rect 28942 4388 28948 4390
rect 29012 4388 29018 4452
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 30189 4314 30255 4317
rect 23062 4312 30255 4314
rect 23062 4256 30194 4312
rect 30250 4256 30255 4312
rect 23062 4254 30255 4256
rect 5717 4178 5783 4181
rect 10133 4178 10199 4181
rect 5717 4176 10199 4178
rect 5717 4120 5722 4176
rect 5778 4120 10138 4176
rect 10194 4120 10199 4176
rect 5717 4118 10199 4120
rect 5717 4115 5783 4118
rect 10133 4115 10199 4118
rect 11513 4178 11579 4181
rect 23062 4178 23122 4254
rect 30189 4251 30255 4254
rect 11513 4176 23122 4178
rect 11513 4120 11518 4176
rect 11574 4120 23122 4176
rect 11513 4118 23122 4120
rect 23197 4178 23263 4181
rect 27981 4178 28047 4181
rect 23197 4176 28047 4178
rect 23197 4120 23202 4176
rect 23258 4120 27986 4176
rect 28042 4120 28047 4176
rect 23197 4118 28047 4120
rect 11513 4115 11579 4118
rect 23197 4115 23263 4118
rect 27981 4115 28047 4118
rect 0 4042 480 4072
rect 2865 4042 2931 4045
rect 0 4040 2931 4042
rect 0 3984 2870 4040
rect 2926 3984 2931 4040
rect 0 3982 2931 3984
rect 0 3952 480 3982
rect 2865 3979 2931 3982
rect 3325 4042 3391 4045
rect 3969 4042 4035 4045
rect 5993 4042 6059 4045
rect 6637 4042 6703 4045
rect 3325 4040 6703 4042
rect 3325 3984 3330 4040
rect 3386 3984 3974 4040
rect 4030 3984 5998 4040
rect 6054 3984 6642 4040
rect 6698 3984 6703 4040
rect 3325 3982 6703 3984
rect 3325 3979 3391 3982
rect 3969 3979 4035 3982
rect 5993 3979 6059 3982
rect 6637 3979 6703 3982
rect 7373 4042 7439 4045
rect 9949 4042 10015 4045
rect 7373 4040 10015 4042
rect 7373 3984 7378 4040
rect 7434 3984 9954 4040
rect 10010 3984 10015 4040
rect 7373 3982 10015 3984
rect 7373 3979 7439 3982
rect 9949 3979 10015 3982
rect 25497 4042 25563 4045
rect 27797 4042 27863 4045
rect 25497 4040 27863 4042
rect 25497 3984 25502 4040
rect 25558 3984 27802 4040
rect 27858 3984 27863 4040
rect 25497 3982 27863 3984
rect 25497 3979 25563 3982
rect 27797 3979 27863 3982
rect 29821 4042 29887 4045
rect 39520 4042 40000 4072
rect 29821 4040 40000 4042
rect 29821 3984 29826 4040
rect 29882 3984 40000 4040
rect 29821 3982 40000 3984
rect 29821 3979 29887 3982
rect 39520 3952 40000 3982
rect 2957 3906 3023 3909
rect 5901 3906 5967 3909
rect 8753 3906 8819 3909
rect 9581 3906 9647 3909
rect 2957 3904 9647 3906
rect 2957 3848 2962 3904
rect 3018 3848 5906 3904
rect 5962 3848 8758 3904
rect 8814 3848 9586 3904
rect 9642 3848 9647 3904
rect 2957 3846 9647 3848
rect 2957 3843 3023 3846
rect 5901 3843 5967 3846
rect 8753 3843 8819 3846
rect 9581 3843 9647 3846
rect 19885 3906 19951 3909
rect 27061 3906 27127 3909
rect 19885 3904 27127 3906
rect 19885 3848 19890 3904
rect 19946 3848 27066 3904
rect 27122 3848 27127 3904
rect 19885 3846 27127 3848
rect 19885 3843 19951 3846
rect 27061 3843 27127 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 3693 3770 3759 3773
rect 6545 3770 6611 3773
rect 9213 3770 9279 3773
rect 12157 3772 12223 3773
rect 12157 3770 12204 3772
rect 3693 3768 9279 3770
rect 3693 3712 3698 3768
rect 3754 3712 6550 3768
rect 6606 3712 9218 3768
rect 9274 3712 9279 3768
rect 3693 3710 9279 3712
rect 12112 3768 12204 3770
rect 12112 3712 12162 3768
rect 12112 3710 12204 3712
rect 3693 3707 3759 3710
rect 6545 3707 6611 3710
rect 9213 3707 9279 3710
rect 12157 3708 12204 3710
rect 12268 3708 12274 3772
rect 15837 3770 15903 3773
rect 20897 3770 20963 3773
rect 26417 3772 26483 3773
rect 15837 3768 20963 3770
rect 15837 3712 15842 3768
rect 15898 3712 20902 3768
rect 20958 3712 20963 3768
rect 15837 3710 20963 3712
rect 12157 3707 12223 3708
rect 15837 3707 15903 3710
rect 20897 3707 20963 3710
rect 26366 3708 26372 3772
rect 26436 3770 26483 3772
rect 26436 3768 26528 3770
rect 26478 3712 26528 3768
rect 26436 3710 26528 3712
rect 26436 3708 26483 3710
rect 26417 3707 26483 3708
rect 6361 3634 6427 3637
rect 8845 3634 8911 3637
rect 6361 3632 8911 3634
rect 6361 3576 6366 3632
rect 6422 3576 8850 3632
rect 8906 3576 8911 3632
rect 6361 3574 8911 3576
rect 6361 3571 6427 3574
rect 8845 3571 8911 3574
rect 9029 3634 9095 3637
rect 12249 3634 12315 3637
rect 21081 3634 21147 3637
rect 9029 3632 21147 3634
rect 9029 3576 9034 3632
rect 9090 3576 12254 3632
rect 12310 3576 21086 3632
rect 21142 3576 21147 3632
rect 9029 3574 21147 3576
rect 9029 3571 9095 3574
rect 12249 3571 12315 3574
rect 21081 3571 21147 3574
rect 22645 3634 22711 3637
rect 30465 3634 30531 3637
rect 22645 3632 30531 3634
rect 22645 3576 22650 3632
rect 22706 3576 30470 3632
rect 30526 3576 30531 3632
rect 22645 3574 30531 3576
rect 22645 3571 22711 3574
rect 30465 3571 30531 3574
rect 1945 3498 2011 3501
rect 4429 3498 4495 3501
rect 6177 3498 6243 3501
rect 10133 3498 10199 3501
rect 1945 3496 10199 3498
rect 1945 3440 1950 3496
rect 2006 3440 4434 3496
rect 4490 3440 6182 3496
rect 6238 3440 10138 3496
rect 10194 3440 10199 3496
rect 1945 3438 10199 3440
rect 1945 3435 2011 3438
rect 4429 3435 4495 3438
rect 6177 3435 6243 3438
rect 10133 3435 10199 3438
rect 14365 3498 14431 3501
rect 19149 3498 19215 3501
rect 14365 3496 19215 3498
rect 14365 3440 14370 3496
rect 14426 3440 19154 3496
rect 19210 3440 19215 3496
rect 14365 3438 19215 3440
rect 14365 3435 14431 3438
rect 19149 3435 19215 3438
rect 26969 3498 27035 3501
rect 29545 3498 29611 3501
rect 26969 3496 29611 3498
rect 26969 3440 26974 3496
rect 27030 3440 29550 3496
rect 29606 3440 29611 3496
rect 26969 3438 29611 3440
rect 26969 3435 27035 3438
rect 29545 3435 29611 3438
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 23841 3226 23907 3229
rect 27613 3226 27679 3229
rect 23841 3224 27679 3226
rect 23841 3168 23846 3224
rect 23902 3168 27618 3224
rect 27674 3168 27679 3224
rect 23841 3166 27679 3168
rect 23841 3163 23907 3166
rect 27613 3163 27679 3166
rect 28942 3164 28948 3228
rect 29012 3226 29018 3228
rect 29012 3166 30482 3226
rect 29012 3164 29018 3166
rect 0 3090 480 3120
rect 3785 3090 3851 3093
rect 0 3088 3851 3090
rect 0 3032 3790 3088
rect 3846 3032 3851 3088
rect 0 3030 3851 3032
rect 0 3000 480 3030
rect 3785 3027 3851 3030
rect 4245 3090 4311 3093
rect 4705 3090 4771 3093
rect 14181 3090 14247 3093
rect 14774 3090 14780 3092
rect 4245 3088 14780 3090
rect 4245 3032 4250 3088
rect 4306 3032 4710 3088
rect 4766 3032 14186 3088
rect 14242 3032 14780 3088
rect 4245 3030 14780 3032
rect 4245 3027 4311 3030
rect 4705 3027 4771 3030
rect 14181 3027 14247 3030
rect 14774 3028 14780 3030
rect 14844 3028 14850 3092
rect 18781 3090 18847 3093
rect 30281 3090 30347 3093
rect 18781 3088 30347 3090
rect 18781 3032 18786 3088
rect 18842 3032 30286 3088
rect 30342 3032 30347 3088
rect 18781 3030 30347 3032
rect 30422 3090 30482 3166
rect 39520 3090 40000 3120
rect 30422 3030 40000 3090
rect 18781 3027 18847 3030
rect 30281 3027 30347 3030
rect 39520 3000 40000 3030
rect 14641 2954 14707 2957
rect 19333 2954 19399 2957
rect 22553 2956 22619 2957
rect 22502 2954 22508 2956
rect 14641 2952 19399 2954
rect 14641 2896 14646 2952
rect 14702 2896 19338 2952
rect 19394 2896 19399 2952
rect 14641 2894 19399 2896
rect 22462 2894 22508 2954
rect 22572 2952 22619 2956
rect 22614 2896 22619 2952
rect 14641 2891 14707 2894
rect 19333 2891 19399 2894
rect 22502 2892 22508 2894
rect 22572 2892 22619 2896
rect 22553 2891 22619 2892
rect 27245 2954 27311 2957
rect 35801 2954 35867 2957
rect 27245 2952 35867 2954
rect 27245 2896 27250 2952
rect 27306 2896 35806 2952
rect 35862 2896 35867 2952
rect 27245 2894 35867 2896
rect 27245 2891 27311 2894
rect 35801 2891 35867 2894
rect 19149 2818 19215 2821
rect 19517 2818 19583 2821
rect 21633 2818 21699 2821
rect 19149 2816 21699 2818
rect 19149 2760 19154 2816
rect 19210 2760 19522 2816
rect 19578 2760 21638 2816
rect 21694 2760 21699 2816
rect 19149 2758 21699 2760
rect 19149 2755 19215 2758
rect 19517 2755 19583 2758
rect 21633 2755 21699 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 4889 2682 4955 2685
rect 8845 2682 8911 2685
rect 26325 2682 26391 2685
rect 4889 2680 8911 2682
rect 4889 2624 4894 2680
rect 4950 2624 8850 2680
rect 8906 2624 8911 2680
rect 4889 2622 8911 2624
rect 4889 2619 4955 2622
rect 8845 2619 8911 2622
rect 15150 2680 26391 2682
rect 15150 2624 26330 2680
rect 26386 2624 26391 2680
rect 15150 2622 26391 2624
rect 13353 2546 13419 2549
rect 15150 2546 15210 2622
rect 26325 2619 26391 2622
rect 33961 2682 34027 2685
rect 33961 2680 37842 2682
rect 33961 2624 33966 2680
rect 34022 2624 37842 2680
rect 33961 2622 37842 2624
rect 33961 2619 34027 2622
rect 13353 2544 15210 2546
rect 13353 2488 13358 2544
rect 13414 2488 15210 2544
rect 13353 2486 15210 2488
rect 20253 2546 20319 2549
rect 22461 2546 22527 2549
rect 20253 2544 22527 2546
rect 20253 2488 20258 2544
rect 20314 2488 22466 2544
rect 22522 2488 22527 2544
rect 20253 2486 22527 2488
rect 13353 2483 13419 2486
rect 20253 2483 20319 2486
rect 22461 2483 22527 2486
rect 24761 2546 24827 2549
rect 27889 2546 27955 2549
rect 35985 2546 36051 2549
rect 24761 2544 27955 2546
rect 24761 2488 24766 2544
rect 24822 2488 27894 2544
rect 27950 2488 27955 2544
rect 24761 2486 27955 2488
rect 24761 2483 24827 2486
rect 27889 2483 27955 2486
rect 28030 2544 36051 2546
rect 28030 2488 35990 2544
rect 36046 2488 36051 2544
rect 28030 2486 36051 2488
rect 1669 2410 1735 2413
rect 15193 2410 15259 2413
rect 1669 2408 15259 2410
rect 1669 2352 1674 2408
rect 1730 2352 15198 2408
rect 15254 2352 15259 2408
rect 1669 2350 15259 2352
rect 1669 2347 1735 2350
rect 15193 2347 15259 2350
rect 21357 2410 21423 2413
rect 26233 2410 26299 2413
rect 21357 2408 26299 2410
rect 21357 2352 21362 2408
rect 21418 2352 26238 2408
rect 26294 2352 26299 2408
rect 21357 2350 26299 2352
rect 21357 2347 21423 2350
rect 26233 2347 26299 2350
rect 0 2274 480 2304
rect 2221 2274 2287 2277
rect 0 2272 2287 2274
rect 0 2216 2226 2272
rect 2282 2216 2287 2272
rect 0 2214 2287 2216
rect 0 2184 480 2214
rect 2221 2211 2287 2214
rect 22461 2274 22527 2277
rect 26509 2274 26575 2277
rect 22461 2272 26575 2274
rect 22461 2216 22466 2272
rect 22522 2216 26514 2272
rect 26570 2216 26575 2272
rect 22461 2214 26575 2216
rect 22461 2211 22527 2214
rect 26509 2211 26575 2214
rect 27429 2274 27495 2277
rect 28030 2274 28090 2486
rect 35985 2483 36051 2486
rect 27429 2272 28090 2274
rect 27429 2216 27434 2272
rect 27490 2216 28090 2272
rect 27429 2214 28090 2216
rect 37782 2274 37842 2622
rect 39520 2274 40000 2304
rect 37782 2214 40000 2274
rect 27429 2211 27495 2214
rect 7610 2208 7930 2209
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 39520 2184 40000 2214
rect 34277 2143 34597 2144
rect 4153 2002 4219 2005
rect 12893 2002 12959 2005
rect 4153 2000 12959 2002
rect 4153 1944 4158 2000
rect 4214 1944 12898 2000
rect 12954 1944 12959 2000
rect 4153 1942 12959 1944
rect 4153 1939 4219 1942
rect 12893 1939 12959 1942
rect 11973 1866 12039 1869
rect 20805 1866 20871 1869
rect 11973 1864 20871 1866
rect 11973 1808 11978 1864
rect 12034 1808 20810 1864
rect 20866 1808 20871 1864
rect 11973 1806 20871 1808
rect 11973 1803 12039 1806
rect 20805 1803 20871 1806
rect 28901 1594 28967 1597
rect 34973 1594 35039 1597
rect 28901 1592 35039 1594
rect 28901 1536 28906 1592
rect 28962 1536 34978 1592
rect 35034 1536 35039 1592
rect 28901 1534 35039 1536
rect 28901 1531 28967 1534
rect 34973 1531 35039 1534
rect 31661 1458 31727 1461
rect 38285 1458 38351 1461
rect 31661 1456 38351 1458
rect 31661 1400 31666 1456
rect 31722 1400 38290 1456
rect 38346 1400 38351 1456
rect 31661 1398 38351 1400
rect 31661 1395 31727 1398
rect 38285 1395 38351 1398
rect 0 1322 480 1352
rect 4153 1322 4219 1325
rect 0 1320 4219 1322
rect 0 1264 4158 1320
rect 4214 1264 4219 1320
rect 0 1262 4219 1264
rect 0 1232 480 1262
rect 4153 1259 4219 1262
rect 35801 1322 35867 1325
rect 39520 1322 40000 1352
rect 35801 1320 40000 1322
rect 35801 1264 35806 1320
rect 35862 1264 40000 1320
rect 35801 1262 40000 1264
rect 35801 1259 35867 1262
rect 39520 1232 40000 1262
rect 0 506 480 536
rect 4245 506 4311 509
rect 0 504 4311 506
rect 0 448 4250 504
rect 4306 448 4311 504
rect 0 446 4311 448
rect 0 416 480 446
rect 4245 443 4311 446
rect 34697 506 34763 509
rect 39520 506 40000 536
rect 34697 504 40000 506
rect 34697 448 34702 504
rect 34758 448 40000 504
rect 34697 446 40000 448
rect 34697 443 34763 446
rect 39520 416 40000 446
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 28948 10916 29012 10980
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 28948 10644 29012 10708
rect 28948 10372 29012 10436
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 28948 9692 29012 9756
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 17908 8196 17972 8260
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 17908 7652 17972 7716
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 28948 4388 29012 4452
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 12204 3768 12268 3772
rect 12204 3712 12218 3768
rect 12218 3712 12268 3768
rect 12204 3708 12268 3712
rect 26372 3768 26436 3772
rect 26372 3712 26422 3768
rect 26422 3712 26436 3768
rect 26372 3708 26436 3712
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 28948 3164 29012 3228
rect 14780 3028 14844 3092
rect 22508 2952 22572 2956
rect 22508 2896 22558 2952
rect 22558 2896 22572 2952
rect 22508 2892 22572 2896
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 17907 8260 17973 8261
rect 17907 8196 17908 8260
rect 17972 8196 17973 8260
rect 17907 8195 17973 8196
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 17910 7717 17970 8195
rect 17907 7716 17973 7717
rect 17907 7652 17908 7716
rect 17972 7652 17973 7716
rect 17907 7651 17973 7652
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 2752 14597 3776
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 28947 10980 29013 10981
rect 28947 10916 28948 10980
rect 29012 10916 29013 10980
rect 28947 10915 29013 10916
rect 28950 10709 29010 10915
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 28947 10708 29013 10709
rect 28947 10644 28948 10708
rect 29012 10644 29013 10708
rect 28947 10643 29013 10644
rect 28947 10436 29013 10437
rect 28947 10372 28948 10436
rect 29012 10372 29013 10436
rect 28947 10371 29013 10372
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 28950 9757 29010 10371
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 28947 9756 29013 9757
rect 28947 9692 28948 9756
rect 29012 9692 29013 9756
rect 28947 9691 29013 9692
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 28947 4452 29013 4453
rect 28947 4388 28948 4452
rect 29012 4388 29013 4452
rect 28947 4387 29013 4388
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 2208 21264 3232
rect 22507 2892 22508 2942
rect 22572 2892 22573 2942
rect 22507 2891 22573 2892
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 2752 27930 3776
rect 28950 3229 29010 4387
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 28947 3228 29013 3229
rect 28947 3164 28948 3228
rect 29012 3164 29013 3228
rect 28947 3163 29013 3164
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
<< via4 >>
rect 12118 3772 12354 3858
rect 12118 3708 12204 3772
rect 12204 3708 12268 3772
rect 12268 3708 12354 3772
rect 12118 3622 12354 3708
rect 26286 3772 26522 3858
rect 26286 3708 26372 3772
rect 26372 3708 26436 3772
rect 26436 3708 26522 3772
rect 26286 3622 26522 3708
rect 14694 3092 14930 3178
rect 14694 3028 14780 3092
rect 14780 3028 14844 3092
rect 14844 3028 14930 3092
rect 14694 2942 14930 3028
rect 22422 2956 22658 3178
rect 22422 2942 22508 2956
rect 22508 2942 22572 2956
rect 22572 2942 22658 2956
<< metal5 >>
rect 12076 3858 26564 3900
rect 12076 3622 12118 3858
rect 12354 3622 26286 3858
rect 26522 3622 26564 3858
rect 12076 3580 26564 3622
rect 14652 3178 22700 3220
rect 14652 2942 14694 3178
rect 14930 2942 22422 3178
rect 22658 2942 22700 3178
rect 14652 2900 22700 2942
use scs8hd_decap_3  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__085__A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_1_8 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 314 592
use scs8hd_nor2_4  _082_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_19 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_18
timestamp 1586364061
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_22
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_31
timestamp 1586364061
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_35
timestamp 1586364061
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_39 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 406 592
use scs8hd_buf_1  _164_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_44
timestamp 1586364061
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_45
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_56
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_66
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__C
timestamp 1586364061
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use scs8hd_inv_8  _067_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _069_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 866 592
use scs8hd_buf_1  _087_
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 8096 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_74
timestamp 1586364061
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_78
timestamp 1586364061
transform 1 0 8280 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_70
timestamp 1586364061
transform 1 0 7544 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_nor2_4  _177_
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 866 592
use scs8hd_nor2_4  _178_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 10580 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_103
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_97
timestamp 1586364061
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_123
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_129
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_130
timestamp 1586364061
transform 1 0 13064 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_125
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12788 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13248 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 314 592
use scs8hd_inv_8  _108_
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 866 592
use scs8hd_or4_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_139
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use scs8hd_inv_8  _073_
timestamp 1586364061
transform 1 0 15548 0 -1 2720
box -38 -48 866 592
use scs8hd_or3_4  _075_
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _093_
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__C
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__D
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 17572 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_177
timestamp 1586364061
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_181
timestamp 1586364061
transform 1 0 17756 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__B
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_buf_1  _076_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_187
timestamp 1586364061
transform 1 0 18308 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_185
timestamp 1586364061
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__137__C
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 18492 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_191
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_192
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_206
timestamp 1586364061
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_210
timestamp 1586364061
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__145__B
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 20792 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__C
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20792 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_225
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_229
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22356 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_240
timestamp 1586364061
transform 1 0 23184 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__C
timestamp 1586364061
transform 1 0 23000 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_247
timestamp 1586364061
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_244
timestamp 1586364061
transform 1 0 23552 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24104 0 -1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 25208 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_256
timestamp 1586364061
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_260
timestamp 1586364061
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_268
timestamp 1586364061
transform 1 0 25760 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_264
timestamp 1586364061
transform 1 0 25392 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_263
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _190_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_270
timestamp 1586364061
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26496 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26128 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26220 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_0_278
timestamp 1586364061
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_286
timestamp 1586364061
transform 1 0 27416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_282
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_283
timestamp 1586364061
transform 1 0 27140 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27232 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27324 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_287
timestamp 1586364061
transform 1 0 27508 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27600 0 1 2720
box -38 -48 222 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 27784 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_293
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_294
timestamp 1586364061
transform 1 0 28152 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 28244 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27876 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_298
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28336 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 28980 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_0_309
timestamp 1586364061
transform 1 0 29532 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_305
timestamp 1586364061
transform 1 0 29164 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29348 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_316
timestamp 1586364061
transform 1 0 30176 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30360 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29348 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _161_
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 866 592
use scs8hd_conb_1  _191_
timestamp 1586364061
transform 1 0 30912 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30728 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_320 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 30544 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_331
timestamp 1586364061
transform 1 0 31556 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_320
timestamp 1586364061
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_327
timestamp 1586364061
transform 1 0 31188 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_335
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_342
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_339
timestamp 1586364061
transform 1 0 32292 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_354
timestamp 1586364061
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_351
timestamp 1586364061
transform 1 0 33396 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_366
timestamp 1586364061
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_1_363
timestamp 1586364061
transform 1 0 34500 0 1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_15
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_19
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_35
timestamp 1586364061
transform 1 0 4324 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_46
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_4  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_1  _084_
timestamp 1586364061
transform 1 0 6348 0 -1 3808
box -38 -48 314 592
use scs8hd_or3_4  _086_
timestamp 1586364061
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__C
timestamp 1586364061
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_56
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_77
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_81
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 590 592
use scs8hd_nor2_4  _176_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 590 592
use scs8hd_inv_8  _068_
timestamp 1586364061
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_112
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use scs8hd_nand2_4  _109_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_126
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_130
timestamp 1586364061
transform 1 0 13064 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_151
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _094_
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__D
timestamp 1586364061
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__B
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_158
timestamp 1586364061
transform 1 0 15640 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__C
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_171
timestamp 1586364061
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_175
timestamp 1586364061
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use scs8hd_or4_4  _137_
timestamp 1586364061
transform 1 0 17756 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__C
timestamp 1586364061
transform 1 0 18768 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_190
timestamp 1586364061
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use scs8hd_or2_4  _145_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19320 0 -1 3808
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_194
timestamp 1586364061
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _156_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__156__B
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 22632 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_228
timestamp 1586364061
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_232
timestamp 1586364061
transform 1 0 22448 0 -1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _158_
timestamp 1586364061
transform 1 0 22816 0 -1 3808
box -38 -48 1234 592
use scs8hd_fill_2  FILLER_2_249
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_8  _159_
timestamp 1586364061
transform 1 0 24748 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24564 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_266
timestamp 1586364061
transform 1 0 25576 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_272
timestamp 1586364061
transform 1 0 26128 0 -1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26956 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_279
timestamp 1586364061
transform 1 0 26772 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_283
timestamp 1586364061
transform 1 0 27140 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_8  FILLER_2_300
timestamp 1586364061
transform 1 0 28704 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_12  FILLER_2_317
timestamp 1586364061
transform 1 0 30268 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_2_329
timestamp 1586364061
transform 1 0 31372 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_335
timestamp 1586364061
transform 1 0 31924 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_nor2_4  _169_
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_17
timestamp 1586364061
transform 1 0 2668 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_21
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_34
timestamp 1586364061
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _081_
timestamp 1586364061
transform 1 0 5704 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 5520 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_42
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_46
timestamp 1586364061
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _083_
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _179_
timestamp 1586364061
transform 1 0 9936 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__080__C
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_92
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _174_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _074_
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_142
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_146
timestamp 1586364061
transform 1 0 14536 0 1 3808
box -38 -48 130 592
use scs8hd_or4_4  _095_
timestamp 1586364061
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__163__B
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_158
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_162
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__C
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_175
timestamp 1586364061
transform 1 0 17204 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_or3_4  _119_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_193
timestamp 1586364061
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use scs8hd_or4_4  _147_
timestamp 1586364061
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_197
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__D
timestamp 1586364061
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_210
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_nor3_4  _155_
timestamp 1586364061
transform 1 0 21620 0 1 3808
box -38 -48 1234 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 23920 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__C
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_236
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_240
timestamp 1586364061
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_250
timestamp 1586364061
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26220 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 25668 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26036 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_265
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 222 592
use scs8hd_buf_1  _130_
timestamp 1586364061
transform 1 0 27784 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_282
timestamp 1586364061
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_286
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 28244 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_293
timestamp 1586364061
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 406 592
use scs8hd_buf_1  _120_
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_309
timestamp 1586364061
transform 1 0 29532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_313
timestamp 1586364061
transform 1 0 29900 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 30728 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_320
timestamp 1586364061
transform 1 0 30544 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_324
timestamp 1586364061
transform 1 0 30912 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_336
timestamp 1586364061
transform 1 0 32016 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_348
timestamp 1586364061
transform 1 0 33120 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_3_360
timestamp 1586364061
transform 1 0 34224 0 1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 130 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3680 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_30
timestamp 1586364061
transform 1 0 3864 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 590 592
use scs8hd_or3_4  _098_
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _090_
timestamp 1586364061
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_58
timestamp 1586364061
transform 1 0 6440 0 -1 4896
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_81
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _080_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_85
timestamp 1586364061
transform 1 0 8924 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_89
timestamp 1586364061
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_106
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_114
timestamp 1586364061
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_128
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_132
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_or2_4  _171_
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_161
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 130 592
use scs8hd_or4_4  _163_
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use scs8hd_fill_1  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _078_
timestamp 1586364061
transform 1 0 19780 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_195
timestamp 1586364061
transform 1 0 19044 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_199
timestamp 1586364061
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_conb_1  _189_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 406 592
use scs8hd_nor3_4  _157_
timestamp 1586364061
transform 1 0 22080 0 -1 4896
box -38 -48 1234 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 21620 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_225
timestamp 1586364061
transform 1 0 21804 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_241
timestamp 1586364061
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_6  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 590 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24472 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_253
timestamp 1586364061
transform 1 0 24380 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_256
timestamp 1586364061
transform 1 0 24656 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_8  _162_
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_266
timestamp 1586364061
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27508 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_285
timestamp 1586364061
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_289
timestamp 1586364061
transform 1 0 27692 0 -1 4896
box -38 -48 406 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_8  FILLER_4_302
timestamp 1586364061
transform 1 0 28888 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29624 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 30084 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_313
timestamp 1586364061
transform 1 0 29900 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_317
timestamp 1586364061
transform 1 0 30268 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_4_329
timestamp 1586364061
transform 1 0 31372 0 -1 4896
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_335
timestamp 1586364061
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_24
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 3680 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_39
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _070_
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_43
timestamp 1586364061
transform 1 0 5060 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_47
timestamp 1586364061
transform 1 0 5428 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_buf_1  _099_
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__165__B
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_68
timestamp 1586364061
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_72
timestamp 1586364061
transform 1 0 7728 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_99
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12052 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_5_121
timestamp 1586364061
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13064 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12880 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_127
timestamp 1586364061
transform 1 0 12788 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14628 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_139
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_143
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _173_
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__173__B
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_156
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_160
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__163__D
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use scs8hd_or2_4  _072_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_191
timestamp 1586364061
transform 1 0 18676 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _160_
timestamp 1586364061
transform 1 0 21252 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_217
timestamp 1586364061
transform 1 0 21068 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_234
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_238
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_242
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 25208 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_254
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_258
timestamp 1586364061
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_271
timestamp 1586364061
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_275
timestamp 1586364061
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_279
timestamp 1586364061
transform 1 0 26772 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28520 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28888 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_291
timestamp 1586364061
transform 1 0 27876 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_295
timestamp 1586364061
transform 1 0 28244 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_300
timestamp 1586364061
transform 1 0 28704 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_304
timestamp 1586364061
transform 1 0 29072 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_309
timestamp 1586364061
transform 1 0 29532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_313
timestamp 1586364061
transform 1 0 29900 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30728 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_320
timestamp 1586364061
transform 1 0 30544 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_324
timestamp 1586364061
transform 1 0 30912 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_331
timestamp 1586364061
transform 1 0 31556 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32108 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_335
timestamp 1586364061
transform 1 0 31924 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_339
timestamp 1586364061
transform 1 0 32292 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33396 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34040 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_353
timestamp 1586364061
transform 1 0 33580 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_357
timestamp 1586364061
transform 1 0 33948 0 1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35328 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34408 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_360
timestamp 1586364061
transform 1 0 34224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_370
timestamp 1586364061
transform 1 0 35144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_374
timestamp 1586364061
transform 1 0 35512 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_378
timestamp 1586364061
transform 1 0 35880 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_381
timestamp 1586364061
transform 1 0 36156 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_393
timestamp 1586364061
transform 1 0 37260 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_405
timestamp 1586364061
transform 1 0 38364 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _200_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_17
timestamp 1586364061
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_21
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_25
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_26
timestamp 1586364061
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_29
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_30
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_43
timestamp 1586364061
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_47
timestamp 1586364061
transform 1 0 5428 0 1 5984
box -38 -48 774 592
use scs8hd_nor2_4  _165_
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _167_
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__167__B
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_85
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_88
timestamp 1586364061
transform 1 0 9200 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_92
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_99
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_116
timestamp 1586364061
transform 1 0 11776 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_113
timestamp 1586364061
transform 1 0 11500 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_117
timestamp 1586364061
transform 1 0 11868 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_120
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13064 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_128
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_132
timestamp 1586364061
transform 1 0 13248 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _071_
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_145
timestamp 1586364061
transform 1 0 14444 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_149
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__D
timestamp 1586364061
transform 1 0 16376 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_168
timestamp 1586364061
transform 1 0 16560 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_7_178
timestamp 1586364061
transform 1 0 17480 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_181
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_184
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_180
timestamp 1586364061
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18584 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_201
timestamp 1586364061
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_216
timestamp 1586364061
transform 1 0 20976 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_220
timestamp 1586364061
transform 1 0 21344 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 21988 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_229
timestamp 1586364061
transform 1 0 22172 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_234
timestamp 1586364061
transform 1 0 22632 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_224
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23184 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_236
timestamp 1586364061
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_240
timestamp 1586364061
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use scs8hd_or2_4  _129_
timestamp 1586364061
transform 1 0 24932 0 -1 5984
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24380 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_255
timestamp 1586364061
transform 1 0 24564 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_256
timestamp 1586364061
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_260
timestamp 1586364061
transform 1 0 25024 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_265
timestamp 1586364061
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_266
timestamp 1586364061
transform 1 0 25576 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26956 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26772 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_290
timestamp 1586364061
transform 1 0 27784 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_280
timestamp 1586364061
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_284
timestamp 1586364061
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28520 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27968 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_294
timestamp 1586364061
transform 1 0 28152 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_297
timestamp 1586364061
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_301
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 30084 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29532 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_307
timestamp 1586364061
transform 1 0 29348 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_311
timestamp 1586364061
transform 1 0 29716 0 -1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_315
timestamp 1586364061
transform 1 0 30084 0 1 5984
box -38 -48 406 592
use scs8hd_nor2_4  _136_
timestamp 1586364061
transform 1 0 31096 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 30912 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 31096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_324
timestamp 1586364061
transform 1 0 30912 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_328
timestamp 1586364061
transform 1 0 31280 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_7_321
timestamp 1586364061
transform 1 0 30636 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_339
timestamp 1586364061
transform 1 0 32292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_335
timestamp 1586364061
transform 1 0 31924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_6  FILLER_6_345
timestamp 1586364061
transform 1 0 32844 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_6_340
timestamp 1586364061
transform 1 0 32384 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 32476 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 32660 0 1 5984
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33396 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33856 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_354
timestamp 1586364061
transform 1 0 33672 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_354
timestamp 1586364061
transform 1 0 33672 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_358
timestamp 1586364061
transform 1 0 34040 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34224 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_371
timestamp 1586364061
transform 1 0 35236 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_362
timestamp 1586364061
transform 1 0 34408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_376
timestamp 1586364061
transform 1 0 35696 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_375
timestamp 1586364061
transform 1 0 35604 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 35972 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_387
timestamp 1586364061
transform 1 0 36708 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_381
timestamp 1586364061
transform 1 0 36156 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_382
timestamp 1586364061
transform 1 0 36248 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36432 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36432 0 1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_386
timestamp 1586364061
transform 1 0 36616 0 -1 5984
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_394
timestamp 1586364061
transform 1 0 37352 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_3
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_8_9
timestamp 1586364061
transform 1 0 1932 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_44
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6532 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_8_56
timestamp 1586364061
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_6  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_88
timestamp 1586364061
transform 1 0 9200 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_12  FILLER_8_104
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11960 0 -1 7072
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_8_116
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_8_135
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15732 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use scs8hd_or2_4  _077_
timestamp 1586364061
transform 1 0 17572 0 -1 7072
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_174
timestamp 1586364061
transform 1 0 17112 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_186
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_190
timestamp 1586364061
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18952 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_8_205
timestamp 1586364061
transform 1 0 19964 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_224
timestamp 1586364061
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_228
timestamp 1586364061
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_235
timestamp 1586364061
transform 1 0 22724 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 23736 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  FILLER_8_243
timestamp 1586364061
transform 1 0 23460 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_255
timestamp 1586364061
transform 1 0 24564 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _122_
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_266
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_8_271
timestamp 1586364061
transform 1 0 26036 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27048 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26680 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_280
timestamp 1586364061
transform 1 0 26864 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_291
timestamp 1586364061
transform 1 0 27876 0 -1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__135__B
timestamp 1586364061
transform 1 0 30268 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_308
timestamp 1586364061
transform 1 0 29440 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_316
timestamp 1586364061
transform 1 0 30176 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _135_
timestamp 1586364061
transform 1 0 30452 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_328
timestamp 1586364061
transform 1 0 31280 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_348
timestamp 1586364061
transform 1 0 33120 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_8_354
timestamp 1586364061
transform 1 0 33672 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_358
timestamp 1586364061
transform 1 0 34040 0 -1 7072
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34408 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_371
timestamp 1586364061
transform 1 0 35236 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35972 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_4  FILLER_8_375
timestamp 1586364061
transform 1 0 35604 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_388
timestamp 1586364061
transform 1 0 36800 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_396
timestamp 1586364061
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 1050 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_23
timestamp 1586364061
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_27
timestamp 1586364061
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 5612 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_44
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_51
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 406 592
use scs8hd_buf_1  _091_
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_65
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_69
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_90
timestamp 1586364061
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_94
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_107
timestamp 1586364061
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12512 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_111
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_131
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_148
timestamp 1586364061
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15548 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_155
timestamp 1586364061
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_159
timestamp 1586364061
transform 1 0 15732 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_180
timestamp 1586364061
transform 1 0 17664 0 1 7072
box -38 -48 314 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20148 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_199
timestamp 1586364061
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_210
timestamp 1586364061
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_214
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_218
timestamp 1586364061
transform 1 0 21160 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_236
timestamp 1586364061
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_240
timestamp 1586364061
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_254
timestamp 1586364061
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_262
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_266
timestamp 1586364061
transform 1 0 25576 0 1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 27048 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_280
timestamp 1586364061
transform 1 0 26864 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_284
timestamp 1586364061
transform 1 0 27232 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28888 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_297
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_301
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_9_304
timestamp 1586364061
transform 1 0 29072 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 30084 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 29900 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29440 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_306
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_310
timestamp 1586364061
transform 1 0 29624 0 1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_9_326
timestamp 1586364061
transform 1 0 31096 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32200 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 32660 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_341
timestamp 1586364061
transform 1 0 32476 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_345
timestamp 1586364061
transform 1 0 32844 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 33028 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_358
timestamp 1586364061
transform 1 0 34040 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 34224 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_362
timestamp 1586364061
transform 1 0 34408 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _209_
timestamp 1586364061
transform 1 0 36432 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 35880 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_376
timestamp 1586364061
transform 1 0 35696 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_380
timestamp 1586364061
transform 1 0 36064 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__209__A
timestamp 1586364061
transform 1 0 36984 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_388
timestamp 1586364061
transform 1 0 36800 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_392
timestamp 1586364061
transform 1 0 37168 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_9_404
timestamp 1586364061
transform 1 0 38272 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2944 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_18
timestamp 1586364061
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_22
timestamp 1586364061
transform 1 0 3128 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_2  _195_
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_53
timestamp 1586364061
transform 1 0 5980 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_57
timestamp 1586364061
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_73
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 314 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_8  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13064 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_128
timestamp 1586364061
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_149
timestamp 1586364061
transform 1 0 14812 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_165
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_169
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_187
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_191
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_204
timestamp 1586364061
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_4  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_8  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 774 592
use scs8hd_or2_4  _121_
timestamp 1586364061
transform 1 0 23000 0 -1 8160
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_249
timestamp 1586364061
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_253
timestamp 1586364061
transform 1 0 24380 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_265
timestamp 1586364061
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27692 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_287
timestamp 1586364061
transform 1 0 27508 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28888 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_10_291
timestamp 1586364061
transform 1 0 27876 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_299
timestamp 1586364061
transform 1 0 28612 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30084 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_313
timestamp 1586364061
transform 1 0 29900 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_317
timestamp 1586364061
transform 1 0 30268 0 -1 8160
box -38 -48 222 592
use scs8hd_conb_1  _187_
timestamp 1586364061
transform 1 0 30636 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 30452 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_324
timestamp 1586364061
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 32476 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 32292 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_344
timestamp 1586364061
transform 1 0 32752 0 -1 8160
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 33488 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_348
timestamp 1586364061
transform 1 0 33120 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_351
timestamp 1586364061
transform 1 0 33396 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 35236 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_363
timestamp 1586364061
transform 1 0 34500 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_10_369
timestamp 1586364061
transform 1 0 35052 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_380
timestamp 1586364061
transform 1 0 36064 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_10_392
timestamp 1586364061
transform 1 0 37168 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_396
timestamp 1586364061
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3588 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_21
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_25
timestamp 1586364061
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use scs8hd_buf_2  _199_
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_33
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_37
timestamp 1586364061
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_41
timestamp 1586364061
transform 1 0 4876 0 1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 6900 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_78
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_82
timestamp 1586364061
transform 1 0 8648 0 1 8160
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_112
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_116
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 590 592
use scs8hd_fill_2  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_138
timestamp 1586364061
transform 1 0 13800 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_142
timestamp 1586364061
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_178
timestamp 1586364061
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_194
timestamp 1586364061
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_198
timestamp 1586364061
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 21436 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 21252 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_217
timestamp 1586364061
transform 1 0 21068 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_230
timestamp 1586364061
transform 1 0 22264 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_234
timestamp 1586364061
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_238
timestamp 1586364061
transform 1 0 23000 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_256
timestamp 1586364061
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_260
timestamp 1586364061
transform 1 0 25024 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25668 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_264
timestamp 1586364061
transform 1 0 25392 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_276
timestamp 1586364061
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _134_
timestamp 1586364061
transform 1 0 27600 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 27416 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 26680 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 27048 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_280
timestamp 1586364061
transform 1 0 26864 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_284
timestamp 1586364061
transform 1 0 27232 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_297
timestamp 1586364061
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_301
timestamp 1586364061
transform 1 0 28796 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29992 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31556 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 31004 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31372 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_323
timestamp 1586364061
transform 1 0 30820 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_327
timestamp 1586364061
transform 1 0 31188 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32752 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 32108 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_334
timestamp 1586364061
transform 1 0 31832 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_339
timestamp 1586364061
transform 1 0 32292 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 33948 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_355
timestamp 1586364061
transform 1 0 33764 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_359
timestamp 1586364061
transform 1 0 34132 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_363
timestamp 1586364061
transform 1 0 34500 0 1 8160
box -38 -48 130 592
use scs8hd_buf_2  _208_
timestamp 1586364061
transform 1 0 36432 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 35880 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 36248 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_376
timestamp 1586364061
transform 1 0 35696 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_380
timestamp 1586364061
transform 1 0 36064 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__208__A
timestamp 1586364061
transform 1 0 36984 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_388
timestamp 1586364061
transform 1 0 36800 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_392
timestamp 1586364061
transform 1 0 37168 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_11_404
timestamp 1586364061
transform 1 0 38272 0 1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_6
timestamp 1586364061
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_10
timestamp 1586364061
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_50
timestamp 1586364061
transform 1 0 5704 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7452 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_67
timestamp 1586364061
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _166_
timestamp 1586364061
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_12_71
timestamp 1586364061
transform 1 0 7636 0 -1 9248
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_96
timestamp 1586364061
transform 1 0 9936 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11040 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10856 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_100
timestamp 1586364061
transform 1 0 10304 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_104
timestamp 1586364061
transform 1 0 10672 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_119
timestamp 1586364061
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_125
timestamp 1586364061
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_133
timestamp 1586364061
transform 1 0 13340 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_158
timestamp 1586364061
transform 1 0 15640 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_181
timestamp 1586364061
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_185
timestamp 1586364061
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_189
timestamp 1586364061
transform 1 0 18492 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_206
timestamp 1586364061
transform 1 0 20056 0 -1 9248
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 21436 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_218
timestamp 1586364061
transform 1 0 21160 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 22264 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 21804 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_223
timestamp 1586364061
transform 1 0 21620 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 23828 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_258
timestamp 1586364061
transform 1 0 24840 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_262
timestamp 1586364061
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25392 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_266
timestamp 1586364061
transform 1 0 25576 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_272
timestamp 1586364061
transform 1 0 26128 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_285
timestamp 1586364061
transform 1 0 27324 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_12_290
timestamp 1586364061
transform 1 0 27784 0 -1 9248
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28612 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_296
timestamp 1586364061
transform 1 0 28336 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 29992 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_310
timestamp 1586364061
transform 1 0 29624 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  FILLER_12_316
timestamp 1586364061
transform 1 0 30176 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 30452 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_12_328
timestamp 1586364061
transform 1 0 31280 0 -1 9248
box -38 -48 774 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 33672 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33120 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 33488 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_346
timestamp 1586364061
transform 1 0 32936 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_350
timestamp 1586364061
transform 1 0 33304 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 34868 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_365
timestamp 1586364061
transform 1 0 34684 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_369
timestamp 1586364061
transform 1 0 35052 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 36616 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_384
timestamp 1586364061
transform 1 0 36432 0 -1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_388
timestamp 1586364061
transform 1 0 36800 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_396
timestamp 1586364061
transform 1 0 37536 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2208 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _168_
timestamp 1586364061
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_21
timestamp 1586364061
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_25
timestamp 1586364061
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_18
timestamp 1586364061
transform 1 0 2760 0 -1 10336
box -38 -48 1142 592
use scs8hd_nor2_4  _170_
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_29
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_42
timestamp 1586364061
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_43
timestamp 1586364061
transform 1 0 5060 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_55
timestamp 1586364061
transform 1 0 6164 0 -1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _180_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use scs8hd_conb_1  _183_
timestamp 1586364061
transform 1 0 6532 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__180__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_62
timestamp 1586364061
transform 1 0 6808 0 -1 10336
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_71
timestamp 1586364061
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_75
timestamp 1586364061
transform 1 0 8004 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_73
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_90
timestamp 1586364061
transform 1 0 9384 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9568 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_94
timestamp 1586364061
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_109
timestamp 1586364061
transform 1 0 11132 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_97
timestamp 1586364061
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_110
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_143
timestamp 1586364061
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_162
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_166
timestamp 1586364061
transform 1 0 16376 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_158
timestamp 1586364061
transform 1 0 15640 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _175_
timestamp 1586364061
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_177
timestamp 1586364061
transform 1 0 17388 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_188
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_189
timestamp 1586364061
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_192
timestamp 1586364061
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _115_
timestamp 1586364061
transform 1 0 19136 0 -1 10336
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20976 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_209
timestamp 1586364061
transform 1 0 20332 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_227
timestamp 1586364061
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_231
timestamp 1586364061
transform 1 0 22356 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_224
timestamp 1586364061
transform 1 0 21712 0 -1 10336
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23000 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_236
timestamp 1586364061
transform 1 0 22816 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_240
timestamp 1586364061
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_236
timestamp 1586364061
transform 1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_248
timestamp 1586364061
transform 1 0 23920 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24656 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24472 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 24104 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24840 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 25208 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_256
timestamp 1586364061
transform 1 0 24656 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_260
timestamp 1586364061
transform 1 0 25024 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_252
timestamp 1586364061
transform 1 0 24288 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 25392 0 1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 26496 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_273
timestamp 1586364061
transform 1 0 26220 0 1 9248
box -38 -48 314 592
use scs8hd_decap_6  FILLER_14_265
timestamp 1586364061
transform 1 0 25484 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_273
timestamp 1586364061
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 27600 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 27416 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 27784 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 27048 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_278
timestamp 1586364061
transform 1 0 26680 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_284
timestamp 1586364061
transform 1 0 27232 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_285
timestamp 1586364061
transform 1 0 27324 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_289
timestamp 1586364061
transform 1 0 27692 0 -1 10336
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 28520 0 -1 10336
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_297
timestamp 1586364061
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_301
timestamp 1586364061
transform 1 0 28796 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_292
timestamp 1586364061
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 29716 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_317
timestamp 1586364061
transform 1 0 30268 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_309
timestamp 1586364061
transform 1 0 29532 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_313
timestamp 1586364061
transform 1 0 29900 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_317
timestamp 1586364061
transform 1 0 30268 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31280 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30452 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 31464 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_321
timestamp 1586364061
transform 1 0 30636 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_325
timestamp 1586364061
transform 1 0 31004 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_331
timestamp 1586364061
transform 1 0 31556 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_327
timestamp 1586364061
transform 1 0 31188 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_14_332
timestamp 1586364061
transform 1 0 31648 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_335
timestamp 1586364061
transform 1 0 31924 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 32292 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 32108 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31740 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_14_345
timestamp 1586364061
transform 1 0 32844 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_341
timestamp 1586364061
transform 1 0 32476 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 32660 0 -1 10336
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 32292 0 1 9248
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 32936 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 33488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33856 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 33948 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_350
timestamp 1586364061
transform 1 0 33304 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_358
timestamp 1586364061
transform 1 0 34040 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_355
timestamp 1586364061
transform 1 0 33764 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_359
timestamp 1586364061
transform 1 0 34132 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34500 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34224 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_362
timestamp 1586364061
transform 1 0 34408 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_372
timestamp 1586364061
transform 1 0 35328 0 -1 10336
box -38 -48 774 592
use scs8hd_buf_2  _202_
timestamp 1586364061
transform 1 0 36064 0 -1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 36432 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 36064 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 36616 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_376
timestamp 1586364061
transform 1 0 35696 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_382
timestamp 1586364061
transform 1 0 36248 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_384
timestamp 1586364061
transform 1 0 36432 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_393
timestamp 1586364061
transform 1 0 37260 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_388
timestamp 1586364061
transform 1 0 36800 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_396
timestamp 1586364061
transform 1 0 37536 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_405
timestamp 1586364061
transform 1 0 38364 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _198_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_7
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_11
timestamp 1586364061
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 3312 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_18
timestamp 1586364061
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_22
timestamp 1586364061
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_33
timestamp 1586364061
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_37
timestamp 1586364061
transform 1 0 4508 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_41
timestamp 1586364061
transform 1 0 4876 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use scs8hd_conb_1  _181_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_15_65
timestamp 1586364061
transform 1 0 7084 0 1 10336
box -38 -48 774 592
use scs8hd_buf_1  _104_
timestamp 1586364061
transform 1 0 8096 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 8556 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_73
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_79
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_83
timestamp 1586364061
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_94
timestamp 1586364061
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_107
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_111
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_114
timestamp 1586364061
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_136
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use scs8hd_conb_1  _182_
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_143
timestamp 1586364061
transform 1 0 14260 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_160
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_164
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 590 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 18400 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19964 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_201
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _138_
timestamp 1586364061
transform 1 0 21528 0 1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_225
timestamp 1586364061
transform 1 0 21804 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23920 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_236
timestamp 1586364061
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_240
timestamp 1586364061
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24472 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 24288 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_250
timestamp 1586364061
transform 1 0 24104 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 26036 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_263
timestamp 1586364061
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_267
timestamp 1586364061
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _140_
timestamp 1586364061
transform 1 0 27600 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 27416 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27048 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_280
timestamp 1586364061
transform 1 0 26864 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_284
timestamp 1586364061
transform 1 0 27232 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 28612 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_297
timestamp 1586364061
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_301
timestamp 1586364061
transform 1 0 28796 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29900 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29716 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_310
timestamp 1586364061
transform 1 0 29624 0 1 10336
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 31280 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30912 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_322
timestamp 1586364061
transform 1 0 30728 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_326
timestamp 1586364061
transform 1 0 31096 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 32844 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__144__B
timestamp 1586364061
transform 1 0 32476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_339
timestamp 1586364061
transform 1 0 32292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_343
timestamp 1586364061
transform 1 0 32660 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _144_
timestamp 1586364061
transform 1 0 33028 0 1 10336
box -38 -48 866 592
use scs8hd_decap_4  FILLER_15_356
timestamp 1586364061
transform 1 0 33856 0 1 10336
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__207__A
timestamp 1586364061
transform 1 0 34316 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_360
timestamp 1586364061
transform 1 0 34224 0 1 10336
box -38 -48 130 592
use scs8hd_decap_3  FILLER_15_363
timestamp 1586364061
transform 1 0 34500 0 1 10336
box -38 -48 314 592
use scs8hd_buf_2  _201_
timestamp 1586364061
transform 1 0 36432 0 1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 35880 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 36248 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_376
timestamp 1586364061
transform 1 0 35696 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_380
timestamp 1586364061
transform 1 0 36064 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 37536 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 36984 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 37996 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_388
timestamp 1586364061
transform 1 0 36800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_392
timestamp 1586364061
transform 1 0 37168 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_399
timestamp 1586364061
transform 1 0 37812 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_buf_2  _197_
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_7
timestamp 1586364061
transform 1 0 1748 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_2  _192_
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_19
timestamp 1586364061
transform 1 0 2852 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_35
timestamp 1586364061
transform 1 0 4324 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_59
timestamp 1586364061
transform 1 0 6532 0 -1 11424
box -38 -48 1142 592
use scs8hd_buf_1  _106_
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_71
timestamp 1586364061
transform 1 0 7636 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_79
timestamp 1586364061
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _107_
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_104
timestamp 1586364061
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_108
timestamp 1586364061
transform 1 0 11040 0 -1 11424
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_121
timestamp 1586364061
transform 1 0 12236 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _113_
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_132
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_144
timestamp 1586364061
transform 1 0 14352 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 15456 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_165
timestamp 1586364061
transform 1 0 16284 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_16_177
timestamp 1586364061
transform 1 0 17388 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18124 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_16_188
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 19136 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20148 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_205
timestamp 1586364061
transform 1 0 19964 0 -1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_209
timestamp 1586364061
transform 1 0 20332 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_224
timestamp 1586364061
transform 1 0 21712 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_16_236
timestamp 1586364061
transform 1 0 22816 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_240
timestamp 1586364061
transform 1 0 23184 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_244
timestamp 1586364061
transform 1 0 23552 0 -1 11424
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 24288 0 -1 11424
box -38 -48 866 592
use scs8hd_decap_12  FILLER_16_261
timestamp 1586364061
transform 1 0 25116 0 -1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_273
timestamp 1586364061
transform 1 0 26220 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 27784 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_279
timestamp 1586364061
transform 1 0 26772 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_287
timestamp 1586364061
transform 1 0 27508 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_299
timestamp 1586364061
transform 1 0 28612 0 -1 11424
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29716 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 31464 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_320
timestamp 1586364061
transform 1 0 30544 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_328
timestamp 1586364061
transform 1 0 31280 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_332
timestamp 1586364061
transform 1 0 31648 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_346
timestamp 1586364061
transform 1 0 32936 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_358
timestamp 1586364061
transform 1 0 34040 0 -1 11424
box -38 -48 314 592
use scs8hd_buf_2  _205_
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 406 592
use scs8hd_buf_2  _207_
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 34868 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 35236 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_365
timestamp 1586364061
transform 1 0 34684 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_369
timestamp 1586364061
transform 1 0 35052 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_2  _206_
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_377
timestamp 1586364061
transform 1 0 35788 0 -1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_389
timestamp 1586364061
transform 1 0 36892 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _196_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_22
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_26
timestamp 1586364061
transform 1 0 3496 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_38
timestamp 1586364061
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_94
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use scs8hd_nor2_4  _105_
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_106
timestamp 1586364061
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _184_
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_155
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_161
timestamp 1586364061
transform 1 0 15916 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_173
timestamp 1586364061
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 18584 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_181
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _185_
timestamp 1586364061
transform 1 0 19688 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_201
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_205
timestamp 1586364061
transform 1 0 19964 0 1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20700 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_216
timestamp 1586364061
transform 1 0 20976 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_251
timestamp 1586364061
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_256
timestamp 1586364061
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_260
timestamp 1586364061
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _186_
timestamp 1586364061
transform 1 0 25392 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_267
timestamp 1586364061
transform 1 0 25668 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_279
timestamp 1586364061
transform 1 0 26772 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_291
timestamp 1586364061
transform 1 0 27876 0 1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_17_303
timestamp 1586364061
transform 1 0 28980 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29992 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_317
timestamp 1586364061
transform 1 0 30268 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 31188 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31648 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30452 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_321
timestamp 1586364061
transform 1 0 30636 0 1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_334
timestamp 1586364061
transform 1 0 31832 0 1 11424
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 33764 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_346
timestamp 1586364061
transform 1 0 32936 0 1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_358
timestamp 1586364061
transform 1 0 34040 0 1 11424
box -38 -48 222 592
use scs8hd_buf_2  _204_
timestamp 1586364061
transform 1 0 35420 0 1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 35236 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34224 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 34592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_362
timestamp 1586364061
transform 1 0 34408 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 36524 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_377
timestamp 1586364061
transform 1 0 35788 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_381
timestamp 1586364061
transform 1 0 36156 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 36984 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_388
timestamp 1586364061
transform 1 0 36800 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_392
timestamp 1586364061
transform 1 0 37168 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_17_404
timestamp 1586364061
transform 1 0 38272 0 1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_9
timestamp 1586364061
transform 1 0 1932 0 -1 12512
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_20
timestamp 1586364061
transform 1 0 2944 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_28
timestamp 1586364061
transform 1 0 3680 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_99
timestamp 1586364061
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_18_110
timestamp 1586364061
transform 1 0 11224 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_122
timestamp 1586364061
transform 1 0 12328 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_134
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_146
timestamp 1586364061
transform 1 0 14536 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_152
timestamp 1586364061
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 590 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 19136 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_199
timestamp 1586364061
transform 1 0 19412 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_211
timestamp 1586364061
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24012 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_247
timestamp 1586364061
transform 1 0 23828 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 25024 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_252
timestamp 1586364061
transform 1 0 24288 0 -1 12512
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 774 592
use scs8hd_conb_1  _188_
timestamp 1586364061
transform 1 0 29532 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_308
timestamp 1586364061
transform 1 0 29440 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_buf_2  _203_
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_364
timestamp 1586364061
transform 1 0 34592 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_372
timestamp 1586364061
transform 1 0 35328 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_377
timestamp 1586364061
transform 1 0 35788 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_389
timestamp 1586364061
transform 1 0 36892 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_buf_2  _193_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_buf_2  _194_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 590 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24196 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_254
timestamp 1586364061
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_258
timestamp 1586364061
transform 1 0 24840 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_270
timestamp 1586364061
transform 1 0 25944 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_282
timestamp 1586364061
transform 1 0 27048 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_294
timestamp 1586364061
transform 1 0 28152 0 1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_302
timestamp 1586364061
transform 1 0 28888 0 1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 4986 0 5042 480 6 address[0]
port 0 nsew default input
rlabel metal2 s 8298 0 8354 480 6 address[1]
port 1 nsew default input
rlabel metal2 s 11610 0 11666 480 6 address[2]
port 2 nsew default input
rlabel metal2 s 15014 0 15070 480 6 address[3]
port 3 nsew default input
rlabel metal2 s 18326 0 18382 480 6 address[4]
port 4 nsew default input
rlabel metal2 s 21638 0 21694 480 6 address[5]
port 5 nsew default input
rlabel metal2 s 24950 0 25006 480 6 address[6]
port 6 nsew default input
rlabel metal2 s 31666 0 31722 480 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal2 s 34978 0 35034 480 6 bottom_grid_pin_4_
port 8 nsew default tristate
rlabel metal2 s 38290 0 38346 480 6 bottom_grid_pin_8_
port 9 nsew default tristate
rlabel metal3 s 0 416 480 536 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 1232 480 1352 6 chanx_left_in[1]
port 11 nsew default input
rlabel metal3 s 0 2184 480 2304 6 chanx_left_in[2]
port 12 nsew default input
rlabel metal3 s 0 3000 480 3120 6 chanx_left_in[3]
port 13 nsew default input
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[4]
port 14 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[5]
port 15 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[6]
port 16 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 17 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 18 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[0]
port 19 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[1]
port 20 nsew default tristate
rlabel metal3 s 0 10208 480 10328 6 chanx_left_out[2]
port 21 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[3]
port 22 nsew default tristate
rlabel metal3 s 0 11976 480 12096 6 chanx_left_out[4]
port 23 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 chanx_left_out[5]
port 24 nsew default tristate
rlabel metal3 s 0 13744 480 13864 6 chanx_left_out[6]
port 25 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[7]
port 26 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[8]
port 27 nsew default tristate
rlabel metal3 s 39520 416 40000 536 6 chanx_right_in[0]
port 28 nsew default input
rlabel metal3 s 39520 1232 40000 1352 6 chanx_right_in[1]
port 29 nsew default input
rlabel metal3 s 39520 2184 40000 2304 6 chanx_right_in[2]
port 30 nsew default input
rlabel metal3 s 39520 3000 40000 3120 6 chanx_right_in[3]
port 31 nsew default input
rlabel metal3 s 39520 3952 40000 4072 6 chanx_right_in[4]
port 32 nsew default input
rlabel metal3 s 39520 4768 40000 4888 6 chanx_right_in[5]
port 33 nsew default input
rlabel metal3 s 39520 5720 40000 5840 6 chanx_right_in[6]
port 34 nsew default input
rlabel metal3 s 39520 6536 40000 6656 6 chanx_right_in[7]
port 35 nsew default input
rlabel metal3 s 39520 7488 40000 7608 6 chanx_right_in[8]
port 36 nsew default input
rlabel metal3 s 39520 8440 40000 8560 6 chanx_right_out[0]
port 37 nsew default tristate
rlabel metal3 s 39520 9256 40000 9376 6 chanx_right_out[1]
port 38 nsew default tristate
rlabel metal3 s 39520 10208 40000 10328 6 chanx_right_out[2]
port 39 nsew default tristate
rlabel metal3 s 39520 11024 40000 11144 6 chanx_right_out[3]
port 40 nsew default tristate
rlabel metal3 s 39520 11976 40000 12096 6 chanx_right_out[4]
port 41 nsew default tristate
rlabel metal3 s 39520 12792 40000 12912 6 chanx_right_out[5]
port 42 nsew default tristate
rlabel metal3 s 39520 13744 40000 13864 6 chanx_right_out[6]
port 43 nsew default tristate
rlabel metal3 s 39520 14560 40000 14680 6 chanx_right_out[7]
port 44 nsew default tristate
rlabel metal3 s 39520 15512 40000 15632 6 chanx_right_out[8]
port 45 nsew default tristate
rlabel metal2 s 28354 0 28410 480 6 data_in
port 46 nsew default input
rlabel metal2 s 1674 0 1730 480 6 enable
port 47 nsew default input
rlabel metal2 s 2502 15520 2558 16000 6 top_grid_pin_0_
port 48 nsew default tristate
rlabel metal2 s 27434 15520 27490 16000 6 top_grid_pin_10_
port 49 nsew default tristate
rlabel metal2 s 32494 15520 32550 16000 6 top_grid_pin_12_
port 50 nsew default tristate
rlabel metal2 s 37462 15520 37518 16000 6 top_grid_pin_14_
port 51 nsew default tristate
rlabel metal2 s 7470 15520 7526 16000 6 top_grid_pin_2_
port 52 nsew default tristate
rlabel metal2 s 12438 15520 12494 16000 6 top_grid_pin_4_
port 53 nsew default tristate
rlabel metal2 s 17498 15520 17554 16000 6 top_grid_pin_6_
port 54 nsew default tristate
rlabel metal2 s 22466 15520 22522 16000 6 top_grid_pin_8_
port 55 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 56 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 57 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
