VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__2_
  CLASS BLOCK ;
  FOREIGN sb_0__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 111.600 28.890 114.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 2.400 ;
    END
  END SC_OUT_BOT
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.650 111.600 85.930 114.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 2.400 57.760 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 18.400 114.000 19.000 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 41.520 114.000 42.120 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 43.560 114.000 44.160 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 46.280 114.000 46.880 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 48.320 114.000 48.920 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 50.360 114.000 50.960 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 53.080 114.000 53.680 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 55.120 114.000 55.720 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 57.840 114.000 58.440 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 59.880 114.000 60.480 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 61.920 114.000 62.520 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 21.120 114.000 21.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 23.160 114.000 23.760 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 25.200 114.000 25.800 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 27.920 114.000 28.520 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 29.960 114.000 30.560 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 32.680 114.000 33.280 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 34.720 114.000 35.320 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 36.760 114.000 37.360 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 39.480 114.000 40.080 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 64.640 114.000 65.240 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 87.080 114.000 87.680 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 89.800 114.000 90.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 91.840 114.000 92.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 93.880 114.000 94.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 96.600 114.000 97.200 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 98.640 114.000 99.240 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 100.680 114.000 101.280 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 103.400 114.000 104.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 105.440 114.000 106.040 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 107.480 114.000 108.080 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 66.680 114.000 67.280 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 68.720 114.000 69.320 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 71.440 114.000 72.040 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 73.480 114.000 74.080 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 75.520 114.000 76.120 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 78.240 114.000 78.840 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 80.280 114.000 80.880 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 82.320 114.000 82.920 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 111.600 85.040 114.000 85.640 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.400 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.400 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.400 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.400 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.400 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.400 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 2.400 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 2.400 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.400 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 2.400 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.400 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 2.400 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 2.400 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 2.400 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 2.400 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 2.400 ;
    END
  END chany_bottom_out[9]
  PIN prog_clk_0_E_in
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 110.200 114.000 110.800 ;
    END
  END prog_clk_0_E_in
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 2.760 114.000 3.360 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 4.800 114.000 5.400 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 7.520 114.000 8.120 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 9.560 114.000 10.160 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 11.600 114.000 12.200 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 14.320 114.000 14.920 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 16.360 114.000 16.960 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 112.240 114.000 112.840 ;
    END
  END right_top_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 3.290 2.760 112.630 100.880 ;
      LAYER met2 ;
        RECT 1.010 111.320 28.330 112.725 ;
        RECT 29.170 111.320 85.370 112.725 ;
        RECT 86.210 111.320 112.600 112.725 ;
        RECT 1.010 2.680 112.600 111.320 ;
        RECT 1.570 0.835 3.030 2.680 ;
        RECT 3.870 0.835 5.790 2.680 ;
        RECT 6.630 0.835 8.550 2.680 ;
        RECT 9.390 0.835 11.310 2.680 ;
        RECT 12.150 0.835 14.070 2.680 ;
        RECT 14.910 0.835 16.830 2.680 ;
        RECT 17.670 0.835 19.590 2.680 ;
        RECT 20.430 0.835 22.350 2.680 ;
        RECT 23.190 0.835 25.110 2.680 ;
        RECT 25.950 0.835 27.870 2.680 ;
        RECT 28.710 0.835 30.170 2.680 ;
        RECT 31.010 0.835 32.930 2.680 ;
        RECT 33.770 0.835 35.690 2.680 ;
        RECT 36.530 0.835 38.450 2.680 ;
        RECT 39.290 0.835 41.210 2.680 ;
        RECT 42.050 0.835 43.970 2.680 ;
        RECT 44.810 0.835 46.730 2.680 ;
        RECT 47.570 0.835 49.490 2.680 ;
        RECT 50.330 0.835 52.250 2.680 ;
        RECT 53.090 0.835 55.010 2.680 ;
        RECT 55.850 0.835 57.770 2.680 ;
        RECT 58.610 0.835 60.070 2.680 ;
        RECT 60.910 0.835 62.830 2.680 ;
        RECT 63.670 0.835 65.590 2.680 ;
        RECT 66.430 0.835 68.350 2.680 ;
        RECT 69.190 0.835 71.110 2.680 ;
        RECT 71.950 0.835 73.870 2.680 ;
        RECT 74.710 0.835 76.630 2.680 ;
        RECT 77.470 0.835 79.390 2.680 ;
        RECT 80.230 0.835 82.150 2.680 ;
        RECT 82.990 0.835 84.910 2.680 ;
        RECT 85.750 0.835 87.210 2.680 ;
        RECT 88.050 0.835 89.970 2.680 ;
        RECT 90.810 0.835 92.730 2.680 ;
        RECT 93.570 0.835 95.490 2.680 ;
        RECT 96.330 0.835 98.250 2.680 ;
        RECT 99.090 0.835 101.010 2.680 ;
        RECT 101.850 0.835 103.770 2.680 ;
        RECT 104.610 0.835 106.530 2.680 ;
        RECT 107.370 0.835 109.290 2.680 ;
        RECT 110.130 0.835 112.050 2.680 ;
      LAYER met3 ;
        RECT 0.985 111.840 111.200 112.705 ;
        RECT 0.985 111.200 111.600 111.840 ;
        RECT 0.985 109.800 111.200 111.200 ;
        RECT 0.985 108.480 111.600 109.800 ;
        RECT 0.985 107.080 111.200 108.480 ;
        RECT 0.985 106.440 111.600 107.080 ;
        RECT 0.985 105.040 111.200 106.440 ;
        RECT 0.985 104.400 111.600 105.040 ;
        RECT 0.985 103.000 111.200 104.400 ;
        RECT 0.985 101.680 111.600 103.000 ;
        RECT 0.985 100.280 111.200 101.680 ;
        RECT 0.985 99.640 111.600 100.280 ;
        RECT 0.985 98.240 111.200 99.640 ;
        RECT 0.985 97.600 111.600 98.240 ;
        RECT 0.985 96.200 111.200 97.600 ;
        RECT 0.985 94.880 111.600 96.200 ;
        RECT 0.985 93.480 111.200 94.880 ;
        RECT 0.985 92.840 111.600 93.480 ;
        RECT 0.985 91.440 111.200 92.840 ;
        RECT 0.985 90.800 111.600 91.440 ;
        RECT 0.985 89.400 111.200 90.800 ;
        RECT 0.985 88.080 111.600 89.400 ;
        RECT 0.985 86.680 111.200 88.080 ;
        RECT 0.985 86.040 111.600 86.680 ;
        RECT 0.985 84.640 111.200 86.040 ;
        RECT 0.985 83.320 111.600 84.640 ;
        RECT 0.985 81.920 111.200 83.320 ;
        RECT 0.985 81.280 111.600 81.920 ;
        RECT 0.985 79.880 111.200 81.280 ;
        RECT 0.985 79.240 111.600 79.880 ;
        RECT 0.985 77.840 111.200 79.240 ;
        RECT 0.985 76.520 111.600 77.840 ;
        RECT 0.985 75.120 111.200 76.520 ;
        RECT 0.985 74.480 111.600 75.120 ;
        RECT 0.985 73.080 111.200 74.480 ;
        RECT 0.985 72.440 111.600 73.080 ;
        RECT 0.985 71.040 111.200 72.440 ;
        RECT 0.985 69.720 111.600 71.040 ;
        RECT 0.985 68.320 111.200 69.720 ;
        RECT 0.985 67.680 111.600 68.320 ;
        RECT 0.985 66.280 111.200 67.680 ;
        RECT 0.985 65.640 111.600 66.280 ;
        RECT 0.985 64.240 111.200 65.640 ;
        RECT 0.985 62.920 111.600 64.240 ;
        RECT 0.985 61.520 111.200 62.920 ;
        RECT 0.985 60.880 111.600 61.520 ;
        RECT 0.985 59.480 111.200 60.880 ;
        RECT 0.985 58.840 111.600 59.480 ;
        RECT 0.985 58.160 111.200 58.840 ;
        RECT 2.800 57.440 111.200 58.160 ;
        RECT 2.800 56.760 111.600 57.440 ;
        RECT 0.985 56.120 111.600 56.760 ;
        RECT 0.985 54.720 111.200 56.120 ;
        RECT 0.985 54.080 111.600 54.720 ;
        RECT 0.985 52.680 111.200 54.080 ;
        RECT 0.985 51.360 111.600 52.680 ;
        RECT 0.985 49.960 111.200 51.360 ;
        RECT 0.985 49.320 111.600 49.960 ;
        RECT 0.985 47.920 111.200 49.320 ;
        RECT 0.985 47.280 111.600 47.920 ;
        RECT 0.985 45.880 111.200 47.280 ;
        RECT 0.985 44.560 111.600 45.880 ;
        RECT 0.985 43.160 111.200 44.560 ;
        RECT 0.985 42.520 111.600 43.160 ;
        RECT 0.985 41.120 111.200 42.520 ;
        RECT 0.985 40.480 111.600 41.120 ;
        RECT 0.985 39.080 111.200 40.480 ;
        RECT 0.985 37.760 111.600 39.080 ;
        RECT 0.985 36.360 111.200 37.760 ;
        RECT 0.985 35.720 111.600 36.360 ;
        RECT 0.985 34.320 111.200 35.720 ;
        RECT 0.985 33.680 111.600 34.320 ;
        RECT 0.985 32.280 111.200 33.680 ;
        RECT 0.985 30.960 111.600 32.280 ;
        RECT 0.985 29.560 111.200 30.960 ;
        RECT 0.985 28.920 111.600 29.560 ;
        RECT 0.985 27.520 111.200 28.920 ;
        RECT 0.985 26.200 111.600 27.520 ;
        RECT 0.985 24.800 111.200 26.200 ;
        RECT 0.985 24.160 111.600 24.800 ;
        RECT 0.985 22.760 111.200 24.160 ;
        RECT 0.985 22.120 111.600 22.760 ;
        RECT 0.985 20.720 111.200 22.120 ;
        RECT 0.985 19.400 111.600 20.720 ;
        RECT 0.985 18.000 111.200 19.400 ;
        RECT 0.985 17.360 111.600 18.000 ;
        RECT 0.985 15.960 111.200 17.360 ;
        RECT 0.985 15.320 111.600 15.960 ;
        RECT 0.985 13.920 111.200 15.320 ;
        RECT 0.985 12.600 111.600 13.920 ;
        RECT 0.985 11.200 111.200 12.600 ;
        RECT 0.985 10.560 111.600 11.200 ;
        RECT 0.985 9.160 111.200 10.560 ;
        RECT 0.985 8.520 111.600 9.160 ;
        RECT 0.985 7.120 111.200 8.520 ;
        RECT 0.985 5.800 111.600 7.120 ;
        RECT 0.985 4.400 111.200 5.800 ;
        RECT 0.985 3.760 111.600 4.400 ;
        RECT 0.985 2.360 111.200 3.760 ;
        RECT 0.985 1.720 111.600 2.360 ;
        RECT 0.985 0.855 111.200 1.720 ;
      LAYER met4 ;
        RECT 56.200 9.695 100.905 100.880 ;
  END
END sb_0__2_
END LIBRARY

