VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO grid_clb
  CLASS BLOCK ;
  FOREIGN grid_clb ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN Test_en
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 2.400 ;
    END
  END Test_en
  PIN bottom_width_0_height_0__pin_16_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 2.400 ;
    END
  END bottom_width_0_height_0__pin_16_
  PIN bottom_width_0_height_0__pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END bottom_width_0_height_0__pin_17_
  PIN bottom_width_0_height_0__pin_18_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.400 ;
    END
  END bottom_width_0_height_0__pin_18_
  PIN bottom_width_0_height_0__pin_19_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 2.400 ;
    END
  END bottom_width_0_height_0__pin_19_
  PIN bottom_width_0_height_0__pin_20_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 2.400 ;
    END
  END bottom_width_0_height_0__pin_20_
  PIN bottom_width_0_height_0__pin_21_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 2.400 ;
    END
  END bottom_width_0_height_0__pin_21_
  PIN bottom_width_0_height_0__pin_22_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END bottom_width_0_height_0__pin_22_
  PIN bottom_width_0_height_0__pin_23_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 2.400 ;
    END
  END bottom_width_0_height_0__pin_23_
  PIN bottom_width_0_height_0__pin_24_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END bottom_width_0_height_0__pin_24_
  PIN bottom_width_0_height_0__pin_25_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 2.400 ;
    END
  END bottom_width_0_height_0__pin_25_
  PIN bottom_width_0_height_0__pin_26_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.400 ;
    END
  END bottom_width_0_height_0__pin_26_
  PIN bottom_width_0_height_0__pin_27_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END bottom_width_0_height_0__pin_27_
  PIN bottom_width_0_height_0__pin_28_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 2.400 ;
    END
  END bottom_width_0_height_0__pin_28_
  PIN bottom_width_0_height_0__pin_29_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 2.400 ;
    END
  END bottom_width_0_height_0__pin_29_
  PIN bottom_width_0_height_0__pin_30_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 2.400 ;
    END
  END bottom_width_0_height_0__pin_30_
  PIN bottom_width_0_height_0__pin_31_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.400 ;
    END
  END bottom_width_0_height_0__pin_31_
  PIN bottom_width_0_height_0__pin_42_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_lower
  PIN bottom_width_0_height_0__pin_42_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 2.400 ;
    END
  END bottom_width_0_height_0__pin_42_upper
  PIN bottom_width_0_height_0__pin_43_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_lower
  PIN bottom_width_0_height_0__pin_43_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.400 ;
    END
  END bottom_width_0_height_0__pin_43_upper
  PIN bottom_width_0_height_0__pin_44_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_lower
  PIN bottom_width_0_height_0__pin_44_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 2.400 ;
    END
  END bottom_width_0_height_0__pin_44_upper
  PIN bottom_width_0_height_0__pin_45_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_lower
  PIN bottom_width_0_height_0__pin_45_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 2.400 ;
    END
  END bottom_width_0_height_0__pin_45_upper
  PIN bottom_width_0_height_0__pin_46_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_lower
  PIN bottom_width_0_height_0__pin_46_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 2.400 ;
    END
  END bottom_width_0_height_0__pin_46_upper
  PIN bottom_width_0_height_0__pin_47_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_lower
  PIN bottom_width_0_height_0__pin_47_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 2.400 ;
    END
  END bottom_width_0_height_0__pin_47_upper
  PIN bottom_width_0_height_0__pin_48_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_lower
  PIN bottom_width_0_height_0__pin_48_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 2.400 ;
    END
  END bottom_width_0_height_0__pin_48_upper
  PIN bottom_width_0_height_0__pin_49_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.150 0.000 212.430 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_lower
  PIN bottom_width_0_height_0__pin_49_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.400 ;
    END
  END bottom_width_0_height_0__pin_49_upper
  PIN bottom_width_0_height_0__pin_50_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 2.400 ;
    END
  END bottom_width_0_height_0__pin_50_
  PIN bottom_width_0_height_0__pin_51_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 2.400 ;
    END
  END bottom_width_0_height_0__pin_51_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 2.400 188.320 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.010 247.600 208.290 250.000 ;
    END
  END ccff_tail
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END clk
  PIN left_width_0_height_0__pin_52_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 2.400 63.200 ;
    END
  END left_width_0_height_0__pin_52_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 2.400 ;
    END
  END prog_clk
  PIN right_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 3.440 250.000 4.040 ;
    END
  END right_width_0_height_0__pin_0_
  PIN right_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 81.640 250.000 82.240 ;
    END
  END right_width_0_height_0__pin_10_
  PIN right_width_0_height_0__pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 89.120 250.000 89.720 ;
    END
  END right_width_0_height_0__pin_11_
  PIN right_width_0_height_0__pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 97.280 250.000 97.880 ;
    END
  END right_width_0_height_0__pin_12_
  PIN right_width_0_height_0__pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 104.760 250.000 105.360 ;
    END
  END right_width_0_height_0__pin_13_
  PIN right_width_0_height_0__pin_14_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 112.920 250.000 113.520 ;
    END
  END right_width_0_height_0__pin_14_
  PIN right_width_0_height_0__pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 120.400 250.000 121.000 ;
    END
  END right_width_0_height_0__pin_15_
  PIN right_width_0_height_0__pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 10.920 250.000 11.520 ;
    END
  END right_width_0_height_0__pin_1_
  PIN right_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 19.080 250.000 19.680 ;
    END
  END right_width_0_height_0__pin_2_
  PIN right_width_0_height_0__pin_34_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 128.560 250.000 129.160 ;
    END
  END right_width_0_height_0__pin_34_lower
  PIN right_width_0_height_0__pin_34_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 136.040 250.000 136.640 ;
    END
  END right_width_0_height_0__pin_34_upper
  PIN right_width_0_height_0__pin_35_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 144.200 250.000 144.800 ;
    END
  END right_width_0_height_0__pin_35_lower
  PIN right_width_0_height_0__pin_35_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 151.680 250.000 152.280 ;
    END
  END right_width_0_height_0__pin_35_upper
  PIN right_width_0_height_0__pin_36_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 159.840 250.000 160.440 ;
    END
  END right_width_0_height_0__pin_36_lower
  PIN right_width_0_height_0__pin_36_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 167.320 250.000 167.920 ;
    END
  END right_width_0_height_0__pin_36_upper
  PIN right_width_0_height_0__pin_37_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 175.480 250.000 176.080 ;
    END
  END right_width_0_height_0__pin_37_lower
  PIN right_width_0_height_0__pin_37_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 182.960 250.000 183.560 ;
    END
  END right_width_0_height_0__pin_37_upper
  PIN right_width_0_height_0__pin_38_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 191.120 250.000 191.720 ;
    END
  END right_width_0_height_0__pin_38_lower
  PIN right_width_0_height_0__pin_38_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 198.600 250.000 199.200 ;
    END
  END right_width_0_height_0__pin_38_upper
  PIN right_width_0_height_0__pin_39_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 206.760 250.000 207.360 ;
    END
  END right_width_0_height_0__pin_39_lower
  PIN right_width_0_height_0__pin_39_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 214.240 250.000 214.840 ;
    END
  END right_width_0_height_0__pin_39_upper
  PIN right_width_0_height_0__pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 26.560 250.000 27.160 ;
    END
  END right_width_0_height_0__pin_3_
  PIN right_width_0_height_0__pin_40_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 222.400 250.000 223.000 ;
    END
  END right_width_0_height_0__pin_40_lower
  PIN right_width_0_height_0__pin_40_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 229.880 250.000 230.480 ;
    END
  END right_width_0_height_0__pin_40_upper
  PIN right_width_0_height_0__pin_41_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 238.040 250.000 238.640 ;
    END
  END right_width_0_height_0__pin_41_lower
  PIN right_width_0_height_0__pin_41_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 247.600 245.520 250.000 246.120 ;
    END
  END right_width_0_height_0__pin_41_upper
  PIN right_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 34.720 250.000 35.320 ;
    END
  END right_width_0_height_0__pin_4_
  PIN right_width_0_height_0__pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 42.200 250.000 42.800 ;
    END
  END right_width_0_height_0__pin_5_
  PIN right_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 50.360 250.000 50.960 ;
    END
  END right_width_0_height_0__pin_6_
  PIN right_width_0_height_0__pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 57.840 250.000 58.440 ;
    END
  END right_width_0_height_0__pin_7_
  PIN right_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 66.000 250.000 66.600 ;
    END
  END right_width_0_height_0__pin_8_
  PIN right_width_0_height_0__pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 247.600 73.480 250.000 74.080 ;
    END
  END right_width_0_height_0__pin_9_
  PIN top_width_0_height_0__pin_32_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.490 247.600 41.770 250.000 ;
    END
  END top_width_0_height_0__pin_32_
  PIN top_width_0_height_0__pin_33_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.750 247.600 125.030 250.000 ;
    END
  END top_width_0_height_0__pin_33_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 236.880 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 236.880 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 244.260 236.725 ;
      LAYER met1 ;
        RECT 5.520 2.760 244.260 236.880 ;
      LAYER met2 ;
        RECT 3.310 247.320 41.210 247.600 ;
        RECT 42.050 247.320 124.470 247.600 ;
        RECT 125.310 247.320 207.730 247.600 ;
        RECT 208.570 247.320 246.470 247.600 ;
        RECT 3.310 2.680 246.470 247.320 ;
        RECT 3.870 0.155 9.470 2.680 ;
        RECT 10.310 0.155 16.370 2.680 ;
        RECT 17.210 0.155 23.270 2.680 ;
        RECT 24.110 0.155 29.710 2.680 ;
        RECT 30.550 0.155 36.610 2.680 ;
        RECT 37.450 0.155 43.510 2.680 ;
        RECT 44.350 0.155 49.950 2.680 ;
        RECT 50.790 0.155 56.850 2.680 ;
        RECT 57.690 0.155 63.750 2.680 ;
        RECT 64.590 0.155 70.190 2.680 ;
        RECT 71.030 0.155 77.090 2.680 ;
        RECT 77.930 0.155 83.990 2.680 ;
        RECT 84.830 0.155 90.430 2.680 ;
        RECT 91.270 0.155 97.330 2.680 ;
        RECT 98.170 0.155 104.230 2.680 ;
        RECT 105.070 0.155 110.670 2.680 ;
        RECT 111.510 0.155 117.570 2.680 ;
        RECT 118.410 0.155 124.470 2.680 ;
        RECT 125.310 0.155 130.910 2.680 ;
        RECT 131.750 0.155 137.810 2.680 ;
        RECT 138.650 0.155 144.710 2.680 ;
        RECT 145.550 0.155 151.150 2.680 ;
        RECT 151.990 0.155 158.050 2.680 ;
        RECT 158.890 0.155 164.950 2.680 ;
        RECT 165.790 0.155 171.390 2.680 ;
        RECT 172.230 0.155 178.290 2.680 ;
        RECT 179.130 0.155 185.190 2.680 ;
        RECT 186.030 0.155 191.630 2.680 ;
        RECT 192.470 0.155 198.530 2.680 ;
        RECT 199.370 0.155 205.430 2.680 ;
        RECT 206.270 0.155 211.870 2.680 ;
        RECT 212.710 0.155 218.770 2.680 ;
        RECT 219.610 0.155 225.670 2.680 ;
        RECT 226.510 0.155 232.110 2.680 ;
        RECT 232.950 0.155 239.010 2.680 ;
        RECT 239.850 0.155 245.910 2.680 ;
      LAYER met3 ;
        RECT 2.400 245.120 247.200 245.985 ;
        RECT 2.400 239.040 247.600 245.120 ;
        RECT 2.400 237.640 247.200 239.040 ;
        RECT 2.400 230.880 247.600 237.640 ;
        RECT 2.400 229.480 247.200 230.880 ;
        RECT 2.400 223.400 247.600 229.480 ;
        RECT 2.400 222.000 247.200 223.400 ;
        RECT 2.400 215.240 247.600 222.000 ;
        RECT 2.400 213.840 247.200 215.240 ;
        RECT 2.400 207.760 247.600 213.840 ;
        RECT 2.400 206.360 247.200 207.760 ;
        RECT 2.400 199.600 247.600 206.360 ;
        RECT 2.400 198.200 247.200 199.600 ;
        RECT 2.400 192.120 247.600 198.200 ;
        RECT 2.400 190.720 247.200 192.120 ;
        RECT 2.400 188.720 247.600 190.720 ;
        RECT 2.800 187.320 247.600 188.720 ;
        RECT 2.400 183.960 247.600 187.320 ;
        RECT 2.400 182.560 247.200 183.960 ;
        RECT 2.400 176.480 247.600 182.560 ;
        RECT 2.400 175.080 247.200 176.480 ;
        RECT 2.400 168.320 247.600 175.080 ;
        RECT 2.400 166.920 247.200 168.320 ;
        RECT 2.400 160.840 247.600 166.920 ;
        RECT 2.400 159.440 247.200 160.840 ;
        RECT 2.400 152.680 247.600 159.440 ;
        RECT 2.400 151.280 247.200 152.680 ;
        RECT 2.400 145.200 247.600 151.280 ;
        RECT 2.400 143.800 247.200 145.200 ;
        RECT 2.400 137.040 247.600 143.800 ;
        RECT 2.400 135.640 247.200 137.040 ;
        RECT 2.400 129.560 247.600 135.640 ;
        RECT 2.400 128.160 247.200 129.560 ;
        RECT 2.400 121.400 247.600 128.160 ;
        RECT 2.400 120.000 247.200 121.400 ;
        RECT 2.400 113.920 247.600 120.000 ;
        RECT 2.400 112.520 247.200 113.920 ;
        RECT 2.400 105.760 247.600 112.520 ;
        RECT 2.400 104.360 247.200 105.760 ;
        RECT 2.400 98.280 247.600 104.360 ;
        RECT 2.400 96.880 247.200 98.280 ;
        RECT 2.400 90.120 247.600 96.880 ;
        RECT 2.400 88.720 247.200 90.120 ;
        RECT 2.400 82.640 247.600 88.720 ;
        RECT 2.400 81.240 247.200 82.640 ;
        RECT 2.400 74.480 247.600 81.240 ;
        RECT 2.400 73.080 247.200 74.480 ;
        RECT 2.400 67.000 247.600 73.080 ;
        RECT 2.400 65.600 247.200 67.000 ;
        RECT 2.400 63.600 247.600 65.600 ;
        RECT 2.800 62.200 247.600 63.600 ;
        RECT 2.400 58.840 247.600 62.200 ;
        RECT 2.400 57.440 247.200 58.840 ;
        RECT 2.400 51.360 247.600 57.440 ;
        RECT 2.400 49.960 247.200 51.360 ;
        RECT 2.400 43.200 247.600 49.960 ;
        RECT 2.400 41.800 247.200 43.200 ;
        RECT 2.400 35.720 247.600 41.800 ;
        RECT 2.400 34.320 247.200 35.720 ;
        RECT 2.400 27.560 247.600 34.320 ;
        RECT 2.400 26.160 247.200 27.560 ;
        RECT 2.400 20.080 247.600 26.160 ;
        RECT 2.400 18.680 247.200 20.080 ;
        RECT 2.400 11.920 247.600 18.680 ;
        RECT 2.400 10.520 247.200 11.920 ;
        RECT 2.400 4.440 247.600 10.520 ;
        RECT 2.400 3.040 247.200 4.440 ;
        RECT 2.400 0.175 247.600 3.040 ;
      LAYER met4 ;
        RECT 3.550 10.640 20.640 236.880 ;
        RECT 23.040 10.640 97.440 236.880 ;
        RECT 99.840 10.640 176.240 236.880 ;
      LAYER met5 ;
        RECT 3.340 14.500 155.820 19.500 ;
  END
END grid_clb
END LIBRARY

