VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.800 140.000 5.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 14.320 140.000 14.920 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END address[5]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 2.400 15.600 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 2.400 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 137.600 4.970 140.000 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 137.600 14.170 140.000 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 2.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 24.520 140.000 25.120 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 137.600 23.370 140.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 137.600 32.570 140.000 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 2.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.400 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 34.720 140.000 35.320 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.400 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 2.400 48.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_right_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 137.600 42.230 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 137.600 51.430 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 54.440 140.000 55.040 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.350 137.600 60.630 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 64.640 140.000 65.240 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 137.600 79.490 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 2.400 91.080 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 2.400 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 137.600 88.690 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 74.840 140.000 75.440 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 2.400 ;
    END
  END enable
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.760 140.000 105.360 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.280 140.000 114.880 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.470 137.600 116.750 140.000 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 84.360 140.000 84.960 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.810 137.600 107.090 140.000 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 94.560 140.000 95.160 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 2.400 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 2.400 ;
    END
  END right_bottom_grid_pin_9_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 2.400 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END top_left_grid_pin_11_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 2.400 123.720 ;
    END
  END top_left_grid_pin_13_
  PIN top_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.870 137.600 135.150 140.000 ;
    END
  END top_left_grid_pin_15_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.670 137.600 125.950 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN top_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 124.480 140.000 125.080 ;
    END
  END top_left_grid_pin_3_
  PIN top_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END top_left_grid_pin_5_
  PIN top_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 134.680 140.000 135.280 ;
    END
  END top_left_grid_pin_7_
  PIN top_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END top_left_grid_pin_9_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 2.400 134.600 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 10.640 138.390 137.660 ;
      LAYER met2 ;
        RECT 0.550 137.320 4.410 137.770 ;
        RECT 5.250 137.320 13.610 137.770 ;
        RECT 14.450 137.320 22.810 137.770 ;
        RECT 23.650 137.320 32.010 137.770 ;
        RECT 32.850 137.320 41.670 137.770 ;
        RECT 42.510 137.320 50.870 137.770 ;
        RECT 51.710 137.320 60.070 137.770 ;
        RECT 60.910 137.320 69.270 137.770 ;
        RECT 70.110 137.320 78.930 137.770 ;
        RECT 79.770 137.320 88.130 137.770 ;
        RECT 88.970 137.320 97.330 137.770 ;
        RECT 98.170 137.320 106.530 137.770 ;
        RECT 107.370 137.320 116.190 137.770 ;
        RECT 117.030 137.320 125.390 137.770 ;
        RECT 126.230 137.320 134.590 137.770 ;
        RECT 135.430 137.320 138.370 137.770 ;
        RECT 0.550 2.680 138.370 137.320 ;
        RECT 0.550 0.155 3.030 2.680 ;
        RECT 3.870 0.155 9.930 2.680 ;
        RECT 10.770 0.155 16.830 2.680 ;
        RECT 17.670 0.155 23.730 2.680 ;
        RECT 24.570 0.155 30.630 2.680 ;
        RECT 31.470 0.155 37.990 2.680 ;
        RECT 38.830 0.155 44.890 2.680 ;
        RECT 45.730 0.155 51.790 2.680 ;
        RECT 52.630 0.155 58.690 2.680 ;
        RECT 59.530 0.155 65.590 2.680 ;
        RECT 66.430 0.155 72.950 2.680 ;
        RECT 73.790 0.155 79.850 2.680 ;
        RECT 80.690 0.155 86.750 2.680 ;
        RECT 87.590 0.155 93.650 2.680 ;
        RECT 94.490 0.155 100.550 2.680 ;
        RECT 101.390 0.155 107.910 2.680 ;
        RECT 108.750 0.155 114.810 2.680 ;
        RECT 115.650 0.155 121.710 2.680 ;
        RECT 122.550 0.155 128.610 2.680 ;
        RECT 129.450 0.155 135.510 2.680 ;
        RECT 136.350 0.155 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 134.280 137.200 134.680 ;
        RECT 2.800 133.600 138.610 134.280 ;
        RECT 0.310 125.480 138.610 133.600 ;
        RECT 0.310 124.120 137.200 125.480 ;
        RECT 2.800 124.080 137.200 124.120 ;
        RECT 2.800 122.720 138.610 124.080 ;
        RECT 0.310 115.280 138.610 122.720 ;
        RECT 0.310 113.880 137.200 115.280 ;
        RECT 0.310 113.240 138.610 113.880 ;
        RECT 2.800 111.840 138.610 113.240 ;
        RECT 0.310 105.760 138.610 111.840 ;
        RECT 0.310 104.360 137.200 105.760 ;
        RECT 0.310 102.360 138.610 104.360 ;
        RECT 2.800 100.960 138.610 102.360 ;
        RECT 0.310 95.560 138.610 100.960 ;
        RECT 0.310 94.160 137.200 95.560 ;
        RECT 0.310 91.480 138.610 94.160 ;
        RECT 2.800 90.080 138.610 91.480 ;
        RECT 0.310 85.360 138.610 90.080 ;
        RECT 0.310 83.960 137.200 85.360 ;
        RECT 0.310 80.600 138.610 83.960 ;
        RECT 2.800 79.200 138.610 80.600 ;
        RECT 0.310 75.840 138.610 79.200 ;
        RECT 0.310 74.440 137.200 75.840 ;
        RECT 0.310 70.400 138.610 74.440 ;
        RECT 2.800 69.000 138.610 70.400 ;
        RECT 0.310 65.640 138.610 69.000 ;
        RECT 0.310 64.240 137.200 65.640 ;
        RECT 0.310 59.520 138.610 64.240 ;
        RECT 2.800 58.120 138.610 59.520 ;
        RECT 0.310 55.440 138.610 58.120 ;
        RECT 0.310 54.040 137.200 55.440 ;
        RECT 0.310 48.640 138.610 54.040 ;
        RECT 2.800 47.240 138.610 48.640 ;
        RECT 0.310 45.240 138.610 47.240 ;
        RECT 0.310 43.840 137.200 45.240 ;
        RECT 0.310 37.760 138.610 43.840 ;
        RECT 2.800 36.360 138.610 37.760 ;
        RECT 0.310 35.720 138.610 36.360 ;
        RECT 0.310 34.320 137.200 35.720 ;
        RECT 0.310 26.880 138.610 34.320 ;
        RECT 2.800 25.520 138.610 26.880 ;
        RECT 2.800 25.480 137.200 25.520 ;
        RECT 0.310 24.120 137.200 25.480 ;
        RECT 0.310 16.000 138.610 24.120 ;
        RECT 2.800 15.320 138.610 16.000 ;
        RECT 2.800 14.600 137.200 15.320 ;
        RECT 0.310 13.920 137.200 14.600 ;
        RECT 0.310 5.800 138.610 13.920 ;
        RECT 2.800 4.400 137.200 5.800 ;
        RECT 0.310 0.175 138.610 4.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_0__0_
END LIBRARY

