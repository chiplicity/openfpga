magic
tech sky130A
magscale 1 2
timestamp 1605198049
<< locali >>
rect 6837 19771 6871 20009
rect 12449 13719 12483 13821
<< viali >>
rect 1961 20553 1995 20587
rect 3065 20553 3099 20587
rect 4629 20485 4663 20519
rect 6929 20485 6963 20519
rect 13829 20485 13863 20519
rect 5089 20417 5123 20451
rect 5181 20417 5215 20451
rect 7481 20417 7515 20451
rect 11253 20417 11287 20451
rect 14473 20417 14507 20451
rect 16037 20417 16071 20451
rect 18521 20417 18555 20451
rect 19901 20417 19935 20451
rect 1777 20349 1811 20383
rect 2881 20349 2915 20383
rect 7389 20349 7423 20383
rect 8585 20349 8619 20383
rect 9781 20349 9815 20383
rect 11069 20349 11103 20383
rect 12725 20349 12759 20383
rect 17141 20349 17175 20383
rect 18337 20349 18371 20383
rect 19717 20349 19751 20383
rect 7297 20281 7331 20315
rect 10057 20281 10091 20315
rect 14197 20281 14231 20315
rect 4997 20213 5031 20247
rect 8769 20213 8803 20247
rect 12909 20213 12943 20247
rect 14289 20213 14323 20247
rect 15485 20213 15519 20247
rect 15853 20213 15887 20247
rect 15945 20213 15979 20247
rect 17325 20213 17359 20247
rect 1961 20009 1995 20043
rect 3065 20009 3099 20043
rect 6837 20009 6871 20043
rect 13185 20009 13219 20043
rect 4528 19941 4562 19975
rect 1777 19873 1811 19907
rect 2881 19873 2915 19907
rect 4261 19805 4295 19839
rect 9956 19941 9990 19975
rect 7185 19873 7219 19907
rect 15669 19873 15703 19907
rect 16865 19873 16899 19907
rect 18153 19873 18187 19907
rect 19533 19873 19567 19907
rect 6929 19805 6963 19839
rect 9696 19805 9730 19839
rect 13277 19805 13311 19839
rect 13461 19805 13495 19839
rect 15761 19805 15795 19839
rect 15945 19805 15979 19839
rect 17049 19805 17083 19839
rect 18337 19805 18371 19839
rect 19717 19805 19751 19839
rect 6837 19737 6871 19771
rect 5641 19669 5675 19703
rect 8309 19669 8343 19703
rect 11069 19669 11103 19703
rect 12817 19669 12851 19703
rect 15301 19669 15335 19703
rect 19625 19465 19659 19499
rect 4813 19397 4847 19431
rect 10977 19329 11011 19363
rect 20177 19329 20211 19363
rect 2329 19261 2363 19295
rect 3433 19261 3467 19295
rect 5641 19261 5675 19295
rect 6837 19261 6871 19295
rect 8125 19261 8159 19295
rect 8392 19261 8426 19295
rect 10701 19261 10735 19295
rect 13185 19261 13219 19295
rect 15393 19261 15427 19295
rect 18061 19261 18095 19295
rect 3700 19193 3734 19227
rect 7113 19193 7147 19227
rect 10793 19193 10827 19227
rect 13452 19193 13486 19227
rect 15638 19193 15672 19227
rect 18337 19193 18371 19227
rect 19993 19193 20027 19227
rect 2513 19125 2547 19159
rect 5825 19125 5859 19159
rect 9505 19125 9539 19159
rect 10333 19125 10367 19159
rect 14565 19125 14599 19159
rect 16773 19125 16807 19159
rect 20085 19125 20119 19159
rect 3065 18921 3099 18955
rect 13921 18921 13955 18955
rect 5702 18853 5736 18887
rect 8401 18853 8435 18887
rect 10600 18853 10634 18887
rect 15301 18853 15335 18887
rect 16580 18853 16614 18887
rect 1777 18785 1811 18819
rect 2881 18785 2915 18819
rect 4169 18785 4203 18819
rect 12797 18785 12831 18819
rect 18889 18785 18923 18819
rect 4445 18717 4479 18751
rect 5457 18717 5491 18751
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 10333 18717 10367 18751
rect 12541 18717 12575 18751
rect 16313 18717 16347 18751
rect 18981 18717 19015 18751
rect 19165 18717 19199 18751
rect 1961 18649 1995 18683
rect 6837 18649 6871 18683
rect 11713 18649 11747 18683
rect 17693 18649 17727 18683
rect 8033 18581 8067 18615
rect 18337 18581 18371 18615
rect 18521 18581 18555 18615
rect 6837 18377 6871 18411
rect 10793 18377 10827 18411
rect 13737 18309 13771 18343
rect 5733 18241 5767 18275
rect 7389 18241 7423 18275
rect 9137 18241 9171 18275
rect 9229 18241 9263 18275
rect 11437 18241 11471 18275
rect 14197 18241 14231 18275
rect 14381 18241 14415 18275
rect 15761 18241 15795 18275
rect 15945 18241 15979 18275
rect 20453 18241 20487 18275
rect 1409 18173 1443 18207
rect 2513 18173 2547 18207
rect 5549 18173 5583 18207
rect 7205 18173 7239 18207
rect 11161 18173 11195 18207
rect 11253 18173 11287 18207
rect 12449 18173 12483 18207
rect 15669 18173 15703 18207
rect 16865 18173 16899 18207
rect 18061 18173 18095 18207
rect 18328 18173 18362 18207
rect 20269 18173 20303 18207
rect 2780 18105 2814 18139
rect 9045 18105 9079 18139
rect 12725 18105 12759 18139
rect 14105 18105 14139 18139
rect 1593 18037 1627 18071
rect 3893 18037 3927 18071
rect 5181 18037 5215 18071
rect 5641 18037 5675 18071
rect 7297 18037 7331 18071
rect 8677 18037 8711 18071
rect 15301 18037 15335 18071
rect 17049 18037 17083 18071
rect 19441 18037 19475 18071
rect 2881 17833 2915 17867
rect 6193 17833 6227 17867
rect 12357 17833 12391 17867
rect 18429 17833 18463 17867
rect 18797 17833 18831 17867
rect 9965 17765 9999 17799
rect 2789 17697 2823 17731
rect 4905 17697 4939 17731
rect 6561 17697 6595 17731
rect 8217 17697 8251 17731
rect 9689 17697 9723 17731
rect 11244 17697 11278 17731
rect 14013 17697 14047 17731
rect 16396 17697 16430 17731
rect 1409 17629 1443 17663
rect 3065 17629 3099 17663
rect 4997 17629 5031 17663
rect 5089 17629 5123 17663
rect 6653 17629 6687 17663
rect 6745 17629 6779 17663
rect 8309 17629 8343 17663
rect 8401 17629 8435 17663
rect 10977 17629 11011 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 16129 17629 16163 17663
rect 18889 17629 18923 17663
rect 18981 17629 19015 17663
rect 17509 17561 17543 17595
rect 2421 17493 2455 17527
rect 4537 17493 4571 17527
rect 7849 17493 7883 17527
rect 13645 17493 13679 17527
rect 3709 17289 3743 17323
rect 6837 17289 6871 17323
rect 9965 17289 9999 17323
rect 15117 17289 15151 17323
rect 19625 17289 19659 17323
rect 10793 17221 10827 17255
rect 14197 17221 14231 17255
rect 5089 17153 5123 17187
rect 7481 17153 7515 17187
rect 8585 17153 8619 17187
rect 11437 17153 11471 17187
rect 13001 17153 13035 17187
rect 15669 17153 15703 17187
rect 18613 17153 18647 17187
rect 20177 17153 20211 17187
rect 2329 17085 2363 17119
rect 2596 17085 2630 17119
rect 4905 17085 4939 17119
rect 7205 17085 7239 17119
rect 12817 17085 12851 17119
rect 14013 17085 14047 17119
rect 16681 17085 16715 17119
rect 18429 17085 18463 17119
rect 18889 17085 18923 17119
rect 20085 17085 20119 17119
rect 8852 17017 8886 17051
rect 11161 17017 11195 17051
rect 16957 17017 16991 17051
rect 18521 17017 18555 17051
rect 19993 17017 20027 17051
rect 4537 16949 4571 16983
rect 4997 16949 5031 16983
rect 7297 16949 7331 16983
rect 11253 16949 11287 16983
rect 12449 16949 12483 16983
rect 12909 16949 12943 16983
rect 15485 16949 15519 16983
rect 15577 16949 15611 16983
rect 18061 16949 18095 16983
rect 1777 16745 1811 16779
rect 4537 16745 4571 16779
rect 11253 16745 11287 16779
rect 11713 16745 11747 16779
rect 14381 16745 14415 16779
rect 19073 16745 19107 16779
rect 2973 16677 3007 16711
rect 4629 16677 4663 16711
rect 16764 16677 16798 16711
rect 1593 16609 1627 16643
rect 2697 16609 2731 16643
rect 6920 16609 6954 16643
rect 10057 16609 10091 16643
rect 10149 16609 10183 16643
rect 11621 16609 11655 16643
rect 13001 16609 13035 16643
rect 13268 16609 13302 16643
rect 15393 16609 15427 16643
rect 4813 16541 4847 16575
rect 6653 16541 6687 16575
rect 10241 16541 10275 16575
rect 11805 16541 11839 16575
rect 16497 16541 16531 16575
rect 19165 16541 19199 16575
rect 19257 16541 19291 16575
rect 4169 16473 4203 16507
rect 15577 16473 15611 16507
rect 18705 16473 18739 16507
rect 8033 16405 8067 16439
rect 9689 16405 9723 16439
rect 17877 16405 17911 16439
rect 5181 16201 5215 16235
rect 12633 16201 12667 16235
rect 15577 16201 15611 16235
rect 18061 16201 18095 16235
rect 19901 16201 19935 16235
rect 9045 16133 9079 16167
rect 4077 16065 4111 16099
rect 4261 16065 4295 16099
rect 5825 16065 5859 16099
rect 7389 16065 7423 16099
rect 9505 16065 9539 16099
rect 9597 16065 9631 16099
rect 11437 16065 11471 16099
rect 13277 16065 13311 16099
rect 14197 16065 14231 16099
rect 16957 16065 16991 16099
rect 18613 16065 18647 16099
rect 20453 16065 20487 16099
rect 2329 15997 2363 16031
rect 3985 15997 4019 16031
rect 5549 15997 5583 16031
rect 8585 15997 8619 16031
rect 9413 15997 9447 16031
rect 16865 15997 16899 16031
rect 18521 15997 18555 16031
rect 2605 15929 2639 15963
rect 7297 15929 7331 15963
rect 11161 15929 11195 15963
rect 13001 15929 13035 15963
rect 14464 15929 14498 15963
rect 18429 15929 18463 15963
rect 20361 15929 20395 15963
rect 3617 15861 3651 15895
rect 5641 15861 5675 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 8401 15861 8435 15895
rect 10793 15861 10827 15895
rect 11253 15861 11287 15895
rect 13093 15861 13127 15895
rect 16405 15861 16439 15895
rect 16773 15861 16807 15895
rect 19809 15861 19843 15895
rect 20269 15861 20303 15895
rect 1777 15657 1811 15691
rect 7297 15657 7331 15691
rect 10609 15657 10643 15691
rect 2973 15589 3007 15623
rect 4721 15589 4755 15623
rect 6184 15589 6218 15623
rect 8585 15589 8619 15623
rect 16313 15589 16347 15623
rect 1593 15521 1627 15555
rect 2697 15521 2731 15555
rect 4813 15521 4847 15555
rect 5917 15521 5951 15555
rect 8309 15521 8343 15555
rect 10517 15521 10551 15555
rect 12061 15521 12095 15555
rect 14105 15521 14139 15555
rect 17776 15521 17810 15555
rect 19717 15521 19751 15555
rect 4997 15453 5031 15487
rect 10701 15453 10735 15487
rect 11805 15453 11839 15487
rect 16405 15453 16439 15487
rect 16497 15453 16531 15487
rect 17509 15453 17543 15487
rect 10149 15385 10183 15419
rect 14289 15385 14323 15419
rect 4353 15317 4387 15351
rect 13185 15317 13219 15351
rect 15945 15317 15979 15351
rect 18889 15317 18923 15351
rect 19901 15317 19935 15351
rect 5089 15113 5123 15147
rect 6377 15113 6411 15147
rect 7665 15113 7699 15147
rect 13829 15113 13863 15147
rect 14657 15113 14691 15147
rect 16221 15113 16255 15147
rect 19993 15113 20027 15147
rect 10609 15045 10643 15079
rect 2789 14977 2823 15011
rect 8309 14977 8343 15011
rect 15301 14977 15335 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 2513 14909 2547 14943
rect 3709 14909 3743 14943
rect 6561 14909 6595 14943
rect 9229 14909 9263 14943
rect 12265 14909 12299 14943
rect 12449 14909 12483 14943
rect 15025 14909 15059 14943
rect 16589 14909 16623 14943
rect 18613 14909 18647 14943
rect 18880 14909 18914 14943
rect 3976 14841 4010 14875
rect 8125 14841 8159 14875
rect 9496 14841 9530 14875
rect 12716 14841 12750 14875
rect 15117 14841 15151 14875
rect 2145 14773 2179 14807
rect 2605 14773 2639 14807
rect 8033 14773 8067 14807
rect 12081 14773 12115 14807
rect 3065 14569 3099 14603
rect 7481 14569 7515 14603
rect 8585 14569 8619 14603
rect 10057 14569 10091 14603
rect 11621 14569 11655 14603
rect 17601 14569 17635 14603
rect 5080 14501 5114 14535
rect 10425 14501 10459 14535
rect 16466 14501 16500 14535
rect 1777 14433 1811 14467
rect 2881 14433 2915 14467
rect 7389 14433 7423 14467
rect 11989 14433 12023 14467
rect 13553 14433 13587 14467
rect 13645 14433 13679 14467
rect 15117 14433 15151 14467
rect 16221 14433 16255 14467
rect 19625 14433 19659 14467
rect 4813 14365 4847 14399
rect 7665 14365 7699 14399
rect 10517 14365 10551 14399
rect 10701 14365 10735 14399
rect 12081 14365 12115 14399
rect 12265 14365 12299 14399
rect 13737 14365 13771 14399
rect 19717 14365 19751 14399
rect 19901 14365 19935 14399
rect 1961 14297 1995 14331
rect 13185 14297 13219 14331
rect 14933 14297 14967 14331
rect 6193 14229 6227 14263
rect 7021 14229 7055 14263
rect 9965 14229 9999 14263
rect 19257 14229 19291 14263
rect 10793 14025 10827 14059
rect 14381 14025 14415 14059
rect 19809 14025 19843 14059
rect 1869 13957 1903 13991
rect 4169 13957 4203 13991
rect 7297 13957 7331 13991
rect 16681 13957 16715 13991
rect 5549 13889 5583 13923
rect 7849 13889 7883 13923
rect 9689 13889 9723 13923
rect 11345 13889 11379 13923
rect 13185 13889 13219 13923
rect 18797 13889 18831 13923
rect 20361 13889 20395 13923
rect 1685 13821 1719 13855
rect 2789 13821 2823 13855
rect 5457 13821 5491 13855
rect 7757 13821 7791 13855
rect 9413 13821 9447 13855
rect 11253 13821 11287 13855
rect 12449 13821 12483 13855
rect 13001 13821 13035 13855
rect 14197 13821 14231 13855
rect 15301 13821 15335 13855
rect 15557 13821 15591 13855
rect 18705 13821 18739 13855
rect 20269 13821 20303 13855
rect 3056 13753 3090 13787
rect 5365 13753 5399 13787
rect 7665 13753 7699 13787
rect 9505 13753 9539 13787
rect 18613 13753 18647 13787
rect 4997 13685 5031 13719
rect 9045 13685 9079 13719
rect 11161 13685 11195 13719
rect 12449 13685 12483 13719
rect 12541 13685 12575 13719
rect 12909 13685 12943 13719
rect 18245 13685 18279 13719
rect 20177 13685 20211 13719
rect 1409 13481 1443 13515
rect 2789 13481 2823 13515
rect 8401 13481 8435 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 10149 13481 10183 13515
rect 11529 13481 11563 13515
rect 13829 13481 13863 13515
rect 14657 13481 14691 13515
rect 18061 13481 18095 13515
rect 19257 13481 19291 13515
rect 15761 13413 15795 13447
rect 4169 13345 4203 13379
rect 5457 13345 5491 13379
rect 5724 13345 5758 13379
rect 7941 13345 7975 13379
rect 11345 13345 11379 13379
rect 12705 13345 12739 13379
rect 14841 13345 14875 13379
rect 15669 13345 15703 13379
rect 19625 13345 19659 13379
rect 2881 13277 2915 13311
rect 3065 13277 3099 13311
rect 4445 13277 4479 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 10241 13277 10275 13311
rect 12449 13277 12483 13311
rect 15853 13277 15887 13311
rect 18153 13277 18187 13311
rect 18337 13277 18371 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 7757 13209 7791 13243
rect 2421 13141 2455 13175
rect 6837 13141 6871 13175
rect 8033 13141 8067 13175
rect 15301 13141 15335 13175
rect 17693 13141 17727 13175
rect 1593 12937 1627 12971
rect 6837 12937 6871 12971
rect 12725 12937 12759 12971
rect 15025 12937 15059 12971
rect 16405 12937 16439 12971
rect 20361 12937 20395 12971
rect 3893 12869 3927 12903
rect 8401 12869 8435 12903
rect 5181 12801 5215 12835
rect 5273 12801 5307 12835
rect 7481 12801 7515 12835
rect 8953 12801 8987 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 13645 12801 13679 12835
rect 17049 12801 17083 12835
rect 1409 12733 1443 12767
rect 2513 12733 2547 12767
rect 2780 12733 2814 12767
rect 12541 12733 12575 12767
rect 16773 12733 16807 12767
rect 18981 12733 19015 12767
rect 19237 12733 19271 12767
rect 13890 12665 13924 12699
rect 4721 12597 4755 12631
rect 5089 12597 5123 12631
rect 7205 12597 7239 12631
rect 7297 12597 7331 12631
rect 8769 12597 8803 12631
rect 8861 12597 8895 12631
rect 9965 12597 9999 12631
rect 10333 12597 10367 12631
rect 16865 12597 16899 12631
rect 4261 12393 4295 12427
rect 8125 12393 8159 12427
rect 13645 12393 13679 12427
rect 15301 12393 15335 12427
rect 16313 12393 16347 12427
rect 16681 12393 16715 12427
rect 19257 12393 19291 12427
rect 1869 12325 1903 12359
rect 4629 12325 4663 12359
rect 4721 12325 4755 12359
rect 9965 12325 9999 12359
rect 2881 12257 2915 12291
rect 6745 12257 6779 12291
rect 7012 12257 7046 12291
rect 9137 12257 9171 12291
rect 9689 12257 9723 12291
rect 10977 12257 11011 12291
rect 11244 12257 11278 12291
rect 13553 12257 13587 12291
rect 14933 12257 14967 12291
rect 17877 12257 17911 12291
rect 18133 12257 18167 12291
rect 4813 12189 4847 12223
rect 13737 12189 13771 12223
rect 16773 12189 16807 12223
rect 16957 12189 16991 12223
rect 3065 12121 3099 12155
rect 12357 12121 12391 12155
rect 13185 12121 13219 12155
rect 8953 12053 8987 12087
rect 14749 12053 14783 12087
rect 3525 11849 3559 11883
rect 5089 11849 5123 11883
rect 8217 11849 8251 11883
rect 9045 11849 9079 11883
rect 10609 11849 10643 11883
rect 13185 11849 13219 11883
rect 14841 11849 14875 11883
rect 16405 11849 16439 11883
rect 20821 11849 20855 11883
rect 1501 11713 1535 11747
rect 2513 11713 2547 11747
rect 4077 11713 4111 11747
rect 5641 11713 5675 11747
rect 6837 11713 6871 11747
rect 9597 11713 9631 11747
rect 11161 11713 11195 11747
rect 13737 11713 13771 11747
rect 15301 11713 15335 11747
rect 15393 11713 15427 11747
rect 17049 11713 17083 11747
rect 18337 11713 18371 11747
rect 3893 11645 3927 11679
rect 3985 11645 4019 11679
rect 11069 11645 11103 11679
rect 18153 11645 18187 11679
rect 19441 11645 19475 11679
rect 19708 11645 19742 11679
rect 7104 11577 7138 11611
rect 9413 11577 9447 11611
rect 9505 11577 9539 11611
rect 10977 11577 11011 11611
rect 13553 11577 13587 11611
rect 5457 11509 5491 11543
rect 5549 11509 5583 11543
rect 13645 11509 13679 11543
rect 15209 11509 15243 11543
rect 16773 11509 16807 11543
rect 16865 11509 16899 11543
rect 1961 11305 1995 11339
rect 4445 11305 4479 11339
rect 5549 11305 5583 11339
rect 6469 11305 6503 11339
rect 6837 11305 6871 11339
rect 9873 11305 9907 11339
rect 12173 11305 12207 11339
rect 13461 11305 13495 11339
rect 13921 11305 13955 11339
rect 15393 11305 15427 11339
rect 18337 11305 18371 11339
rect 19717 11305 19751 11339
rect 2973 11237 3007 11271
rect 10885 11237 10919 11271
rect 17202 11237 17236 11271
rect 19073 11237 19107 11271
rect 19625 11237 19659 11271
rect 4261 11169 4295 11203
rect 5365 11169 5399 11203
rect 8401 11169 8435 11203
rect 9689 11169 9723 11203
rect 13829 11169 13863 11203
rect 15761 11169 15795 11203
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 8493 11101 8527 11135
rect 8677 11101 8711 11135
rect 14013 11101 14047 11135
rect 15853 11101 15887 11135
rect 15945 11101 15979 11135
rect 16957 11101 16991 11135
rect 19901 11101 19935 11135
rect 8033 11033 8067 11067
rect 19257 11033 19291 11067
rect 9505 10761 9539 10795
rect 9965 10761 9999 10795
rect 13829 10761 13863 10795
rect 16865 10761 16899 10795
rect 17693 10761 17727 10795
rect 18245 10761 18279 10795
rect 5825 10693 5859 10727
rect 12173 10693 12207 10727
rect 3617 10625 3651 10659
rect 10609 10625 10643 10659
rect 19165 10625 19199 10659
rect 2605 10557 2639 10591
rect 5641 10557 5675 10591
rect 6837 10557 6871 10591
rect 8125 10557 8159 10591
rect 10425 10557 10459 10591
rect 10793 10557 10827 10591
rect 12449 10557 12483 10591
rect 15485 10557 15519 10591
rect 15752 10557 15786 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 4537 10489 4571 10523
rect 4629 10489 4663 10523
rect 7113 10489 7147 10523
rect 8392 10489 8426 10523
rect 11060 10489 11094 10523
rect 12694 10489 12728 10523
rect 19432 10489 19466 10523
rect 10333 10421 10367 10455
rect 20545 10421 20579 10455
rect 4721 10217 4755 10251
rect 4813 10217 4847 10251
rect 6009 10217 6043 10251
rect 8033 10217 8067 10251
rect 8493 10217 8527 10251
rect 12173 10217 12207 10251
rect 13921 10217 13955 10251
rect 15568 10149 15602 10183
rect 19165 10149 19199 10183
rect 5825 10081 5859 10115
rect 6929 10081 6963 10115
rect 8401 10081 8435 10115
rect 10232 10081 10266 10115
rect 12541 10081 12575 10115
rect 13737 10081 13771 10115
rect 15025 10081 15059 10115
rect 17509 10081 17543 10115
rect 19257 10081 19291 10115
rect 8677 10013 8711 10047
rect 9965 10013 9999 10047
rect 12633 10013 12667 10047
rect 12725 10013 12759 10047
rect 15301 10013 15335 10047
rect 17693 10013 17727 10047
rect 19349 10013 19383 10047
rect 11345 9945 11379 9979
rect 16681 9945 16715 9979
rect 7113 9877 7147 9911
rect 14841 9877 14875 9911
rect 18797 9877 18831 9911
rect 10517 9673 10551 9707
rect 12633 9605 12667 9639
rect 16865 9605 16899 9639
rect 18521 9605 18555 9639
rect 20821 9605 20855 9639
rect 5733 9537 5767 9571
rect 11345 9537 11379 9571
rect 14197 9537 14231 9571
rect 15761 9537 15795 9571
rect 19441 9537 19475 9571
rect 6929 9469 6963 9503
rect 9137 9469 9171 9503
rect 12449 9469 12483 9503
rect 14013 9469 14047 9503
rect 16681 9469 16715 9503
rect 18337 9469 18371 9503
rect 3617 9401 3651 9435
rect 3709 9401 3743 9435
rect 7196 9401 7230 9435
rect 9404 9401 9438 9435
rect 15485 9401 15519 9435
rect 15577 9401 15611 9435
rect 19708 9401 19742 9435
rect 4721 9333 4755 9367
rect 8309 9333 8343 9367
rect 13553 9333 13587 9367
rect 13921 9333 13955 9367
rect 15117 9333 15151 9367
rect 4629 9129 4663 9163
rect 8033 9129 8067 9163
rect 13645 9129 13679 9163
rect 16405 9129 16439 9163
rect 16865 9129 16899 9163
rect 19349 9129 19383 9163
rect 5641 9061 5675 9095
rect 16773 9061 16807 9095
rect 6653 8993 6687 9027
rect 6920 8993 6954 9027
rect 9045 8993 9079 9027
rect 10701 8993 10735 9027
rect 10968 8993 11002 9027
rect 14013 8993 14047 9027
rect 14105 8993 14139 9027
rect 15301 8993 15335 9027
rect 18225 8993 18259 9027
rect 9689 8925 9723 8959
rect 14197 8925 14231 8959
rect 17049 8925 17083 8959
rect 17969 8925 18003 8959
rect 15485 8857 15519 8891
rect 8861 8789 8895 8823
rect 12081 8789 12115 8823
rect 11437 8585 11471 8619
rect 16405 8585 16439 8619
rect 7941 8517 7975 8551
rect 14197 8517 14231 8551
rect 17233 8517 17267 8551
rect 8493 8449 8527 8483
rect 10057 8449 10091 8483
rect 18613 8449 18647 8483
rect 20545 8449 20579 8483
rect 20637 8449 20671 8483
rect 9873 8381 9907 8415
rect 11253 8381 11287 8415
rect 12817 8381 12851 8415
rect 15025 8381 15059 8415
rect 15281 8381 15315 8415
rect 17417 8381 17451 8415
rect 18429 8381 18463 8415
rect 4721 8313 4755 8347
rect 5733 8313 5767 8347
rect 13062 8313 13096 8347
rect 18521 8313 18555 8347
rect 19901 8313 19935 8347
rect 20453 8313 20487 8347
rect 6929 8245 6963 8279
rect 8309 8245 8343 8279
rect 8401 8245 8435 8279
rect 9505 8245 9539 8279
rect 9965 8245 9999 8279
rect 18061 8245 18095 8279
rect 20085 8245 20119 8279
rect 4445 8041 4479 8075
rect 6837 8041 6871 8075
rect 8033 8041 8067 8075
rect 9229 8041 9263 8075
rect 12449 8041 12483 8075
rect 13553 8041 13587 8075
rect 13921 8041 13955 8075
rect 18797 8041 18831 8075
rect 15945 7973 15979 8007
rect 16037 7973 16071 8007
rect 19165 7973 19199 8007
rect 5457 7905 5491 7939
rect 5724 7905 5758 7939
rect 9413 7905 9447 7939
rect 10048 7905 10082 7939
rect 12357 7905 12391 7939
rect 17601 7905 17635 7939
rect 8125 7837 8159 7871
rect 8217 7837 8251 7871
rect 9781 7837 9815 7871
rect 12541 7837 12575 7871
rect 14013 7837 14047 7871
rect 14105 7837 14139 7871
rect 16129 7837 16163 7871
rect 17693 7837 17727 7871
rect 17785 7837 17819 7871
rect 19257 7837 19291 7871
rect 19349 7837 19383 7871
rect 7665 7769 7699 7803
rect 11161 7701 11195 7735
rect 11989 7701 12023 7735
rect 15577 7701 15611 7735
rect 17233 7701 17267 7735
rect 6469 7497 6503 7531
rect 10701 7497 10735 7531
rect 12449 7497 12483 7531
rect 19441 7497 19475 7531
rect 9873 7429 9907 7463
rect 7021 7361 7055 7395
rect 11253 7361 11287 7395
rect 13093 7361 13127 7395
rect 14473 7361 14507 7395
rect 14657 7361 14691 7395
rect 16037 7361 16071 7395
rect 16221 7361 16255 7395
rect 18061 7361 18095 7395
rect 2973 7293 3007 7327
rect 5181 7293 5215 7327
rect 5457 7293 5491 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 8493 7293 8527 7327
rect 12817 7293 12851 7327
rect 14381 7293 14415 7327
rect 15945 7293 15979 7327
rect 20545 7293 20579 7327
rect 3218 7225 3252 7259
rect 8760 7225 8794 7259
rect 11069 7225 11103 7259
rect 18328 7225 18362 7259
rect 4353 7157 4387 7191
rect 11161 7157 11195 7191
rect 12909 7157 12943 7191
rect 14013 7157 14047 7191
rect 15577 7157 15611 7191
rect 20729 7157 20763 7191
rect 6009 6953 6043 6987
rect 7757 6953 7791 6987
rect 10885 6953 10919 6987
rect 12081 6953 12115 6987
rect 14105 6953 14139 6987
rect 8125 6885 8159 6919
rect 12449 6885 12483 6919
rect 14013 6885 14047 6919
rect 15568 6885 15602 6919
rect 4997 6817 5031 6851
rect 6377 6817 6411 6851
rect 15301 6817 15335 6851
rect 17693 6817 17727 6851
rect 17960 6817 17994 6851
rect 6469 6749 6503 6783
rect 6653 6749 6687 6783
rect 8217 6749 8251 6783
rect 8401 6749 8435 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 12541 6749 12575 6783
rect 12633 6749 12667 6783
rect 14289 6749 14323 6783
rect 10517 6681 10551 6715
rect 13645 6681 13679 6715
rect 16681 6613 16715 6647
rect 19073 6613 19107 6647
rect 3801 6409 3835 6443
rect 16589 6409 16623 6443
rect 10701 6341 10735 6375
rect 4353 6273 4387 6307
rect 6837 6273 6871 6307
rect 9321 6273 9355 6307
rect 12909 6273 12943 6307
rect 13001 6273 13035 6307
rect 15209 6273 15243 6307
rect 18613 6273 18647 6307
rect 18797 6273 18831 6307
rect 20361 6273 20395 6307
rect 2789 6205 2823 6239
rect 9588 6205 9622 6239
rect 14105 6205 14139 6239
rect 15476 6205 15510 6239
rect 18521 6205 18555 6239
rect 7104 6137 7138 6171
rect 20177 6137 20211 6171
rect 4169 6069 4203 6103
rect 4261 6069 4295 6103
rect 5733 6069 5767 6103
rect 8217 6069 8251 6103
rect 12449 6069 12483 6103
rect 12817 6069 12851 6103
rect 14289 6069 14323 6103
rect 18153 6069 18187 6103
rect 19717 6069 19751 6103
rect 20085 6069 20119 6103
rect 2973 5865 3007 5899
rect 7665 5865 7699 5899
rect 8677 5865 8711 5899
rect 12265 5865 12299 5899
rect 12357 5865 12391 5899
rect 13461 5865 13495 5899
rect 13829 5865 13863 5899
rect 19257 5865 19291 5899
rect 1869 5797 1903 5831
rect 1961 5797 1995 5831
rect 6530 5797 6564 5831
rect 17040 5797 17074 5831
rect 19625 5797 19659 5831
rect 4344 5729 4378 5763
rect 8493 5729 8527 5763
rect 9689 5729 9723 5763
rect 9956 5729 9990 5763
rect 15669 5729 15703 5763
rect 4077 5661 4111 5695
rect 6285 5661 6319 5695
rect 12449 5661 12483 5695
rect 13921 5661 13955 5695
rect 14105 5661 14139 5695
rect 16773 5661 16807 5695
rect 19717 5661 19751 5695
rect 19901 5661 19935 5695
rect 5457 5593 5491 5627
rect 11069 5525 11103 5559
rect 11897 5525 11931 5559
rect 15853 5525 15887 5559
rect 18153 5525 18187 5559
rect 4537 5321 4571 5355
rect 8769 5321 8803 5355
rect 20821 5321 20855 5355
rect 12817 5253 12851 5287
rect 17049 5253 17083 5287
rect 3157 5185 3191 5219
rect 7389 5185 7423 5219
rect 11345 5185 11379 5219
rect 14197 5185 14231 5219
rect 14289 5185 14323 5219
rect 15853 5185 15887 5219
rect 19441 5185 19475 5219
rect 5641 5117 5675 5151
rect 7656 5117 7690 5151
rect 9689 5117 9723 5151
rect 11161 5117 11195 5151
rect 11253 5117 11287 5151
rect 12633 5117 12667 5151
rect 15669 5117 15703 5151
rect 16865 5117 16899 5151
rect 18337 5117 18371 5151
rect 3424 5049 3458 5083
rect 19708 5049 19742 5083
rect 2145 4981 2179 5015
rect 5825 4981 5859 5015
rect 9873 4981 9907 5015
rect 10793 4981 10827 5015
rect 13737 4981 13771 5015
rect 14105 4981 14139 5015
rect 15301 4981 15335 5015
rect 15761 4981 15795 5015
rect 18521 4981 18555 5015
rect 2421 4777 2455 4811
rect 4905 4777 4939 4811
rect 6469 4777 6503 4811
rect 8493 4777 8527 4811
rect 12265 4777 12299 4811
rect 14105 4777 14139 4811
rect 15301 4777 15335 4811
rect 15761 4777 15795 4811
rect 17325 4777 17359 4811
rect 6929 4709 6963 4743
rect 8401 4709 8435 4743
rect 11130 4709 11164 4743
rect 14013 4709 14047 4743
rect 17417 4709 17451 4743
rect 18766 4709 18800 4743
rect 2789 4641 2823 4675
rect 5273 4641 5307 4675
rect 6837 4641 6871 4675
rect 9781 4641 9815 4675
rect 15669 4641 15703 4675
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 7113 4573 7147 4607
rect 8677 4573 8711 4607
rect 10885 4573 10919 4607
rect 14289 4573 14323 4607
rect 15853 4573 15887 4607
rect 17601 4573 17635 4607
rect 18521 4573 18555 4607
rect 8033 4505 8067 4539
rect 9965 4437 9999 4471
rect 13645 4437 13679 4471
rect 16957 4437 16991 4471
rect 19901 4437 19935 4471
rect 4169 4233 4203 4267
rect 7021 4165 7055 4199
rect 13829 4165 13863 4199
rect 2789 4097 2823 4131
rect 5733 4097 5767 4131
rect 7573 4097 7607 4131
rect 15209 4097 15243 4131
rect 17049 4097 17083 4131
rect 3056 4029 3090 4063
rect 7481 4029 7515 4063
rect 8585 4029 8619 4063
rect 8852 4029 8886 4063
rect 10793 4029 10827 4063
rect 12449 4029 12483 4063
rect 12705 4029 12739 4063
rect 15025 4029 15059 4063
rect 18337 4029 18371 4063
rect 19441 4029 19475 4063
rect 19697 4029 19731 4063
rect 5549 3961 5583 3995
rect 11069 3961 11103 3995
rect 15117 3961 15151 3995
rect 1777 3893 1811 3927
rect 5181 3893 5215 3927
rect 5641 3893 5675 3927
rect 7389 3893 7423 3927
rect 9965 3893 9999 3927
rect 14657 3893 14691 3927
rect 16405 3893 16439 3927
rect 16773 3893 16807 3927
rect 16865 3893 16899 3927
rect 18521 3893 18555 3927
rect 20821 3893 20855 3927
rect 5825 3689 5859 3723
rect 11069 3689 11103 3723
rect 14013 3689 14047 3723
rect 14105 3689 14139 3723
rect 17969 3689 18003 3723
rect 18429 3689 18463 3723
rect 17785 3621 17819 3655
rect 18337 3621 18371 3655
rect 1777 3553 1811 3587
rect 2881 3553 2915 3587
rect 4712 3553 4746 3587
rect 6745 3553 6779 3587
rect 7012 3553 7046 3587
rect 9956 3553 9990 3587
rect 11897 3553 11931 3587
rect 16017 3553 16051 3587
rect 19533 3553 19567 3587
rect 4445 3485 4479 3519
rect 9689 3485 9723 3519
rect 12081 3485 12115 3519
rect 14289 3485 14323 3519
rect 15761 3485 15795 3519
rect 18613 3485 18647 3519
rect 19717 3485 19751 3519
rect 17141 3417 17175 3451
rect 1961 3349 1995 3383
rect 3065 3349 3099 3383
rect 8125 3349 8159 3383
rect 13645 3349 13679 3383
rect 5457 3145 5491 3179
rect 8217 3145 8251 3179
rect 9689 3145 9723 3179
rect 11437 3145 11471 3179
rect 15761 3145 15795 3179
rect 18061 3145 18095 3179
rect 2053 3077 2087 3111
rect 3157 3077 3191 3111
rect 6837 3009 6871 3043
rect 10241 3009 10275 3043
rect 14381 3009 14415 3043
rect 16865 3009 16899 3043
rect 18613 3009 18647 3043
rect 20177 3009 20211 3043
rect 1869 2941 1903 2975
rect 2973 2941 3007 2975
rect 4077 2941 4111 2975
rect 11253 2941 11287 2975
rect 12725 2941 12759 2975
rect 16681 2941 16715 2975
rect 18521 2941 18555 2975
rect 19993 2941 20027 2975
rect 4344 2873 4378 2907
rect 7104 2873 7138 2907
rect 13001 2873 13035 2907
rect 14648 2873 14682 2907
rect 18429 2873 18463 2907
rect 10057 2805 10091 2839
rect 10149 2805 10183 2839
rect 19625 2805 19659 2839
rect 20085 2805 20119 2839
rect 4905 2601 4939 2635
rect 7205 2601 7239 2635
rect 7665 2601 7699 2635
rect 9781 2601 9815 2635
rect 11621 2601 11655 2635
rect 14197 2533 14231 2567
rect 2881 2465 2915 2499
rect 5273 2465 5307 2499
rect 7573 2465 7607 2499
rect 10149 2465 10183 2499
rect 10241 2465 10275 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 13921 2465 13955 2499
rect 16037 2465 16071 2499
rect 17141 2465 17175 2499
rect 18981 2465 19015 2499
rect 1869 2397 1903 2431
rect 5365 2397 5399 2431
rect 5457 2397 5491 2431
rect 7757 2397 7791 2431
rect 10333 2397 10367 2431
rect 12817 2397 12851 2431
rect 19165 2397 19199 2431
rect 16221 2329 16255 2363
rect 3065 2261 3099 2295
rect 17325 2261 17359 2295
<< metal1 >>
rect 10226 21088 10232 21140
rect 10284 21128 10290 21140
rect 18322 21128 18328 21140
rect 10284 21100 18328 21128
rect 10284 21088 10290 21100
rect 18322 21088 18328 21100
rect 18380 21088 18386 21140
rect 3142 20952 3148 21004
rect 3200 20992 3206 21004
rect 18690 20992 18696 21004
rect 3200 20964 18696 20992
rect 3200 20952 3206 20964
rect 18690 20952 18696 20964
rect 18748 20952 18754 21004
rect 2866 20884 2872 20936
rect 2924 20924 2930 20936
rect 17954 20924 17960 20936
rect 2924 20896 17960 20924
rect 2924 20884 2930 20896
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 2222 20816 2228 20868
rect 2280 20856 2286 20868
rect 18046 20856 18052 20868
rect 2280 20828 18052 20856
rect 2280 20816 2286 20828
rect 18046 20816 18052 20828
rect 18104 20816 18110 20868
rect 1946 20748 1952 20800
rect 2004 20788 2010 20800
rect 18138 20788 18144 20800
rect 2004 20760 18144 20788
rect 2004 20748 2010 20760
rect 18138 20748 18144 20760
rect 18196 20748 18202 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 1946 20584 1952 20596
rect 1907 20556 1952 20584
rect 1946 20544 1952 20556
rect 2004 20544 2010 20596
rect 3053 20587 3111 20593
rect 3053 20553 3065 20587
rect 3099 20584 3111 20587
rect 3142 20584 3148 20596
rect 3099 20556 3148 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 18138 20584 18144 20596
rect 3292 20556 18144 20584
rect 3292 20544 3298 20556
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 4617 20519 4675 20525
rect 4617 20485 4629 20519
rect 4663 20516 4675 20519
rect 5442 20516 5448 20528
rect 4663 20488 5448 20516
rect 4663 20485 4675 20488
rect 4617 20479 4675 20485
rect 5442 20476 5448 20488
rect 5500 20476 5506 20528
rect 6914 20516 6920 20528
rect 6875 20488 6920 20516
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 7558 20476 7564 20528
rect 7616 20516 7622 20528
rect 11054 20516 11060 20528
rect 7616 20488 11060 20516
rect 7616 20476 7622 20488
rect 11054 20476 11060 20488
rect 11112 20476 11118 20528
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 13817 20519 13875 20525
rect 13817 20516 13829 20519
rect 11204 20488 13829 20516
rect 11204 20476 11210 20488
rect 13817 20485 13829 20488
rect 13863 20485 13875 20519
rect 20346 20516 20352 20528
rect 13817 20479 13875 20485
rect 13924 20488 20352 20516
rect 1780 20420 4752 20448
rect 1780 20389 1808 20420
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20349 1823 20383
rect 1765 20343 1823 20349
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 3142 20380 3148 20392
rect 2915 20352 3148 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 3142 20340 3148 20352
rect 3200 20340 3206 20392
rect 4724 20380 4752 20420
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4856 20420 5089 20448
rect 4856 20408 4862 20420
rect 5077 20417 5089 20420
rect 5123 20417 5135 20451
rect 5077 20411 5135 20417
rect 5166 20408 5172 20460
rect 5224 20448 5230 20460
rect 5224 20420 5269 20448
rect 5224 20408 5230 20420
rect 6822 20408 6828 20460
rect 6880 20448 6886 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 6880 20420 7481 20448
rect 6880 20408 6886 20420
rect 7469 20417 7481 20420
rect 7515 20417 7527 20451
rect 7469 20411 7527 20417
rect 8478 20408 8484 20460
rect 8536 20448 8542 20460
rect 11241 20451 11299 20457
rect 11241 20448 11253 20451
rect 8536 20420 11253 20448
rect 8536 20408 8542 20420
rect 11241 20417 11253 20420
rect 11287 20417 11299 20451
rect 11241 20411 11299 20417
rect 5718 20380 5724 20392
rect 4724 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 6178 20340 6184 20392
rect 6236 20380 6242 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 6236 20352 7389 20380
rect 6236 20340 6242 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 8570 20380 8576 20392
rect 8531 20352 8576 20380
rect 7377 20343 7435 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 9769 20383 9827 20389
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 10318 20380 10324 20392
rect 9815 20352 10324 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 10318 20340 10324 20352
rect 10376 20340 10382 20392
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20349 11115 20383
rect 11057 20343 11115 20349
rect 12713 20383 12771 20389
rect 12713 20349 12725 20383
rect 12759 20380 12771 20383
rect 13924 20380 13952 20488
rect 20346 20476 20352 20488
rect 20404 20476 20410 20528
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20448 14519 20451
rect 14734 20448 14740 20460
rect 14507 20420 14740 20448
rect 14507 20417 14519 20420
rect 14461 20411 14519 20417
rect 14734 20408 14740 20420
rect 14792 20448 14798 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 14792 20420 16037 20448
rect 14792 20408 14798 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 16025 20411 16083 20417
rect 17144 20420 18521 20448
rect 12759 20352 13952 20380
rect 14200 20380 14228 20408
rect 17144 20389 17172 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 19889 20451 19947 20457
rect 19889 20448 19901 20451
rect 19668 20420 19901 20448
rect 19668 20408 19674 20420
rect 19889 20417 19901 20420
rect 19935 20417 19947 20451
rect 19889 20411 19947 20417
rect 17129 20383 17187 20389
rect 14200 20352 15516 20380
rect 12759 20349 12771 20352
rect 12713 20343 12771 20349
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 7285 20315 7343 20321
rect 7285 20312 7297 20315
rect 6788 20284 7297 20312
rect 6788 20272 6794 20284
rect 7285 20281 7297 20284
rect 7331 20281 7343 20315
rect 9858 20312 9864 20324
rect 7285 20275 7343 20281
rect 7392 20284 9864 20312
rect 2498 20204 2504 20256
rect 2556 20244 2562 20256
rect 2866 20244 2872 20256
rect 2556 20216 2872 20244
rect 2556 20204 2562 20216
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 4985 20247 5043 20253
rect 4985 20213 4997 20247
rect 5031 20244 5043 20247
rect 5074 20244 5080 20256
rect 5031 20216 5080 20244
rect 5031 20213 5043 20216
rect 4985 20207 5043 20213
rect 5074 20204 5080 20216
rect 5132 20244 5138 20256
rect 5258 20244 5264 20256
rect 5132 20216 5264 20244
rect 5132 20204 5138 20216
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 6362 20204 6368 20256
rect 6420 20244 6426 20256
rect 7392 20244 7420 20284
rect 9858 20272 9864 20284
rect 9916 20272 9922 20324
rect 10045 20315 10103 20321
rect 10045 20281 10057 20315
rect 10091 20312 10103 20315
rect 10134 20312 10140 20324
rect 10091 20284 10140 20312
rect 10091 20281 10103 20284
rect 10045 20275 10103 20281
rect 10134 20272 10140 20284
rect 10192 20272 10198 20324
rect 6420 20216 7420 20244
rect 8757 20247 8815 20253
rect 6420 20204 6426 20216
rect 8757 20213 8769 20247
rect 8803 20244 8815 20247
rect 10594 20244 10600 20256
rect 8803 20216 10600 20244
rect 8803 20213 8815 20216
rect 8757 20207 8815 20213
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 11082 20244 11110 20343
rect 11790 20272 11796 20324
rect 11848 20312 11854 20324
rect 13998 20312 14004 20324
rect 11848 20284 14004 20312
rect 11848 20272 11854 20284
rect 13998 20272 14004 20284
rect 14056 20272 14062 20324
rect 14185 20315 14243 20321
rect 14185 20281 14197 20315
rect 14231 20312 14243 20315
rect 14366 20312 14372 20324
rect 14231 20284 14372 20312
rect 14231 20281 14243 20284
rect 14185 20275 14243 20281
rect 14366 20272 14372 20284
rect 14424 20272 14430 20324
rect 12250 20244 12256 20256
rect 11082 20216 12256 20244
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 12897 20247 12955 20253
rect 12897 20213 12909 20247
rect 12943 20244 12955 20247
rect 13262 20244 13268 20256
rect 12943 20216 13268 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15488 20253 15516 20352
rect 17129 20349 17141 20383
rect 17175 20349 17187 20383
rect 17129 20343 17187 20349
rect 17218 20340 17224 20392
rect 17276 20380 17282 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 17276 20352 18337 20380
rect 17276 20340 17282 20352
rect 18325 20349 18337 20352
rect 18371 20349 18383 20383
rect 19702 20380 19708 20392
rect 19663 20352 19708 20380
rect 18325 20343 18383 20349
rect 19702 20340 19708 20352
rect 19760 20340 19766 20392
rect 15562 20272 15568 20324
rect 15620 20312 15626 20324
rect 15620 20284 15976 20312
rect 15620 20272 15626 20284
rect 14277 20247 14335 20253
rect 14277 20244 14289 20247
rect 13872 20216 14289 20244
rect 13872 20204 13878 20216
rect 14277 20213 14289 20216
rect 14323 20213 14335 20247
rect 14277 20207 14335 20213
rect 15473 20247 15531 20253
rect 15473 20213 15485 20247
rect 15519 20213 15531 20247
rect 15473 20207 15531 20213
rect 15654 20204 15660 20256
rect 15712 20244 15718 20256
rect 15948 20253 15976 20284
rect 15841 20247 15899 20253
rect 15841 20244 15853 20247
rect 15712 20216 15853 20244
rect 15712 20204 15718 20216
rect 15841 20213 15853 20216
rect 15887 20213 15899 20247
rect 15841 20207 15899 20213
rect 15933 20247 15991 20253
rect 15933 20213 15945 20247
rect 15979 20244 15991 20247
rect 16206 20244 16212 20256
rect 15979 20216 16212 20244
rect 15979 20213 15991 20216
rect 15933 20207 15991 20213
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 17313 20247 17371 20253
rect 17313 20213 17325 20247
rect 17359 20244 17371 20247
rect 17770 20244 17776 20256
rect 17359 20216 17776 20244
rect 17359 20213 17371 20216
rect 17313 20207 17371 20213
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2222 20040 2228 20052
rect 1995 20012 2228 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2222 20000 2228 20012
rect 2280 20000 2286 20052
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 6825 20043 6883 20049
rect 3099 20012 6408 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 4516 19975 4574 19981
rect 4516 19941 4528 19975
rect 4562 19972 4574 19975
rect 4798 19972 4804 19984
rect 4562 19944 4804 19972
rect 4562 19941 4574 19944
rect 4516 19935 4574 19941
rect 4798 19932 4804 19944
rect 4856 19972 4862 19984
rect 5166 19972 5172 19984
rect 4856 19944 5172 19972
rect 4856 19932 4862 19944
rect 5166 19932 5172 19944
rect 5224 19932 5230 19984
rect 6380 19972 6408 20012
rect 6825 20009 6837 20043
rect 6871 20040 6883 20043
rect 9674 20040 9680 20052
rect 6871 20012 9680 20040
rect 6871 20009 6883 20012
rect 6825 20003 6883 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 11698 20000 11704 20052
rect 11756 20040 11762 20052
rect 13173 20043 13231 20049
rect 13173 20040 13185 20043
rect 11756 20012 13185 20040
rect 11756 20000 11762 20012
rect 13173 20009 13185 20012
rect 13219 20009 13231 20043
rect 13173 20003 13231 20009
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 17862 20040 17868 20052
rect 13320 20012 17868 20040
rect 13320 20000 13326 20012
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 9766 19972 9772 19984
rect 6380 19944 9772 19972
rect 9766 19932 9772 19944
rect 9824 19932 9830 19984
rect 9950 19981 9956 19984
rect 9944 19935 9956 19981
rect 10008 19972 10014 19984
rect 10008 19944 10044 19972
rect 9950 19932 9956 19935
rect 10008 19932 10014 19944
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 1765 19867 1823 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 6638 19904 6644 19916
rect 2915 19876 6644 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 1780 19700 1808 19867
rect 6638 19864 6644 19876
rect 6696 19864 6702 19916
rect 6822 19864 6828 19916
rect 6880 19904 6886 19916
rect 7173 19907 7231 19913
rect 7173 19904 7185 19907
rect 6880 19876 7185 19904
rect 6880 19864 6886 19876
rect 7173 19873 7185 19876
rect 7219 19873 7231 19907
rect 7173 19867 7231 19873
rect 7466 19864 7472 19916
rect 7524 19904 7530 19916
rect 13354 19904 13360 19916
rect 7524 19876 13360 19904
rect 7524 19864 7530 19876
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 4246 19836 4252 19848
rect 4207 19808 4252 19836
rect 4246 19796 4252 19808
rect 4304 19796 4310 19848
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 6825 19771 6883 19777
rect 6825 19768 6837 19771
rect 5552 19740 6837 19768
rect 5552 19700 5580 19740
rect 6825 19737 6837 19740
rect 6871 19737 6883 19771
rect 6825 19731 6883 19737
rect 1780 19672 5580 19700
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 6932 19700 6960 19799
rect 9674 19796 9680 19848
rect 9732 19845 9738 19848
rect 9732 19836 9742 19845
rect 9732 19808 9777 19836
rect 9732 19799 9742 19808
rect 9732 19796 9738 19799
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 11882 19836 11888 19848
rect 11112 19808 11888 19836
rect 11112 19796 11118 19808
rect 11882 19796 11888 19808
rect 11940 19836 11946 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 11940 19808 13277 19836
rect 11940 19796 11946 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13446 19836 13452 19848
rect 13407 19808 13452 19836
rect 13265 19799 13323 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 13630 19796 13636 19848
rect 13688 19836 13694 19848
rect 15672 19836 15700 19867
rect 16022 19864 16028 19916
rect 16080 19904 16086 19916
rect 16853 19907 16911 19913
rect 16853 19904 16865 19907
rect 16080 19876 16865 19904
rect 16080 19864 16086 19876
rect 16853 19873 16865 19876
rect 16899 19873 16911 19907
rect 16853 19867 16911 19873
rect 18046 19864 18052 19916
rect 18104 19904 18110 19916
rect 18141 19907 18199 19913
rect 18141 19904 18153 19907
rect 18104 19876 18153 19904
rect 18104 19864 18110 19876
rect 18141 19873 18153 19876
rect 18187 19873 18199 19907
rect 19518 19904 19524 19916
rect 19479 19876 19524 19904
rect 18141 19867 18199 19873
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 13688 19808 15700 19836
rect 15749 19839 15807 19845
rect 13688 19796 13694 19808
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15749 19799 15807 19805
rect 15856 19808 15945 19836
rect 8018 19728 8024 19780
rect 8076 19768 8082 19780
rect 15764 19768 15792 19799
rect 15856 19780 15884 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 16172 19808 17049 19836
rect 16172 19796 16178 19808
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17126 19796 17132 19848
rect 17184 19836 17190 19848
rect 18325 19839 18383 19845
rect 18325 19836 18337 19839
rect 17184 19808 18337 19836
rect 17184 19796 17190 19808
rect 18325 19805 18337 19808
rect 18371 19805 18383 19839
rect 18325 19799 18383 19805
rect 19705 19839 19763 19845
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 8076 19740 8524 19768
rect 8076 19728 8082 19740
rect 8110 19700 8116 19712
rect 5684 19672 5729 19700
rect 6932 19672 8116 19700
rect 5684 19660 5690 19672
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 8386 19700 8392 19712
rect 8343 19672 8392 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 8496 19700 8524 19740
rect 10888 19740 15792 19768
rect 10888 19700 10916 19740
rect 15838 19728 15844 19780
rect 15896 19728 15902 19780
rect 17310 19728 17316 19780
rect 17368 19768 17374 19780
rect 19720 19768 19748 19799
rect 17368 19740 19748 19768
rect 17368 19728 17374 19740
rect 8496 19672 10916 19700
rect 10962 19660 10968 19712
rect 11020 19700 11026 19712
rect 11057 19703 11115 19709
rect 11057 19700 11069 19703
rect 11020 19672 11069 19700
rect 11020 19660 11026 19672
rect 11057 19669 11069 19672
rect 11103 19669 11115 19703
rect 11057 19663 11115 19669
rect 12805 19703 12863 19709
rect 12805 19669 12817 19703
rect 12851 19700 12863 19703
rect 14182 19700 14188 19712
rect 12851 19672 14188 19700
rect 12851 19669 12863 19672
rect 12805 19663 12863 19669
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 1452 19468 9076 19496
rect 1452 19456 1458 19468
rect 4798 19428 4804 19440
rect 4759 19400 4804 19428
rect 4798 19388 4804 19400
rect 4856 19388 4862 19440
rect 7558 19388 7564 19440
rect 7616 19428 7622 19440
rect 8018 19428 8024 19440
rect 7616 19400 8024 19428
rect 7616 19388 7622 19400
rect 8018 19388 8024 19400
rect 8076 19388 8082 19440
rect 9048 19428 9076 19468
rect 9950 19456 9956 19508
rect 10008 19496 10014 19508
rect 10134 19496 10140 19508
rect 10008 19468 10140 19496
rect 10008 19456 10014 19468
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 10594 19456 10600 19508
rect 10652 19496 10658 19508
rect 13078 19496 13084 19508
rect 10652 19468 13084 19496
rect 10652 19456 10658 19468
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 17126 19496 17132 19508
rect 13188 19468 17132 19496
rect 13188 19428 13216 19468
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19576 19468 19625 19496
rect 19576 19456 19582 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 9048 19400 13216 19428
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 7466 19360 7472 19372
rect 3384 19332 3556 19360
rect 3384 19320 3390 19332
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2406 19292 2412 19304
rect 2363 19264 2412 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2406 19252 2412 19264
rect 2464 19252 2470 19304
rect 2590 19252 2596 19304
rect 2648 19292 2654 19304
rect 3421 19295 3479 19301
rect 3421 19292 3433 19295
rect 2648 19264 3433 19292
rect 2648 19252 2654 19264
rect 3421 19261 3433 19264
rect 3467 19261 3479 19295
rect 3528 19292 3556 19332
rect 4448 19332 7472 19360
rect 4448 19292 4476 19332
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 9674 19360 9680 19372
rect 9140 19332 9680 19360
rect 3528 19264 4476 19292
rect 5629 19295 5687 19301
rect 3421 19255 3479 19261
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 5902 19292 5908 19304
rect 5675 19264 5908 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 842 19184 848 19236
rect 900 19224 906 19236
rect 2866 19224 2872 19236
rect 900 19196 2872 19224
rect 900 19184 906 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 2498 19156 2504 19168
rect 2459 19128 2504 19156
rect 2498 19116 2504 19128
rect 2556 19116 2562 19168
rect 3436 19156 3464 19255
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6086 19252 6092 19304
rect 6144 19292 6150 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6144 19264 6837 19292
rect 6144 19252 6150 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 8110 19292 8116 19304
rect 8023 19264 8116 19292
rect 6825 19255 6883 19261
rect 8110 19252 8116 19264
rect 8168 19252 8174 19304
rect 8386 19301 8392 19304
rect 8380 19292 8392 19301
rect 8347 19264 8392 19292
rect 8380 19255 8392 19264
rect 8444 19292 8450 19304
rect 8662 19292 8668 19304
rect 8444 19264 8668 19292
rect 8386 19252 8392 19255
rect 8444 19252 8450 19264
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 3688 19227 3746 19233
rect 3688 19193 3700 19227
rect 3734 19224 3746 19227
rect 4154 19224 4160 19236
rect 3734 19196 4160 19224
rect 3734 19193 3746 19196
rect 3688 19187 3746 19193
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 6638 19184 6644 19236
rect 6696 19224 6702 19236
rect 7101 19227 7159 19233
rect 7101 19224 7113 19227
rect 6696 19196 7113 19224
rect 6696 19184 6702 19196
rect 7101 19193 7113 19196
rect 7147 19193 7159 19227
rect 8128 19224 8156 19252
rect 8294 19224 8300 19236
rect 8128 19196 8300 19224
rect 7101 19187 7159 19193
rect 8294 19184 8300 19196
rect 8352 19224 8358 19236
rect 9140 19224 9168 19332
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10962 19360 10968 19372
rect 10468 19332 10824 19360
rect 10923 19332 10968 19360
rect 10468 19320 10474 19332
rect 9214 19252 9220 19304
rect 9272 19292 9278 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 9272 19264 10701 19292
rect 9272 19252 9278 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10796 19292 10824 19332
rect 10962 19320 10968 19332
rect 11020 19320 11026 19372
rect 20162 19360 20168 19372
rect 20123 19332 20168 19360
rect 20162 19320 20168 19332
rect 20220 19320 20226 19372
rect 12618 19292 12624 19304
rect 10796 19264 12624 19292
rect 10689 19255 10747 19261
rect 12618 19252 12624 19264
rect 12676 19252 12682 19304
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13173 19295 13231 19301
rect 13173 19292 13185 19295
rect 12952 19264 13185 19292
rect 12952 19252 12958 19264
rect 13173 19261 13185 19264
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 13262 19252 13268 19304
rect 13320 19292 13326 19304
rect 15102 19292 15108 19304
rect 13320 19264 15108 19292
rect 13320 19252 13326 19264
rect 15102 19252 15108 19264
rect 15160 19252 15166 19304
rect 15381 19295 15439 19301
rect 15381 19261 15393 19295
rect 15427 19292 15439 19295
rect 16114 19292 16120 19304
rect 15427 19264 16120 19292
rect 15427 19261 15439 19264
rect 15381 19255 15439 19261
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16942 19252 16948 19304
rect 17000 19292 17006 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17000 19264 18061 19292
rect 17000 19252 17006 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 13446 19233 13452 19236
rect 8352 19196 9168 19224
rect 10781 19227 10839 19233
rect 8352 19184 8358 19196
rect 10781 19193 10793 19227
rect 10827 19224 10839 19227
rect 13440 19224 13452 19233
rect 10827 19196 10916 19224
rect 13407 19196 13452 19224
rect 10827 19193 10839 19196
rect 10781 19187 10839 19193
rect 10888 19168 10916 19196
rect 13440 19187 13452 19196
rect 13446 19184 13452 19187
rect 13504 19184 13510 19236
rect 15626 19227 15684 19233
rect 15626 19224 15638 19227
rect 14568 19196 15638 19224
rect 4338 19156 4344 19168
rect 3436 19128 4344 19156
rect 4338 19116 4344 19128
rect 4396 19156 4402 19168
rect 5534 19156 5540 19168
rect 4396 19128 5540 19156
rect 4396 19116 4402 19128
rect 5534 19116 5540 19128
rect 5592 19116 5598 19168
rect 5810 19156 5816 19168
rect 5771 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 9306 19156 9312 19168
rect 6512 19128 9312 19156
rect 6512 19116 6518 19128
rect 9306 19116 9312 19128
rect 9364 19116 9370 19168
rect 9490 19156 9496 19168
rect 9451 19128 9496 19156
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10318 19156 10324 19168
rect 10279 19128 10324 19156
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10870 19116 10876 19168
rect 10928 19116 10934 19168
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 14568 19165 14596 19196
rect 15626 19193 15638 19196
rect 15672 19224 15684 19227
rect 15838 19224 15844 19236
rect 15672 19196 15844 19224
rect 15672 19193 15684 19196
rect 15626 19187 15684 19193
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 17126 19184 17132 19236
rect 17184 19224 17190 19236
rect 18325 19227 18383 19233
rect 18325 19224 18337 19227
rect 17184 19196 18337 19224
rect 17184 19184 17190 19196
rect 18325 19193 18337 19196
rect 18371 19193 18383 19227
rect 19978 19224 19984 19236
rect 19939 19196 19984 19224
rect 18325 19187 18383 19193
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 14553 19159 14611 19165
rect 14553 19156 14565 19159
rect 14424 19128 14565 19156
rect 14424 19116 14430 19128
rect 14553 19125 14565 19128
rect 14599 19125 14611 19159
rect 16758 19156 16764 19168
rect 16719 19128 16764 19156
rect 14553 19119 14611 19125
rect 16758 19116 16764 19128
rect 16816 19116 16822 19168
rect 20070 19156 20076 19168
rect 20031 19128 20076 19156
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 3053 18955 3111 18961
rect 3053 18921 3065 18955
rect 3099 18952 3111 18955
rect 3234 18952 3240 18964
rect 3099 18924 3240 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 5810 18912 5816 18964
rect 5868 18952 5874 18964
rect 13262 18952 13268 18964
rect 5868 18924 13268 18952
rect 5868 18912 5874 18924
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13504 18924 13921 18952
rect 13504 18912 13510 18924
rect 13909 18921 13921 18924
rect 13955 18921 13967 18955
rect 13909 18915 13967 18921
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 17218 18952 17224 18964
rect 15528 18924 17224 18952
rect 15528 18912 15534 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 5166 18884 5172 18896
rect 4172 18856 5172 18884
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 2590 18816 2596 18828
rect 1811 18788 2596 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18816 2927 18819
rect 4062 18816 4068 18828
rect 2915 18788 4068 18816
rect 2915 18785 2927 18788
rect 2869 18779 2927 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4172 18825 4200 18856
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 5626 18844 5632 18896
rect 5684 18893 5690 18896
rect 5684 18887 5748 18893
rect 5684 18853 5702 18887
rect 5736 18853 5748 18887
rect 5684 18847 5748 18853
rect 5684 18844 5690 18847
rect 5994 18844 6000 18896
rect 6052 18884 6058 18896
rect 6638 18884 6644 18896
rect 6052 18856 6644 18884
rect 6052 18844 6058 18856
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 7006 18844 7012 18896
rect 7064 18884 7070 18896
rect 8389 18887 8447 18893
rect 8389 18884 8401 18887
rect 7064 18856 8401 18884
rect 7064 18844 7070 18856
rect 8389 18853 8401 18856
rect 8435 18853 8447 18887
rect 10410 18884 10416 18896
rect 8389 18847 8447 18853
rect 8496 18856 10416 18884
rect 4157 18819 4215 18825
rect 4157 18785 4169 18819
rect 4203 18785 4215 18819
rect 4157 18779 4215 18785
rect 5534 18776 5540 18828
rect 5592 18776 5598 18828
rect 8496 18816 8524 18856
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 10588 18887 10646 18893
rect 10588 18853 10600 18887
rect 10634 18884 10646 18887
rect 10962 18884 10968 18896
rect 10634 18856 10968 18884
rect 10634 18853 10646 18856
rect 10588 18847 10646 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 11054 18844 11060 18896
rect 11112 18884 11118 18896
rect 11974 18884 11980 18896
rect 11112 18856 11980 18884
rect 11112 18844 11118 18856
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 12066 18844 12072 18896
rect 12124 18884 12130 18896
rect 15289 18887 15347 18893
rect 15289 18884 15301 18887
rect 12124 18856 15301 18884
rect 12124 18844 12130 18856
rect 15289 18853 15301 18856
rect 15335 18853 15347 18887
rect 15289 18847 15347 18853
rect 16568 18887 16626 18893
rect 16568 18853 16580 18887
rect 16614 18884 16626 18887
rect 16758 18884 16764 18896
rect 16614 18856 16764 18884
rect 16614 18853 16626 18856
rect 16568 18847 16626 18853
rect 16758 18844 16764 18856
rect 16816 18844 16822 18896
rect 20990 18884 20996 18896
rect 18064 18856 20996 18884
rect 8662 18816 8668 18828
rect 8220 18788 8524 18816
rect 8588 18788 8668 18816
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 5350 18748 5356 18760
rect 4479 18720 5356 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5552 18748 5580 18776
rect 5491 18720 5580 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 7006 18748 7012 18760
rect 6696 18720 7012 18748
rect 6696 18708 6702 18720
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 8220 18748 8248 18788
rect 8588 18757 8616 18788
rect 8662 18776 8668 18788
rect 8720 18776 8726 18828
rect 8938 18776 8944 18828
rect 8996 18816 9002 18828
rect 12342 18816 12348 18828
rect 8996 18788 12348 18816
rect 8996 18776 9002 18788
rect 12342 18776 12348 18788
rect 12400 18776 12406 18828
rect 12618 18776 12624 18828
rect 12676 18816 12682 18828
rect 12785 18819 12843 18825
rect 12785 18816 12797 18819
rect 12676 18788 12797 18816
rect 12676 18776 12682 18788
rect 12785 18785 12797 18788
rect 12831 18785 12843 18819
rect 12785 18779 12843 18785
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 17954 18816 17960 18828
rect 13136 18788 17960 18816
rect 13136 18776 13142 18788
rect 17954 18776 17960 18788
rect 18012 18776 18018 18828
rect 7116 18720 8248 18748
rect 8481 18751 8539 18757
rect 1949 18683 2007 18689
rect 1949 18649 1961 18683
rect 1995 18680 2007 18683
rect 5258 18680 5264 18692
rect 1995 18652 5264 18680
rect 1995 18649 2007 18652
rect 1949 18643 2007 18649
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 6822 18680 6828 18692
rect 6783 18652 6828 18680
rect 6822 18640 6828 18652
rect 6880 18640 6886 18692
rect 1486 18572 1492 18624
rect 1544 18612 1550 18624
rect 2958 18612 2964 18624
rect 1544 18584 2964 18612
rect 1544 18572 1550 18584
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3786 18572 3792 18624
rect 3844 18612 3850 18624
rect 7116 18612 7144 18720
rect 8481 18717 8493 18751
rect 8527 18717 8539 18751
rect 8481 18711 8539 18717
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 8573 18711 8631 18717
rect 7190 18640 7196 18692
rect 7248 18680 7254 18692
rect 8496 18680 8524 18711
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 9732 18720 10333 18748
rect 9732 18708 9738 18720
rect 10321 18717 10333 18720
rect 10367 18717 10379 18751
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 10321 18711 10379 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 16114 18708 16120 18760
rect 16172 18748 16178 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 16172 18720 16313 18748
rect 16172 18708 16178 18720
rect 16301 18717 16313 18720
rect 16347 18717 16359 18751
rect 18064 18748 18092 18856
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 18138 18776 18144 18828
rect 18196 18816 18202 18828
rect 18877 18819 18935 18825
rect 18877 18816 18889 18819
rect 18196 18788 18889 18816
rect 18196 18776 18202 18788
rect 18877 18785 18889 18788
rect 18923 18785 18935 18819
rect 18877 18779 18935 18785
rect 18966 18748 18972 18760
rect 16301 18711 16359 18717
rect 17328 18720 18092 18748
rect 18927 18720 18972 18748
rect 8754 18680 8760 18692
rect 7248 18652 8760 18680
rect 7248 18640 7254 18652
rect 8754 18640 8760 18652
rect 8812 18640 8818 18692
rect 11330 18640 11336 18692
rect 11388 18680 11394 18692
rect 11701 18683 11759 18689
rect 11701 18680 11713 18683
rect 11388 18652 11713 18680
rect 11388 18640 11394 18652
rect 11701 18649 11713 18652
rect 11747 18649 11759 18683
rect 11701 18643 11759 18649
rect 13538 18640 13544 18692
rect 13596 18680 13602 18692
rect 13596 18652 14780 18680
rect 13596 18640 13602 18652
rect 3844 18584 7144 18612
rect 8021 18615 8079 18621
rect 3844 18572 3850 18584
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 9122 18612 9128 18624
rect 8067 18584 9128 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 9306 18572 9312 18624
rect 9364 18612 9370 18624
rect 13170 18612 13176 18624
rect 9364 18584 13176 18612
rect 9364 18572 9370 18584
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 14642 18612 14648 18624
rect 13320 18584 14648 18612
rect 13320 18572 13326 18584
rect 14642 18572 14648 18584
rect 14700 18572 14706 18624
rect 14752 18612 14780 18652
rect 17328 18612 17356 18720
rect 18966 18708 18972 18720
rect 19024 18708 19030 18760
rect 19150 18748 19156 18760
rect 19111 18720 19156 18748
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 17681 18683 17739 18689
rect 17681 18649 17693 18683
rect 17727 18680 17739 18683
rect 19168 18680 19196 18708
rect 17727 18652 19196 18680
rect 17727 18649 17739 18652
rect 17681 18643 17739 18649
rect 14752 18584 17356 18612
rect 17586 18572 17592 18624
rect 17644 18612 17650 18624
rect 18138 18612 18144 18624
rect 17644 18584 18144 18612
rect 17644 18572 17650 18584
rect 18138 18572 18144 18584
rect 18196 18612 18202 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 18196 18584 18337 18612
rect 18196 18572 18202 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 18509 18615 18567 18621
rect 18509 18581 18521 18615
rect 18555 18612 18567 18615
rect 18782 18612 18788 18624
rect 18555 18584 18788 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 18782 18572 18788 18584
rect 18840 18572 18846 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 5166 18368 5172 18420
rect 5224 18408 5230 18420
rect 6638 18408 6644 18420
rect 5224 18380 6644 18408
rect 5224 18368 5230 18380
rect 6638 18368 6644 18380
rect 6696 18368 6702 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 6825 18411 6883 18417
rect 6825 18408 6837 18411
rect 6788 18380 6837 18408
rect 6788 18368 6794 18380
rect 6825 18377 6837 18380
rect 6871 18377 6883 18411
rect 6825 18371 6883 18377
rect 8202 18368 8208 18420
rect 8260 18408 8266 18420
rect 10686 18408 10692 18420
rect 8260 18380 10692 18408
rect 8260 18368 8266 18380
rect 10686 18368 10692 18380
rect 10744 18368 10750 18420
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 16022 18408 16028 18420
rect 10827 18380 16028 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 13725 18343 13783 18349
rect 5408 18312 13216 18340
rect 5408 18300 5414 18312
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 5810 18272 5816 18284
rect 5767 18244 5816 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 5810 18232 5816 18244
rect 5868 18232 5874 18284
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 6788 18244 7389 18272
rect 6788 18232 6794 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 9122 18272 9128 18284
rect 9083 18244 9128 18272
rect 7377 18235 7435 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9217 18275 9275 18281
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9490 18272 9496 18284
rect 9263 18244 9496 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 1394 18204 1400 18216
rect 1355 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18164 1458 18216
rect 2498 18204 2504 18216
rect 2459 18176 2504 18204
rect 2498 18164 2504 18176
rect 2556 18164 2562 18216
rect 2590 18164 2596 18216
rect 2648 18204 2654 18216
rect 5534 18204 5540 18216
rect 2648 18176 5304 18204
rect 5495 18176 5540 18204
rect 2648 18164 2654 18176
rect 2768 18139 2826 18145
rect 2768 18105 2780 18139
rect 2814 18136 2826 18139
rect 3510 18136 3516 18148
rect 2814 18108 3516 18136
rect 2814 18105 2826 18108
rect 2768 18099 2826 18105
rect 3510 18096 3516 18108
rect 3568 18096 3574 18148
rect 5276 18136 5304 18176
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 5994 18164 6000 18216
rect 6052 18204 6058 18216
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6052 18176 7205 18204
rect 6052 18164 6058 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7340 18176 8616 18204
rect 7340 18164 7346 18176
rect 8478 18136 8484 18148
rect 5276 18108 8484 18136
rect 8478 18096 8484 18108
rect 8536 18096 8542 18148
rect 8588 18136 8616 18176
rect 8846 18164 8852 18216
rect 8904 18204 8910 18216
rect 9232 18204 9260 18235
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 11054 18272 11060 18284
rect 9640 18244 11060 18272
rect 9640 18232 9646 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 11882 18272 11888 18284
rect 11471 18244 11888 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 13188 18272 13216 18312
rect 13725 18309 13737 18343
rect 13771 18340 13783 18343
rect 13771 18312 15792 18340
rect 13771 18309 13783 18312
rect 13725 18303 13783 18309
rect 13998 18272 14004 18284
rect 13188 18244 14004 18272
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14182 18272 14188 18284
rect 14143 18244 14188 18272
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 15764 18281 15792 18312
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16758 18272 16764 18284
rect 15979 18244 16764 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 20346 18232 20352 18284
rect 20404 18272 20410 18284
rect 20441 18275 20499 18281
rect 20441 18272 20453 18275
rect 20404 18244 20453 18272
rect 20404 18232 20410 18244
rect 20441 18241 20453 18244
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 11146 18204 11152 18216
rect 8904 18176 9260 18204
rect 11107 18176 11152 18204
rect 8904 18164 8910 18176
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 11790 18204 11796 18216
rect 11287 18176 11796 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 12434 18164 12440 18216
rect 12492 18204 12498 18216
rect 13078 18204 13084 18216
rect 12492 18176 12537 18204
rect 12636 18176 13084 18204
rect 12492 18164 12498 18176
rect 9033 18139 9091 18145
rect 9033 18136 9045 18139
rect 8588 18108 9045 18136
rect 9033 18105 9045 18108
rect 9079 18105 9091 18139
rect 9033 18099 9091 18105
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 12636 18136 12664 18176
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 15286 18164 15292 18216
rect 15344 18204 15350 18216
rect 15657 18207 15715 18213
rect 15657 18204 15669 18207
rect 15344 18176 15669 18204
rect 15344 18164 15350 18176
rect 15657 18173 15669 18176
rect 15703 18173 15715 18207
rect 15657 18167 15715 18173
rect 15838 18164 15844 18216
rect 15896 18204 15902 18216
rect 16853 18207 16911 18213
rect 16853 18204 16865 18207
rect 15896 18176 16865 18204
rect 15896 18164 15902 18176
rect 16853 18173 16865 18176
rect 16899 18173 16911 18207
rect 16853 18167 16911 18173
rect 17494 18164 17500 18216
rect 17552 18204 17558 18216
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17552 18176 18061 18204
rect 17552 18164 17558 18176
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18316 18207 18374 18213
rect 18316 18173 18328 18207
rect 18362 18204 18374 18207
rect 19150 18204 19156 18216
rect 18362 18176 19156 18204
rect 18362 18173 18374 18176
rect 18316 18167 18374 18173
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 20254 18204 20260 18216
rect 20215 18176 20260 18204
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 10928 18108 12664 18136
rect 12713 18139 12771 18145
rect 10928 18096 10934 18108
rect 12713 18105 12725 18139
rect 12759 18136 12771 18139
rect 13538 18136 13544 18148
rect 12759 18108 13544 18136
rect 12759 18105 12771 18108
rect 12713 18099 12771 18105
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 14090 18136 14096 18148
rect 14051 18108 14096 18136
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 15470 18136 15476 18148
rect 15304 18108 15476 18136
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 3786 18068 3792 18080
rect 1627 18040 3792 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 3786 18028 3792 18040
rect 3844 18028 3850 18080
rect 3881 18071 3939 18077
rect 3881 18037 3893 18071
rect 3927 18068 3939 18071
rect 4154 18068 4160 18080
rect 3927 18040 4160 18068
rect 3927 18037 3939 18040
rect 3881 18031 3939 18037
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5408 18040 5641 18068
rect 5408 18028 5414 18040
rect 5629 18037 5641 18040
rect 5675 18068 5687 18071
rect 7006 18068 7012 18080
rect 5675 18040 7012 18068
rect 5675 18037 5687 18040
rect 5629 18031 5687 18037
rect 7006 18028 7012 18040
rect 7064 18028 7070 18080
rect 7098 18028 7104 18080
rect 7156 18068 7162 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7156 18040 7297 18068
rect 7156 18028 7162 18040
rect 7285 18037 7297 18040
rect 7331 18037 7343 18071
rect 8662 18068 8668 18080
rect 8623 18040 8668 18068
rect 7285 18031 7343 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 12158 18068 12164 18080
rect 9180 18040 12164 18068
rect 9180 18028 9186 18040
rect 12158 18028 12164 18040
rect 12216 18028 12222 18080
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 13722 18068 13728 18080
rect 12584 18040 13728 18068
rect 12584 18028 12590 18040
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 15304 18077 15332 18108
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 15562 18096 15568 18148
rect 15620 18136 15626 18148
rect 19518 18136 19524 18148
rect 15620 18108 19524 18136
rect 15620 18096 15626 18108
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 15289 18071 15347 18077
rect 15289 18037 15301 18071
rect 15335 18037 15347 18071
rect 15289 18031 15347 18037
rect 17037 18071 17095 18077
rect 17037 18037 17049 18071
rect 17083 18068 17095 18071
rect 18138 18068 18144 18080
rect 17083 18040 18144 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 19426 18068 19432 18080
rect 19387 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 2869 17867 2927 17873
rect 2869 17864 2881 17867
rect 2832 17836 2881 17864
rect 2832 17824 2838 17836
rect 2869 17833 2881 17836
rect 2915 17833 2927 17867
rect 4338 17864 4344 17876
rect 2869 17827 2927 17833
rect 3344 17836 4344 17864
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 3344 17728 3372 17836
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 6178 17864 6184 17876
rect 6139 17836 6184 17864
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 12345 17867 12403 17873
rect 6328 17836 11468 17864
rect 6328 17824 6334 17836
rect 5534 17796 5540 17808
rect 2823 17700 3372 17728
rect 3436 17768 5540 17796
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 1412 17592 1440 17623
rect 2590 17620 2596 17672
rect 2648 17660 2654 17672
rect 3053 17663 3111 17669
rect 3053 17660 3065 17663
rect 2648 17632 3065 17660
rect 2648 17620 2654 17632
rect 3053 17629 3065 17632
rect 3099 17660 3111 17663
rect 3326 17660 3332 17672
rect 3099 17632 3332 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 3326 17620 3332 17632
rect 3384 17620 3390 17672
rect 3436 17592 3464 17768
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 5626 17756 5632 17808
rect 5684 17796 5690 17808
rect 6730 17796 6736 17808
rect 5684 17768 6736 17796
rect 5684 17756 5690 17768
rect 6730 17756 6736 17768
rect 6788 17756 6794 17808
rect 7006 17756 7012 17808
rect 7064 17796 7070 17808
rect 9953 17799 10011 17805
rect 9953 17796 9965 17799
rect 7064 17768 9965 17796
rect 7064 17756 7070 17768
rect 9953 17765 9965 17768
rect 9999 17765 10011 17799
rect 11440 17796 11468 17836
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 12618 17864 12624 17876
rect 12391 17836 12624 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 18417 17867 18475 17873
rect 18417 17833 18429 17867
rect 18463 17833 18475 17867
rect 18782 17864 18788 17876
rect 18743 17836 18788 17864
rect 18417 17827 18475 17833
rect 15194 17796 15200 17808
rect 11440 17768 15200 17796
rect 9953 17759 10011 17765
rect 15194 17756 15200 17768
rect 15252 17756 15258 17808
rect 18432 17796 18460 17827
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 19702 17796 19708 17808
rect 18432 17768 19708 17796
rect 19702 17756 19708 17768
rect 19760 17756 19766 17808
rect 4893 17731 4951 17737
rect 4893 17697 4905 17731
rect 4939 17728 4951 17731
rect 6454 17728 6460 17740
rect 4939 17700 6460 17728
rect 4939 17697 4951 17700
rect 4893 17691 4951 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6604 17700 6649 17728
rect 6604 17688 6610 17700
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5077 17623 5135 17629
rect 1412 17564 3464 17592
rect 3510 17552 3516 17604
rect 3568 17592 3574 17604
rect 4798 17592 4804 17604
rect 3568 17564 4804 17592
rect 3568 17552 3574 17564
rect 4798 17552 4804 17564
rect 4856 17592 4862 17604
rect 5092 17592 5120 17623
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 6748 17669 6776 17756
rect 7466 17688 7472 17740
rect 7524 17728 7530 17740
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 7524 17700 8217 17728
rect 7524 17688 7530 17700
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 9677 17731 9735 17737
rect 9677 17697 9689 17731
rect 9723 17728 9735 17731
rect 10134 17728 10140 17740
rect 9723 17700 10140 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 11238 17737 11244 17740
rect 11232 17728 11244 17737
rect 11199 17700 11244 17728
rect 11232 17691 11244 17700
rect 11238 17688 11244 17691
rect 11296 17688 11302 17740
rect 14001 17731 14059 17737
rect 14001 17697 14013 17731
rect 14047 17728 14059 17731
rect 14182 17728 14188 17740
rect 14047 17700 14188 17728
rect 14047 17697 14059 17700
rect 14001 17691 14059 17697
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 16384 17731 16442 17737
rect 16384 17697 16396 17731
rect 16430 17728 16442 17731
rect 19426 17728 19432 17740
rect 16430 17700 19432 17728
rect 16430 17697 16442 17700
rect 16384 17691 16442 17697
rect 6641 17663 6699 17669
rect 6641 17660 6653 17663
rect 5500 17632 6653 17660
rect 5500 17620 5506 17632
rect 6641 17629 6653 17632
rect 6687 17629 6699 17663
rect 6641 17623 6699 17629
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17629 6791 17663
rect 6733 17623 6791 17629
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7432 17632 8309 17660
rect 7432 17620 7438 17632
rect 8297 17629 8309 17632
rect 8343 17629 8355 17663
rect 8297 17623 8355 17629
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 10962 17660 10968 17672
rect 10923 17632 10968 17660
rect 8389 17623 8447 17629
rect 4856 17564 5120 17592
rect 4856 17552 4862 17564
rect 5258 17552 5264 17604
rect 5316 17592 5322 17604
rect 8404 17592 8432 17623
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 14090 17660 14096 17672
rect 14051 17632 14096 17660
rect 14090 17620 14096 17632
rect 14148 17620 14154 17672
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 16022 17660 16028 17672
rect 14323 17632 16028 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 16022 17620 16028 17632
rect 16080 17620 16086 17672
rect 16114 17620 16120 17672
rect 16172 17660 16178 17672
rect 18874 17660 18880 17672
rect 16172 17632 16217 17660
rect 18835 17632 18880 17660
rect 16172 17620 16178 17632
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 18984 17669 19012 17700
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 18969 17663 19027 17669
rect 18969 17629 18981 17663
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 5316 17564 8432 17592
rect 17497 17595 17555 17601
rect 5316 17552 5322 17564
rect 17497 17561 17509 17595
rect 17543 17592 17555 17595
rect 18598 17592 18604 17604
rect 17543 17564 18604 17592
rect 17543 17561 17555 17564
rect 17497 17555 17555 17561
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 2409 17527 2467 17533
rect 2409 17493 2421 17527
rect 2455 17524 2467 17527
rect 3694 17524 3700 17536
rect 2455 17496 3700 17524
rect 2455 17493 2467 17496
rect 2409 17487 2467 17493
rect 3694 17484 3700 17496
rect 3752 17484 3758 17536
rect 4525 17527 4583 17533
rect 4525 17493 4537 17527
rect 4571 17524 4583 17527
rect 4890 17524 4896 17536
rect 4571 17496 4896 17524
rect 4571 17493 4583 17496
rect 4525 17487 4583 17493
rect 4890 17484 4896 17496
rect 4948 17484 4954 17536
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 7837 17527 7895 17533
rect 7837 17524 7849 17527
rect 7708 17496 7849 17524
rect 7708 17484 7714 17496
rect 7837 17493 7849 17496
rect 7883 17493 7895 17527
rect 7837 17487 7895 17493
rect 8202 17484 8208 17536
rect 8260 17524 8266 17536
rect 12802 17524 12808 17536
rect 8260 17496 12808 17524
rect 8260 17484 8266 17496
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 13633 17527 13691 17533
rect 13633 17493 13645 17527
rect 13679 17524 13691 17527
rect 16482 17524 16488 17536
rect 13679 17496 16488 17524
rect 13679 17493 13691 17496
rect 13633 17487 13691 17493
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 17218 17484 17224 17536
rect 17276 17524 17282 17536
rect 17678 17524 17684 17536
rect 17276 17496 17684 17524
rect 17276 17484 17282 17496
rect 17678 17484 17684 17496
rect 17736 17484 17742 17536
rect 19794 17484 19800 17536
rect 19852 17524 19858 17536
rect 20438 17524 20444 17536
rect 19852 17496 20444 17524
rect 19852 17484 19858 17496
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20806 17484 20812 17536
rect 20864 17524 20870 17536
rect 22094 17524 22100 17536
rect 20864 17496 22100 17524
rect 20864 17484 20870 17496
rect 22094 17484 22100 17496
rect 22152 17484 22158 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3568 17292 3709 17320
rect 3568 17280 3574 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 3786 17280 3792 17332
rect 3844 17320 3850 17332
rect 6270 17320 6276 17332
rect 3844 17292 6276 17320
rect 3844 17280 3850 17292
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 6825 17323 6883 17329
rect 6825 17320 6837 17323
rect 6512 17292 6837 17320
rect 6512 17280 6518 17292
rect 6825 17289 6837 17292
rect 6871 17289 6883 17323
rect 9953 17323 10011 17329
rect 6825 17283 6883 17289
rect 7484 17292 9536 17320
rect 3326 17212 3332 17264
rect 3384 17252 3390 17264
rect 3384 17224 5856 17252
rect 3384 17212 3390 17224
rect 5828 17196 5856 17224
rect 6638 17212 6644 17264
rect 6696 17252 6702 17264
rect 7484 17252 7512 17292
rect 6696 17224 7512 17252
rect 9508 17252 9536 17292
rect 9953 17289 9965 17323
rect 9999 17320 10011 17323
rect 10042 17320 10048 17332
rect 9999 17292 10048 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 10686 17280 10692 17332
rect 10744 17320 10750 17332
rect 10744 17292 14044 17320
rect 10744 17280 10750 17292
rect 10781 17255 10839 17261
rect 10781 17252 10793 17255
rect 9508 17224 10793 17252
rect 6696 17212 6702 17224
rect 10781 17221 10793 17224
rect 10827 17221 10839 17255
rect 10781 17215 10839 17221
rect 11238 17212 11244 17264
rect 11296 17252 11302 17264
rect 11790 17252 11796 17264
rect 11296 17224 11796 17252
rect 11296 17212 11302 17224
rect 11790 17212 11796 17224
rect 11848 17252 11854 17264
rect 14016 17252 14044 17292
rect 14090 17280 14096 17332
rect 14148 17320 14154 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14148 17292 15117 17320
rect 14148 17280 14154 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 19613 17323 19671 17329
rect 19613 17320 19625 17323
rect 18932 17292 19625 17320
rect 18932 17280 18938 17292
rect 19613 17289 19625 17292
rect 19659 17289 19671 17323
rect 19613 17283 19671 17289
rect 20990 17280 20996 17332
rect 21048 17320 21054 17332
rect 22646 17320 22652 17332
rect 21048 17292 22652 17320
rect 21048 17280 21054 17292
rect 22646 17280 22652 17292
rect 22704 17280 22710 17332
rect 14185 17255 14243 17261
rect 11848 17224 13032 17252
rect 14016 17224 14136 17252
rect 11848 17212 11854 17224
rect 4154 17144 4160 17196
rect 4212 17184 4218 17196
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 4212 17156 5089 17184
rect 4212 17144 4218 17156
rect 5077 17153 5089 17156
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 5810 17144 5816 17196
rect 5868 17184 5874 17196
rect 7469 17187 7527 17193
rect 7469 17184 7481 17187
rect 5868 17156 7481 17184
rect 5868 17144 5874 17156
rect 7469 17153 7481 17156
rect 7515 17184 7527 17187
rect 7742 17184 7748 17196
rect 7515 17156 7748 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 8352 17156 8585 17184
rect 8352 17144 8358 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 11425 17187 11483 17193
rect 11425 17153 11437 17187
rect 11471 17184 11483 17187
rect 12618 17184 12624 17196
rect 11471 17156 12624 17184
rect 11471 17153 11483 17156
rect 11425 17147 11483 17153
rect 12618 17144 12624 17156
rect 12676 17144 12682 17196
rect 13004 17193 13032 17224
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 2590 17125 2596 17128
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2584 17079 2596 17125
rect 2648 17116 2654 17128
rect 4890 17116 4896 17128
rect 2648 17088 2684 17116
rect 4851 17088 4896 17116
rect 2332 17048 2360 17079
rect 2590 17076 2596 17079
rect 2648 17076 2654 17088
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 7098 17116 7104 17128
rect 5368 17088 7104 17116
rect 2498 17048 2504 17060
rect 2332 17020 2504 17048
rect 2498 17008 2504 17020
rect 2556 17048 2562 17060
rect 2866 17048 2872 17060
rect 2556 17020 2872 17048
rect 2556 17008 2562 17020
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 5368 17048 5396 17088
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 8478 17116 8484 17128
rect 7239 17088 8484 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 8478 17076 8484 17088
rect 8536 17076 8542 17128
rect 12802 17116 12808 17128
rect 8588 17088 12664 17116
rect 12763 17088 12808 17116
rect 4080 17020 5396 17048
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 4080 16980 4108 17020
rect 5442 17008 5448 17060
rect 5500 17048 5506 17060
rect 8588 17048 8616 17088
rect 8846 17057 8852 17060
rect 8840 17048 8852 17057
rect 5500 17020 8616 17048
rect 8807 17020 8852 17048
rect 5500 17008 5506 17020
rect 8840 17011 8852 17020
rect 8846 17008 8852 17011
rect 8904 17008 8910 17060
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 12636 17048 12664 17088
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13998 17116 14004 17128
rect 13959 17088 14004 17116
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 14108 17116 14136 17224
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 17862 17252 17868 17264
rect 14231 17224 17868 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 17972 17224 19012 17252
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 14608 17156 15669 17184
rect 14608 17144 14614 17156
rect 15657 17153 15669 17156
rect 15703 17153 15715 17187
rect 17972 17184 18000 17224
rect 18598 17184 18604 17196
rect 15657 17147 15715 17153
rect 15764 17156 18000 17184
rect 18559 17156 18604 17184
rect 14458 17116 14464 17128
rect 14108 17088 14464 17116
rect 14458 17076 14464 17088
rect 14516 17116 14522 17128
rect 15764 17116 15792 17156
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 14516 17088 15792 17116
rect 14516 17076 14522 17088
rect 16482 17076 16488 17128
rect 16540 17116 16546 17128
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16540 17088 16681 17116
rect 16540 17076 16546 17088
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 18417 17119 18475 17125
rect 18417 17116 18429 17119
rect 16669 17079 16727 17085
rect 16776 17088 18429 17116
rect 16776 17048 16804 17088
rect 18417 17085 18429 17088
rect 18463 17116 18475 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 18463 17088 18889 17116
rect 18463 17085 18475 17088
rect 18417 17079 18475 17085
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 18984 17116 19012 17224
rect 19334 17212 19340 17264
rect 19392 17252 19398 17264
rect 20438 17252 20444 17264
rect 19392 17224 20444 17252
rect 19392 17212 19398 17224
rect 20438 17212 20444 17224
rect 20496 17212 20502 17264
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19208 17156 20177 17184
rect 19208 17144 19214 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 20073 17119 20131 17125
rect 20073 17116 20085 17119
rect 18984 17088 20085 17116
rect 18877 17079 18935 17085
rect 20073 17085 20085 17088
rect 20119 17085 20131 17119
rect 20073 17079 20131 17085
rect 11195 17020 12480 17048
rect 12636 17020 16804 17048
rect 16945 17051 17003 17057
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 1636 16952 4108 16980
rect 1636 16940 1642 16952
rect 4154 16940 4160 16992
rect 4212 16980 4218 16992
rect 4525 16983 4583 16989
rect 4525 16980 4537 16983
rect 4212 16952 4537 16980
rect 4212 16940 4218 16952
rect 4525 16949 4537 16952
rect 4571 16949 4583 16983
rect 4525 16943 4583 16949
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 4985 16983 5043 16989
rect 4985 16980 4997 16983
rect 4948 16952 4997 16980
rect 4948 16940 4954 16952
rect 4985 16949 4997 16952
rect 5031 16949 5043 16983
rect 4985 16943 5043 16949
rect 6270 16940 6276 16992
rect 6328 16980 6334 16992
rect 7006 16980 7012 16992
rect 6328 16952 7012 16980
rect 6328 16940 6334 16952
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 7285 16983 7343 16989
rect 7285 16949 7297 16983
rect 7331 16980 7343 16983
rect 10410 16980 10416 16992
rect 7331 16952 10416 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 12452 16989 12480 17020
rect 16945 17017 16957 17051
rect 16991 17048 17003 17051
rect 17034 17048 17040 17060
rect 16991 17020 17040 17048
rect 16991 17017 17003 17020
rect 16945 17011 17003 17017
rect 17034 17008 17040 17020
rect 17092 17008 17098 17060
rect 17586 17008 17592 17060
rect 17644 17048 17650 17060
rect 18509 17051 18567 17057
rect 18509 17048 18521 17051
rect 17644 17020 18521 17048
rect 17644 17008 17650 17020
rect 18509 17017 18521 17020
rect 18555 17017 18567 17051
rect 18509 17011 18567 17017
rect 19981 17051 20039 17057
rect 19981 17017 19993 17051
rect 20027 17048 20039 17051
rect 20346 17048 20352 17060
rect 20027 17020 20352 17048
rect 20027 17017 20039 17020
rect 19981 17011 20039 17017
rect 20346 17008 20352 17020
rect 20404 17008 20410 17060
rect 12437 16983 12495 16989
rect 11296 16952 11341 16980
rect 11296 16940 11302 16952
rect 12437 16949 12449 16983
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 12897 16983 12955 16989
rect 12897 16949 12909 16983
rect 12943 16980 12955 16983
rect 13354 16980 13360 16992
rect 12943 16952 13360 16980
rect 12943 16949 12955 16952
rect 12897 16943 12955 16949
rect 13354 16940 13360 16952
rect 13412 16940 13418 16992
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 15473 16983 15531 16989
rect 15473 16980 15485 16983
rect 14424 16952 15485 16980
rect 14424 16940 14430 16952
rect 15473 16949 15485 16952
rect 15519 16949 15531 16983
rect 15473 16943 15531 16949
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 18046 16980 18052 16992
rect 15620 16952 15665 16980
rect 18007 16952 18052 16980
rect 15620 16940 15626 16952
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 1762 16776 1768 16788
rect 1723 16748 1768 16776
rect 1762 16736 1768 16748
rect 1820 16736 1826 16788
rect 4525 16779 4583 16785
rect 4525 16745 4537 16779
rect 4571 16776 4583 16779
rect 11238 16776 11244 16788
rect 4571 16748 4752 16776
rect 11199 16748 11244 16776
rect 4571 16745 4583 16748
rect 4525 16739 4583 16745
rect 2961 16711 3019 16717
rect 2961 16677 2973 16711
rect 3007 16708 3019 16711
rect 3786 16708 3792 16720
rect 3007 16680 3792 16708
rect 3007 16677 3019 16680
rect 2961 16671 3019 16677
rect 3786 16668 3792 16680
rect 3844 16668 3850 16720
rect 4617 16711 4675 16717
rect 4617 16708 4629 16711
rect 4540 16680 4629 16708
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 2498 16640 2504 16652
rect 1627 16612 2504 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16609 2743 16643
rect 2685 16603 2743 16609
rect 2700 16572 2728 16603
rect 3694 16600 3700 16652
rect 3752 16640 3758 16652
rect 4540 16640 4568 16680
rect 4617 16677 4629 16680
rect 4663 16677 4675 16711
rect 4724 16708 4752 16748
rect 11238 16736 11244 16748
rect 11296 16736 11302 16788
rect 11698 16776 11704 16788
rect 11659 16748 11704 16776
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 11940 16748 14381 16776
rect 11940 16736 11946 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 19061 16779 19119 16785
rect 19061 16776 19073 16779
rect 18104 16748 19073 16776
rect 18104 16736 18110 16748
rect 19061 16745 19073 16748
rect 19107 16745 19119 16779
rect 19061 16739 19119 16745
rect 5166 16708 5172 16720
rect 4724 16680 5172 16708
rect 4617 16671 4675 16677
rect 5166 16668 5172 16680
rect 5224 16668 5230 16720
rect 6822 16668 6828 16720
rect 6880 16668 6886 16720
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 15562 16708 15568 16720
rect 7064 16680 15568 16708
rect 7064 16668 7070 16680
rect 15562 16668 15568 16680
rect 15620 16668 15626 16720
rect 16752 16711 16810 16717
rect 16752 16677 16764 16711
rect 16798 16708 16810 16711
rect 18598 16708 18604 16720
rect 16798 16680 18604 16708
rect 16798 16677 16810 16680
rect 16752 16671 16810 16677
rect 18598 16668 18604 16680
rect 18656 16668 18662 16720
rect 6840 16640 6868 16668
rect 3752 16612 4568 16640
rect 4632 16612 6868 16640
rect 6908 16643 6966 16649
rect 3752 16600 3758 16612
rect 4632 16572 4660 16612
rect 6908 16609 6920 16643
rect 6954 16640 6966 16643
rect 7282 16640 7288 16652
rect 6954 16612 7288 16640
rect 6954 16609 6966 16612
rect 6908 16603 6966 16609
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7834 16600 7840 16652
rect 7892 16640 7898 16652
rect 8202 16640 8208 16652
rect 7892 16612 8208 16640
rect 7892 16600 7898 16612
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 8444 16612 10057 16640
rect 8444 16600 8450 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16640 10195 16643
rect 11146 16640 11152 16652
rect 10183 16612 11152 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11296 16612 11621 16640
rect 11296 16600 11302 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12894 16640 12900 16652
rect 11756 16612 12900 16640
rect 11756 16600 11762 16612
rect 12894 16600 12900 16612
rect 12952 16640 12958 16652
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 12952 16612 13001 16640
rect 12952 16600 12958 16612
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 13256 16643 13314 16649
rect 13256 16609 13268 16643
rect 13302 16640 13314 16643
rect 13302 16612 14044 16640
rect 13302 16609 13314 16612
rect 13256 16603 13314 16609
rect 4798 16572 4804 16584
rect 2700 16544 4660 16572
rect 4759 16544 4804 16572
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 5626 16532 5632 16584
rect 5684 16572 5690 16584
rect 6641 16575 6699 16581
rect 6641 16572 6653 16575
rect 5684 16544 6653 16572
rect 5684 16532 5690 16544
rect 6641 16541 6653 16544
rect 6687 16541 6699 16575
rect 6641 16535 6699 16541
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 8904 16544 10241 16572
rect 8904 16532 8910 16544
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 10229 16535 10287 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 14016 16572 14044 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 15252 16612 15393 16640
rect 15252 16600 15258 16612
rect 15381 16609 15393 16612
rect 15427 16609 15439 16643
rect 18046 16640 18052 16652
rect 15381 16603 15439 16609
rect 15580 16612 18052 16640
rect 14734 16572 14740 16584
rect 14016 16544 14740 16572
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 4157 16507 4215 16513
rect 4157 16473 4169 16507
rect 4203 16504 4215 16507
rect 4890 16504 4896 16516
rect 4203 16476 4896 16504
rect 4203 16473 4215 16476
rect 4157 16467 4215 16473
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 15580 16513 15608 16612
rect 18046 16600 18052 16612
rect 18104 16600 18110 16652
rect 20254 16640 20260 16652
rect 18708 16612 20260 16640
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16482 16572 16488 16584
rect 16172 16544 16488 16572
rect 16172 16532 16178 16544
rect 16482 16532 16488 16544
rect 16540 16532 16546 16584
rect 18708 16513 18736 16612
rect 20254 16600 20260 16612
rect 20312 16600 20318 16652
rect 19150 16572 19156 16584
rect 19111 16544 19156 16572
rect 19150 16532 19156 16544
rect 19208 16532 19214 16584
rect 19245 16575 19303 16581
rect 19245 16541 19257 16575
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 15565 16507 15623 16513
rect 7576 16476 13032 16504
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 7576 16436 7604 16476
rect 1820 16408 7604 16436
rect 1820 16396 1826 16408
rect 7742 16396 7748 16448
rect 7800 16436 7806 16448
rect 8021 16439 8079 16445
rect 8021 16436 8033 16439
rect 7800 16408 8033 16436
rect 7800 16396 7806 16408
rect 8021 16405 8033 16408
rect 8067 16405 8079 16439
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 8021 16399 8079 16405
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9858 16396 9864 16448
rect 9916 16436 9922 16448
rect 11238 16436 11244 16448
rect 9916 16408 11244 16436
rect 9916 16396 9922 16408
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 13004 16436 13032 16476
rect 15565 16473 15577 16507
rect 15611 16473 15623 16507
rect 15565 16467 15623 16473
rect 18693 16507 18751 16513
rect 18693 16473 18705 16507
rect 18739 16473 18751 16507
rect 18693 16467 18751 16473
rect 16850 16436 16856 16448
rect 13004 16408 16856 16436
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 17865 16439 17923 16445
rect 17865 16436 17877 16439
rect 17828 16408 17877 16436
rect 17828 16396 17834 16408
rect 17865 16405 17877 16408
rect 17911 16436 17923 16439
rect 19260 16436 19288 16535
rect 17911 16408 19288 16436
rect 17911 16405 17923 16408
rect 17865 16399 17923 16405
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 5040 16204 5181 16232
rect 5040 16192 5046 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6362 16232 6368 16244
rect 6052 16204 6368 16232
rect 6052 16192 6058 16204
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 6454 16192 6460 16244
rect 6512 16232 6518 16244
rect 7006 16232 7012 16244
rect 6512 16204 7012 16232
rect 6512 16192 6518 16204
rect 7006 16192 7012 16204
rect 7064 16232 7070 16244
rect 12621 16235 12679 16241
rect 7064 16204 10364 16232
rect 7064 16192 7070 16204
rect 9033 16167 9091 16173
rect 9033 16164 9045 16167
rect 2332 16136 9045 16164
rect 2332 16037 2360 16136
rect 9033 16133 9045 16136
rect 9079 16133 9091 16167
rect 9033 16127 9091 16133
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 4065 16099 4123 16105
rect 4065 16096 4077 16099
rect 3016 16068 4077 16096
rect 3016 16056 3022 16068
rect 4065 16065 4077 16068
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 5258 16096 5264 16108
rect 4295 16068 5264 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5810 16096 5816 16108
rect 5771 16068 5816 16096
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 6236 16068 7389 16096
rect 6236 16056 6242 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 8662 16056 8668 16108
rect 8720 16096 8726 16108
rect 9493 16099 9551 16105
rect 9493 16096 9505 16099
rect 8720 16068 9505 16096
rect 8720 16056 8726 16068
rect 9493 16065 9505 16068
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 9950 16096 9956 16108
rect 9631 16068 9956 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 2317 15991 2375 15997
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 3970 16028 3976 16040
rect 3660 16000 3976 16028
rect 3660 15988 3666 16000
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 5537 16031 5595 16037
rect 5537 15997 5549 16031
rect 5583 16028 5595 16031
rect 5718 16028 5724 16040
rect 5583 16000 5724 16028
rect 5583 15997 5595 16000
rect 5537 15991 5595 15997
rect 5718 15988 5724 16000
rect 5776 16028 5782 16040
rect 6362 16028 6368 16040
rect 5776 16000 6368 16028
rect 5776 15988 5782 16000
rect 6362 15988 6368 16000
rect 6420 15988 6426 16040
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 8573 16031 8631 16037
rect 8573 16028 8585 16031
rect 6972 16000 8585 16028
rect 6972 15988 6978 16000
rect 8573 15997 8585 16000
rect 8619 15997 8631 16031
rect 8573 15991 8631 15997
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 16028 9459 16031
rect 9674 16028 9680 16040
rect 9447 16000 9680 16028
rect 9447 15997 9459 16000
rect 9401 15991 9459 15997
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 10336 16028 10364 16204
rect 12621 16201 12633 16235
rect 12667 16232 12679 16235
rect 14366 16232 14372 16244
rect 12667 16204 14372 16232
rect 12667 16201 12679 16204
rect 12621 16195 12679 16201
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15565 16235 15623 16241
rect 15565 16232 15577 16235
rect 14884 16204 15577 16232
rect 14884 16192 14890 16204
rect 15565 16201 15577 16204
rect 15611 16201 15623 16235
rect 15565 16195 15623 16201
rect 16482 16192 16488 16244
rect 16540 16232 16546 16244
rect 17494 16232 17500 16244
rect 16540 16204 17500 16232
rect 16540 16192 16546 16204
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18049 16235 18107 16241
rect 18049 16201 18061 16235
rect 18095 16232 18107 16235
rect 19150 16232 19156 16244
rect 18095 16204 19156 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 19978 16232 19984 16244
rect 19935 16204 19984 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 12952 16136 14228 16164
rect 12952 16124 12958 16136
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11422 16096 11428 16108
rect 10928 16068 11428 16096
rect 10928 16056 10934 16068
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 13265 16099 13323 16105
rect 13265 16065 13277 16099
rect 13311 16096 13323 16099
rect 13722 16096 13728 16108
rect 13311 16068 13728 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 14200 16105 14228 16136
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 20162 16164 20168 16176
rect 15344 16136 20168 16164
rect 15344 16124 15350 16136
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 16482 16056 16488 16108
rect 16540 16096 16546 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16540 16068 16957 16096
rect 16540 16056 16546 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 18598 16096 18604 16108
rect 18559 16068 18604 16096
rect 16945 16059 17003 16065
rect 18598 16056 18604 16068
rect 18656 16056 18662 16108
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 10336 16000 14688 16028
rect 2590 15960 2596 15972
rect 2551 15932 2596 15960
rect 2590 15920 2596 15932
rect 2648 15920 2654 15972
rect 7285 15963 7343 15969
rect 7285 15960 7297 15963
rect 3620 15932 7297 15960
rect 3620 15901 3648 15932
rect 7285 15929 7297 15932
rect 7331 15929 7343 15963
rect 7285 15923 7343 15929
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 11698 15960 11704 15972
rect 11195 15932 11704 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 11698 15920 11704 15932
rect 11756 15920 11762 15972
rect 14458 15969 14464 15972
rect 12989 15963 13047 15969
rect 12989 15929 13001 15963
rect 13035 15960 13047 15963
rect 13035 15932 14412 15960
rect 13035 15929 13047 15932
rect 12989 15923 13047 15929
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15861 3663 15895
rect 3605 15855 3663 15861
rect 5629 15895 5687 15901
rect 5629 15861 5641 15895
rect 5675 15892 5687 15895
rect 6454 15892 6460 15904
rect 5675 15864 6460 15892
rect 5675 15861 5687 15864
rect 5629 15855 5687 15861
rect 6454 15852 6460 15864
rect 6512 15852 6518 15904
rect 6822 15892 6828 15904
rect 6783 15864 6828 15892
rect 6822 15852 6828 15864
rect 6880 15852 6886 15904
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 8294 15852 8300 15904
rect 8352 15892 8358 15904
rect 8389 15895 8447 15901
rect 8389 15892 8401 15895
rect 8352 15864 8401 15892
rect 8352 15852 8358 15864
rect 8389 15861 8401 15864
rect 8435 15892 8447 15895
rect 9214 15892 9220 15904
rect 8435 15864 9220 15892
rect 8435 15861 8447 15864
rect 8389 15855 8447 15861
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 9950 15852 9956 15904
rect 10008 15892 10014 15904
rect 10502 15892 10508 15904
rect 10008 15864 10508 15892
rect 10008 15852 10014 15864
rect 10502 15852 10508 15864
rect 10560 15852 10566 15904
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 10781 15895 10839 15901
rect 10781 15892 10793 15895
rect 10652 15864 10793 15892
rect 10652 15852 10658 15864
rect 10781 15861 10793 15864
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11296 15864 11341 15892
rect 11296 15852 11302 15864
rect 11422 15852 11428 15904
rect 11480 15892 11486 15904
rect 12618 15892 12624 15904
rect 11480 15864 12624 15892
rect 11480 15852 11486 15864
rect 12618 15852 12624 15864
rect 12676 15852 12682 15904
rect 13081 15895 13139 15901
rect 13081 15861 13093 15895
rect 13127 15892 13139 15895
rect 13998 15892 14004 15904
rect 13127 15864 14004 15892
rect 13127 15861 13139 15864
rect 13081 15855 13139 15861
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 14384 15892 14412 15932
rect 14452 15923 14464 15969
rect 14516 15960 14522 15972
rect 14660 15960 14688 16000
rect 16758 15988 16764 16040
rect 16816 16028 16822 16040
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16816 16000 16865 16028
rect 16816 15988 16822 16000
rect 16853 15997 16865 16000
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 17460 16000 18521 16028
rect 17460 15988 17466 16000
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 20456 16028 20484 16059
rect 19300 16000 20484 16028
rect 19300 15988 19306 16000
rect 18417 15963 18475 15969
rect 18417 15960 18429 15963
rect 14516 15932 14552 15960
rect 14660 15932 18429 15960
rect 14458 15920 14464 15923
rect 14516 15920 14522 15932
rect 18417 15929 18429 15932
rect 18463 15929 18475 15963
rect 18417 15923 18475 15929
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 20349 15963 20407 15969
rect 20349 15960 20361 15963
rect 19392 15932 20361 15960
rect 19392 15920 19398 15932
rect 20349 15929 20361 15932
rect 20395 15929 20407 15963
rect 20349 15923 20407 15929
rect 15562 15892 15568 15904
rect 14384 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 16393 15895 16451 15901
rect 16393 15861 16405 15895
rect 16439 15892 16451 15895
rect 16666 15892 16672 15904
rect 16439 15864 16672 15892
rect 16439 15861 16451 15864
rect 16393 15855 16451 15861
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 16850 15892 16856 15904
rect 16807 15864 16856 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 16850 15852 16856 15864
rect 16908 15852 16914 15904
rect 19797 15895 19855 15901
rect 19797 15861 19809 15895
rect 19843 15892 19855 15895
rect 20254 15892 20260 15904
rect 19843 15864 20260 15892
rect 19843 15861 19855 15864
rect 19797 15855 19855 15861
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 1762 15688 1768 15700
rect 1723 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7098 15688 7104 15700
rect 6880 15660 7104 15688
rect 6880 15648 6886 15660
rect 7098 15648 7104 15660
rect 7156 15648 7162 15700
rect 7282 15688 7288 15700
rect 7243 15660 7288 15688
rect 7282 15648 7288 15660
rect 7340 15688 7346 15700
rect 7558 15688 7564 15700
rect 7340 15660 7564 15688
rect 7340 15648 7346 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 10594 15688 10600 15700
rect 10555 15660 10600 15688
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 16850 15688 16856 15700
rect 15252 15660 16856 15688
rect 15252 15648 15258 15660
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 17862 15648 17868 15700
rect 17920 15688 17926 15700
rect 19610 15688 19616 15700
rect 17920 15660 19616 15688
rect 17920 15648 17926 15660
rect 19610 15648 19616 15660
rect 19668 15648 19674 15700
rect 2961 15623 3019 15629
rect 2961 15589 2973 15623
rect 3007 15620 3019 15623
rect 3326 15620 3332 15632
rect 3007 15592 3332 15620
rect 3007 15589 3019 15592
rect 2961 15583 3019 15589
rect 3326 15580 3332 15592
rect 3384 15580 3390 15632
rect 4709 15623 4767 15629
rect 4709 15589 4721 15623
rect 4755 15620 4767 15623
rect 5534 15620 5540 15632
rect 4755 15592 5540 15620
rect 4755 15589 4767 15592
rect 4709 15583 4767 15589
rect 5534 15580 5540 15592
rect 5592 15580 5598 15632
rect 6178 15629 6184 15632
rect 6172 15583 6184 15629
rect 6236 15620 6242 15632
rect 8570 15620 8576 15632
rect 6236 15592 6272 15620
rect 8531 15592 8576 15620
rect 6178 15580 6184 15583
rect 6236 15580 6242 15592
rect 8570 15580 8576 15592
rect 8628 15580 8634 15632
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 15838 15620 15844 15632
rect 8720 15592 15844 15620
rect 8720 15580 8726 15592
rect 15838 15580 15844 15592
rect 15896 15580 15902 15632
rect 16301 15623 16359 15629
rect 16301 15620 16313 15623
rect 16224 15592 16313 15620
rect 1578 15552 1584 15564
rect 1539 15524 1584 15552
rect 1578 15512 1584 15524
rect 1636 15512 1642 15564
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15552 2743 15555
rect 4154 15552 4160 15564
rect 2731 15524 4160 15552
rect 2731 15521 2743 15524
rect 2685 15515 2743 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4801 15555 4859 15561
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5350 15552 5356 15564
rect 4847 15524 5356 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 8202 15552 8208 15564
rect 5951 15524 8208 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 10502 15552 10508 15564
rect 10463 15524 10508 15552
rect 8297 15515 8355 15521
rect 4985 15487 5043 15493
rect 4985 15453 4997 15487
rect 5031 15484 5043 15487
rect 5258 15484 5264 15496
rect 5031 15456 5264 15484
rect 5031 15453 5043 15456
rect 4985 15447 5043 15453
rect 5258 15444 5264 15456
rect 5316 15444 5322 15496
rect 2958 15376 2964 15428
rect 3016 15416 3022 15428
rect 5442 15416 5448 15428
rect 3016 15388 5448 15416
rect 3016 15376 3022 15388
rect 5442 15376 5448 15388
rect 5500 15376 5506 15428
rect 8312 15416 8340 15515
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 12049 15555 12107 15561
rect 12049 15552 12061 15555
rect 11940 15524 12061 15552
rect 11940 15512 11946 15524
rect 12049 15521 12061 15524
rect 12095 15521 12107 15555
rect 12049 15515 12107 15521
rect 14093 15555 14151 15561
rect 14093 15521 14105 15555
rect 14139 15552 14151 15555
rect 14274 15552 14280 15564
rect 14139 15524 14280 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 15286 15552 15292 15564
rect 14516 15524 15292 15552
rect 14516 15512 14522 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 16224 15552 16252 15592
rect 16301 15589 16313 15592
rect 16347 15589 16359 15623
rect 16301 15583 16359 15589
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 17460 15592 19748 15620
rect 17460 15580 17466 15592
rect 17770 15561 17776 15564
rect 17764 15552 17776 15561
rect 15436 15524 16252 15552
rect 17731 15524 17776 15552
rect 15436 15512 15442 15524
rect 17764 15515 17776 15524
rect 17770 15512 17776 15515
rect 17828 15512 17834 15564
rect 19720 15561 19748 15592
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 10689 15487 10747 15493
rect 10689 15484 10701 15487
rect 10652 15456 10701 15484
rect 10652 15444 10658 15456
rect 10689 15453 10701 15456
rect 10735 15453 10747 15487
rect 11790 15484 11796 15496
rect 11751 15456 11796 15484
rect 10689 15447 10747 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16482 15444 16488 15496
rect 16540 15484 16546 15496
rect 17494 15484 17500 15496
rect 16540 15456 16585 15484
rect 17455 15456 17500 15484
rect 16540 15444 16546 15456
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 10137 15419 10195 15425
rect 10137 15416 10149 15419
rect 8312 15388 10149 15416
rect 10137 15385 10149 15388
rect 10183 15385 10195 15419
rect 14277 15419 14335 15425
rect 10137 15379 10195 15385
rect 13004 15388 13299 15416
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 6822 15348 6828 15360
rect 4387 15320 6828 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 6822 15308 6828 15320
rect 6880 15308 6886 15360
rect 7282 15308 7288 15360
rect 7340 15348 7346 15360
rect 13004 15348 13032 15388
rect 13170 15348 13176 15360
rect 7340 15320 13032 15348
rect 13131 15320 13176 15348
rect 7340 15308 7346 15320
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13271 15348 13299 15388
rect 14277 15385 14289 15419
rect 14323 15416 14335 15419
rect 14323 15388 17540 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 15654 15348 15660 15360
rect 13271 15320 15660 15348
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 15933 15351 15991 15357
rect 15933 15317 15945 15351
rect 15979 15348 15991 15351
rect 16574 15348 16580 15360
rect 15979 15320 16580 15348
rect 15979 15317 15991 15320
rect 15933 15311 15991 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 17512 15348 17540 15388
rect 18782 15348 18788 15360
rect 17512 15320 18788 15348
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 18877 15351 18935 15357
rect 18877 15317 18889 15351
rect 18923 15348 18935 15351
rect 19242 15348 19248 15360
rect 18923 15320 19248 15348
rect 18923 15317 18935 15320
rect 18877 15311 18935 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 19886 15348 19892 15360
rect 19847 15320 19892 15348
rect 19886 15308 19892 15320
rect 19944 15308 19950 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 5077 15147 5135 15153
rect 5077 15144 5089 15147
rect 2792 15116 5089 15144
rect 2792 15017 2820 15116
rect 5077 15113 5089 15116
rect 5123 15144 5135 15147
rect 5258 15144 5264 15156
rect 5123 15116 5264 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 5776 15116 6377 15144
rect 5776 15104 5782 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 7282 15144 7288 15156
rect 6512 15116 7288 15144
rect 6512 15104 6518 15116
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 7653 15147 7711 15153
rect 7653 15113 7665 15147
rect 7699 15144 7711 15147
rect 11238 15144 11244 15156
rect 7699 15116 11244 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 12676 15116 13829 15144
rect 12676 15104 12682 15116
rect 13817 15113 13829 15116
rect 13863 15113 13875 15147
rect 13817 15107 13875 15113
rect 14645 15147 14703 15153
rect 14645 15113 14657 15147
rect 14691 15144 14703 15147
rect 15194 15144 15200 15156
rect 14691 15116 15200 15144
rect 14691 15113 14703 15116
rect 14645 15107 14703 15113
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15144 16267 15147
rect 16942 15144 16948 15156
rect 16255 15116 16948 15144
rect 16255 15113 16267 15116
rect 16209 15107 16267 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20162 15144 20168 15156
rect 20027 15116 20168 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 10594 15076 10600 15088
rect 10555 15048 10600 15076
rect 10594 15036 10600 15048
rect 10652 15036 10658 15088
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 7190 15008 7196 15020
rect 2777 14971 2835 14977
rect 4724 14980 7196 15008
rect 2501 14943 2559 14949
rect 2501 14909 2513 14943
rect 2547 14940 2559 14943
rect 3418 14940 3424 14952
rect 2547 14912 3424 14940
rect 2547 14909 2559 14912
rect 2501 14903 2559 14909
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 3694 14940 3700 14952
rect 3655 14912 3700 14940
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 4724 14940 4752 14980
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 8297 15011 8355 15017
rect 8297 14977 8309 15011
rect 8343 15008 8355 15011
rect 15286 15008 15292 15020
rect 8343 14980 9352 15008
rect 8343 14977 8355 14980
rect 8297 14971 8355 14977
rect 9324 14952 9352 14980
rect 12268 14980 12572 15008
rect 15247 14980 15292 15008
rect 3896 14912 4752 14940
rect 6549 14943 6607 14949
rect 3896 14872 3924 14912
rect 6549 14909 6561 14943
rect 6595 14940 6607 14943
rect 6914 14940 6920 14952
rect 6595 14912 6920 14940
rect 6595 14909 6607 14912
rect 6549 14903 6607 14909
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 9214 14940 9220 14952
rect 9175 14912 9220 14940
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 9306 14900 9312 14952
rect 9364 14900 9370 14952
rect 10778 14940 10784 14952
rect 9416 14912 10784 14940
rect 2148 14844 3924 14872
rect 3964 14875 4022 14881
rect 2148 14813 2176 14844
rect 3964 14841 3976 14875
rect 4010 14872 4022 14875
rect 4062 14872 4068 14884
rect 4010 14844 4068 14872
rect 4010 14841 4022 14844
rect 3964 14835 4022 14841
rect 4062 14832 4068 14844
rect 4120 14832 4126 14884
rect 4816 14844 6592 14872
rect 2133 14807 2191 14813
rect 2133 14773 2145 14807
rect 2179 14773 2191 14807
rect 2133 14767 2191 14773
rect 2593 14807 2651 14813
rect 2593 14773 2605 14807
rect 2639 14804 2651 14807
rect 4816 14804 4844 14844
rect 6564 14816 6592 14844
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 7742 14872 7748 14884
rect 7248 14844 7748 14872
rect 7248 14832 7254 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 8113 14875 8171 14881
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 9416 14872 9444 14912
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 12268 14949 12296 14980
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14909 12311 14943
rect 12253 14903 12311 14909
rect 12342 14900 12348 14952
rect 12400 14940 12406 14952
rect 12437 14943 12495 14949
rect 12437 14940 12449 14943
rect 12400 14912 12449 14940
rect 12400 14900 12406 14912
rect 12437 14909 12449 14912
rect 12483 14909 12495 14943
rect 12544 14940 12572 14980
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 16666 15008 16672 15020
rect 16627 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 16850 15008 16856 15020
rect 16811 14980 16856 15008
rect 16850 14968 16856 14980
rect 16908 14968 16914 15020
rect 12544 14912 13400 14940
rect 12437 14903 12495 14909
rect 8159 14844 9444 14872
rect 9484 14875 9542 14881
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 9484 14841 9496 14875
rect 9530 14841 9542 14875
rect 9484 14835 9542 14841
rect 2639 14776 4844 14804
rect 2639 14773 2651 14776
rect 2593 14767 2651 14773
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 6454 14804 6460 14816
rect 4948 14776 6460 14804
rect 4948 14764 4954 14776
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 6604 14776 8033 14804
rect 6604 14764 6610 14776
rect 8021 14773 8033 14776
rect 8067 14804 8079 14807
rect 8846 14804 8852 14816
rect 8067 14776 8852 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 9508 14804 9536 14835
rect 9582 14832 9588 14884
rect 9640 14872 9646 14884
rect 12704 14875 12762 14881
rect 12704 14872 12716 14875
rect 9640 14844 12716 14872
rect 9640 14832 9646 14844
rect 12704 14841 12716 14844
rect 12750 14872 12762 14875
rect 13170 14872 13176 14884
rect 12750 14844 13176 14872
rect 12750 14841 12762 14844
rect 12704 14835 12762 14841
rect 13170 14832 13176 14844
rect 13228 14832 13234 14884
rect 13372 14872 13400 14912
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 13504 14912 15025 14940
rect 13504 14900 13510 14912
rect 15013 14909 15025 14912
rect 15059 14909 15071 14943
rect 16574 14940 16580 14952
rect 16535 14912 16580 14940
rect 15013 14903 15071 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 17494 14900 17500 14952
rect 17552 14940 17558 14952
rect 17862 14940 17868 14952
rect 17552 14912 17868 14940
rect 17552 14900 17558 14912
rect 17862 14900 17868 14912
rect 17920 14940 17926 14952
rect 18601 14943 18659 14949
rect 18601 14940 18613 14943
rect 17920 14912 18613 14940
rect 17920 14900 17926 14912
rect 18601 14909 18613 14912
rect 18647 14909 18659 14943
rect 18601 14903 18659 14909
rect 18868 14943 18926 14949
rect 18868 14909 18880 14943
rect 18914 14940 18926 14943
rect 19242 14940 19248 14952
rect 18914 14912 19248 14940
rect 18914 14909 18926 14912
rect 18868 14903 18926 14909
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 14458 14872 14464 14884
rect 13372 14844 14464 14872
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 14642 14832 14648 14884
rect 14700 14872 14706 14884
rect 15105 14875 15163 14881
rect 15105 14872 15117 14875
rect 14700 14844 15117 14872
rect 14700 14832 14706 14844
rect 15105 14841 15117 14844
rect 15151 14841 15163 14875
rect 15105 14835 15163 14841
rect 10870 14804 10876 14816
rect 9508 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 11790 14764 11796 14816
rect 11848 14804 11854 14816
rect 12069 14807 12127 14813
rect 12069 14804 12081 14807
rect 11848 14776 12081 14804
rect 11848 14764 11854 14776
rect 12069 14773 12081 14776
rect 12115 14804 12127 14807
rect 12342 14804 12348 14816
rect 12115 14776 12348 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 18690 14804 18696 14816
rect 12676 14776 18696 14804
rect 12676 14764 12682 14776
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 3053 14603 3111 14609
rect 3053 14569 3065 14603
rect 3099 14600 3111 14603
rect 4890 14600 4896 14612
rect 3099 14572 4896 14600
rect 3099 14569 3111 14572
rect 3053 14563 3111 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 5258 14600 5264 14612
rect 5092 14572 5264 14600
rect 5092 14541 5120 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7156 14572 7481 14600
rect 7156 14560 7162 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 7576 14572 7972 14600
rect 5068 14535 5126 14541
rect 5068 14501 5080 14535
rect 5114 14501 5126 14535
rect 5068 14495 5126 14501
rect 6454 14492 6460 14544
rect 6512 14532 6518 14544
rect 7576 14532 7604 14572
rect 6512 14504 7604 14532
rect 6512 14492 6518 14504
rect 7650 14492 7656 14544
rect 7708 14532 7714 14544
rect 7834 14532 7840 14544
rect 7708 14504 7840 14532
rect 7708 14492 7714 14504
rect 7834 14492 7840 14504
rect 7892 14492 7898 14544
rect 7944 14532 7972 14572
rect 8478 14560 8484 14612
rect 8536 14600 8542 14612
rect 8573 14603 8631 14609
rect 8573 14600 8585 14603
rect 8536 14572 8585 14600
rect 8536 14560 8542 14572
rect 8573 14569 8585 14572
rect 8619 14569 8631 14603
rect 8573 14563 8631 14569
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10502 14600 10508 14612
rect 10091 14572 10508 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 11609 14603 11667 14609
rect 11609 14569 11621 14603
rect 11655 14600 11667 14603
rect 14182 14600 14188 14612
rect 11655 14572 14188 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 15838 14600 15844 14612
rect 15344 14572 15844 14600
rect 15344 14560 15350 14572
rect 15838 14560 15844 14572
rect 15896 14600 15902 14612
rect 17589 14603 17647 14609
rect 17589 14600 17601 14603
rect 15896 14572 17601 14600
rect 15896 14560 15902 14572
rect 17589 14569 17601 14572
rect 17635 14569 17647 14603
rect 17589 14563 17647 14569
rect 9950 14532 9956 14544
rect 7944 14504 9956 14532
rect 9950 14492 9956 14504
rect 10008 14492 10014 14544
rect 10413 14535 10471 14541
rect 10413 14501 10425 14535
rect 10459 14532 10471 14535
rect 12066 14532 12072 14544
rect 10459 14504 12072 14532
rect 10459 14501 10471 14504
rect 10413 14495 10471 14501
rect 12066 14492 12072 14504
rect 12124 14492 12130 14544
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 13170 14532 13176 14544
rect 13044 14504 13176 14532
rect 13044 14492 13050 14504
rect 13170 14492 13176 14504
rect 13228 14492 13234 14544
rect 16022 14492 16028 14544
rect 16080 14532 16086 14544
rect 16390 14532 16396 14544
rect 16080 14504 16396 14532
rect 16080 14492 16086 14504
rect 16390 14492 16396 14504
rect 16448 14541 16454 14544
rect 16448 14535 16512 14541
rect 16448 14501 16466 14535
rect 16500 14501 16512 14535
rect 16448 14495 16512 14501
rect 16448 14492 16454 14495
rect 1762 14464 1768 14476
rect 1723 14436 1768 14464
rect 1762 14424 1768 14436
rect 1820 14424 1826 14476
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14464 2927 14467
rect 2915 14436 7236 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 4798 14396 4804 14408
rect 4759 14368 4804 14396
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 7208 14396 7236 14436
rect 7282 14424 7288 14476
rect 7340 14464 7346 14476
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 7340 14436 7389 14464
rect 7340 14424 7346 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 10318 14464 10324 14476
rect 7377 14427 7435 14433
rect 7484 14436 10324 14464
rect 7484 14396 7512 14436
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 10870 14464 10876 14476
rect 10796 14436 10876 14464
rect 7650 14396 7656 14408
rect 7208 14368 7512 14396
rect 7611 14368 7656 14396
rect 7650 14356 7656 14368
rect 7708 14356 7714 14408
rect 7742 14356 7748 14408
rect 7800 14396 7806 14408
rect 9858 14396 9864 14408
rect 7800 14368 9864 14396
rect 7800 14356 7806 14368
rect 9858 14356 9864 14368
rect 9916 14356 9922 14408
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10284 14368 10517 14396
rect 10284 14356 10290 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10689 14399 10747 14405
rect 10689 14365 10701 14399
rect 10735 14396 10747 14399
rect 10796 14396 10824 14436
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11940 14436 11989 14464
rect 11940 14424 11946 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12802 14424 12808 14476
rect 12860 14464 12866 14476
rect 13541 14467 13599 14473
rect 13541 14464 13553 14467
rect 12860 14436 13553 14464
rect 12860 14424 12866 14436
rect 13541 14433 13553 14436
rect 13587 14433 13599 14467
rect 13541 14427 13599 14433
rect 13633 14467 13691 14473
rect 13633 14433 13645 14467
rect 13679 14464 13691 14467
rect 13814 14464 13820 14476
rect 13679 14436 13820 14464
rect 13679 14433 13691 14436
rect 13633 14427 13691 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 14458 14424 14464 14476
rect 14516 14464 14522 14476
rect 14734 14464 14740 14476
rect 14516 14436 14740 14464
rect 14516 14424 14522 14436
rect 14734 14424 14740 14436
rect 14792 14464 14798 14476
rect 15105 14467 15163 14473
rect 15105 14464 15117 14467
rect 14792 14436 15117 14464
rect 14792 14424 14798 14436
rect 15105 14433 15117 14436
rect 15151 14433 15163 14467
rect 15105 14427 15163 14433
rect 15286 14424 15292 14476
rect 15344 14464 15350 14476
rect 16209 14467 16267 14473
rect 16209 14464 16221 14467
rect 15344 14436 16221 14464
rect 15344 14424 15350 14436
rect 16209 14433 16221 14436
rect 16255 14464 16267 14467
rect 17862 14464 17868 14476
rect 16255 14436 17868 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 19610 14464 19616 14476
rect 19571 14436 19616 14464
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 12066 14396 12072 14408
rect 10735 14368 10824 14396
rect 12027 14368 12072 14396
rect 10735 14365 10747 14368
rect 10689 14359 10747 14365
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12253 14399 12311 14405
rect 12253 14365 12265 14399
rect 12299 14396 12311 14399
rect 12894 14396 12900 14408
rect 12299 14368 12900 14396
rect 12299 14365 12311 14368
rect 12253 14359 12311 14365
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13504 14368 13737 14396
rect 13504 14356 13510 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 19702 14396 19708 14408
rect 19663 14368 19708 14396
rect 13725 14359 13783 14365
rect 19702 14356 19708 14368
rect 19760 14356 19766 14408
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14396 19947 14399
rect 20162 14396 20168 14408
rect 19935 14368 20168 14396
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 1949 14331 2007 14337
rect 1949 14297 1961 14331
rect 1995 14328 2007 14331
rect 10962 14328 10968 14340
rect 1995 14300 4844 14328
rect 1995 14297 2007 14300
rect 1949 14291 2007 14297
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 3694 14260 3700 14272
rect 2096 14232 3700 14260
rect 2096 14220 2102 14232
rect 3694 14220 3700 14232
rect 3752 14220 3758 14272
rect 4816 14260 4844 14300
rect 5736 14300 10968 14328
rect 5736 14260 5764 14300
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 11054 14288 11060 14340
rect 11112 14328 11118 14340
rect 11974 14328 11980 14340
rect 11112 14300 11980 14328
rect 11112 14288 11118 14300
rect 11974 14288 11980 14300
rect 12032 14288 12038 14340
rect 12158 14288 12164 14340
rect 12216 14328 12222 14340
rect 13173 14331 13231 14337
rect 13173 14328 13185 14331
rect 12216 14300 13185 14328
rect 12216 14288 12222 14300
rect 13173 14297 13185 14300
rect 13219 14297 13231 14331
rect 13173 14291 13231 14297
rect 14921 14331 14979 14337
rect 14921 14297 14933 14331
rect 14967 14328 14979 14331
rect 15286 14328 15292 14340
rect 14967 14300 15292 14328
rect 14967 14297 14979 14300
rect 14921 14291 14979 14297
rect 15286 14288 15292 14300
rect 15344 14288 15350 14340
rect 6178 14260 6184 14272
rect 4816 14232 5764 14260
rect 6139 14232 6184 14260
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 7009 14263 7067 14269
rect 7009 14229 7021 14263
rect 7055 14260 7067 14263
rect 9674 14260 9680 14272
rect 7055 14232 9680 14260
rect 7055 14229 7067 14232
rect 7009 14223 7067 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14260 10011 14263
rect 10226 14260 10232 14272
rect 9999 14232 10232 14260
rect 9999 14229 10011 14232
rect 9953 14223 10011 14229
rect 10226 14220 10232 14232
rect 10284 14220 10290 14272
rect 10318 14220 10324 14272
rect 10376 14260 10382 14272
rect 17126 14260 17132 14272
rect 10376 14232 17132 14260
rect 10376 14220 10382 14232
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 19245 14263 19303 14269
rect 19245 14260 19257 14263
rect 18196 14232 19257 14260
rect 18196 14220 18202 14232
rect 19245 14229 19257 14232
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 9858 14056 9864 14068
rect 3752 14028 7972 14056
rect 3752 14016 3758 14028
rect 1854 13988 1860 14000
rect 1815 13960 1860 13988
rect 1854 13948 1860 13960
rect 1912 13948 1918 14000
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4157 13991 4215 13997
rect 4157 13988 4169 13991
rect 4120 13960 4169 13988
rect 4120 13948 4126 13960
rect 4157 13957 4169 13960
rect 4203 13957 4215 13991
rect 7282 13988 7288 14000
rect 7243 13960 7288 13988
rect 4157 13951 4215 13957
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 4448 13892 5549 13920
rect 1670 13852 1676 13864
rect 1631 13824 1676 13852
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2740 13824 2789 13852
rect 2740 13812 2746 13824
rect 2777 13821 2789 13824
rect 2823 13852 2835 13855
rect 2866 13852 2872 13864
rect 2823 13824 2872 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 3044 13787 3102 13793
rect 3044 13753 3056 13787
rect 3090 13784 3102 13787
rect 3878 13784 3884 13796
rect 3090 13756 3884 13784
rect 3090 13753 3102 13756
rect 3044 13747 3102 13753
rect 3878 13744 3884 13756
rect 3936 13784 3942 13796
rect 4448 13784 4476 13892
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 6236 13892 7849 13920
rect 6236 13880 6242 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7944 13920 7972 14028
rect 9784 14028 9864 14056
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8260 13960 9628 13988
rect 8260 13948 8266 13960
rect 9030 13920 9036 13932
rect 7944 13892 9036 13920
rect 7837 13883 7895 13889
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 6822 13852 6828 13864
rect 5491 13824 6828 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 6972 13824 7757 13852
rect 6972 13812 6978 13824
rect 7745 13821 7757 13824
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13821 9459 13855
rect 9600 13852 9628 13960
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9784 13920 9812 14028
rect 9858 14016 9864 14028
rect 9916 14016 9922 14068
rect 10781 14059 10839 14065
rect 10781 14025 10793 14059
rect 10827 14056 10839 14059
rect 12066 14056 12072 14068
rect 10827 14028 12072 14056
rect 10827 14025 10839 14028
rect 10781 14019 10839 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 18782 14056 18788 14068
rect 14415 14028 18788 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 20070 14056 20076 14068
rect 19843 14028 20076 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 12894 13948 12900 14000
rect 12952 13988 12958 14000
rect 12952 13960 14596 13988
rect 12952 13948 12958 13960
rect 14568 13932 14596 13960
rect 16390 13948 16396 14000
rect 16448 13988 16454 14000
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 16448 13960 16681 13988
rect 16448 13948 16454 13960
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 16669 13951 16727 13957
rect 9723 13892 9812 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 10686 13880 10692 13932
rect 10744 13920 10750 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 10744 13892 11345 13920
rect 10744 13880 10750 13892
rect 11333 13889 11345 13892
rect 11379 13889 11391 13923
rect 11333 13883 11391 13889
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13920 13231 13923
rect 13722 13920 13728 13932
rect 13219 13892 13728 13920
rect 13219 13889 13231 13892
rect 13173 13883 13231 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 14550 13880 14556 13932
rect 14608 13920 14614 13932
rect 15194 13920 15200 13932
rect 14608 13892 15200 13920
rect 14608 13880 14614 13892
rect 15194 13880 15200 13892
rect 15252 13920 15258 13932
rect 18782 13920 18788 13932
rect 15252 13892 15424 13920
rect 18743 13892 18788 13920
rect 15252 13880 15258 13892
rect 9600 13824 9720 13852
rect 9401 13815 9459 13821
rect 3936 13756 4476 13784
rect 3936 13744 3942 13756
rect 4798 13744 4804 13796
rect 4856 13784 4862 13796
rect 5353 13787 5411 13793
rect 5353 13784 5365 13787
rect 4856 13756 5365 13784
rect 4856 13744 4862 13756
rect 5353 13753 5365 13756
rect 5399 13753 5411 13787
rect 5353 13747 5411 13753
rect 7653 13787 7711 13793
rect 7653 13753 7665 13787
rect 7699 13784 7711 13787
rect 7834 13784 7840 13796
rect 7699 13756 7840 13784
rect 7699 13753 7711 13756
rect 7653 13747 7711 13753
rect 7834 13744 7840 13756
rect 7892 13744 7898 13796
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 9407 13784 9435 13815
rect 8904 13756 9435 13784
rect 9493 13787 9551 13793
rect 8904 13744 8910 13756
rect 9493 13753 9505 13787
rect 9539 13784 9551 13787
rect 9582 13784 9588 13796
rect 9539 13756 9588 13784
rect 9539 13753 9551 13756
rect 9493 13747 9551 13753
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 9692 13784 9720 13824
rect 10410 13812 10416 13864
rect 10468 13852 10474 13864
rect 11238 13852 11244 13864
rect 10468 13824 11244 13852
rect 10468 13812 10474 13824
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 11698 13812 11704 13864
rect 11756 13852 11762 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 11756 13824 12449 13852
rect 11756 13812 11762 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12986 13852 12992 13864
rect 12947 13824 12992 13852
rect 12437 13815 12495 13821
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 14185 13855 14243 13861
rect 14185 13821 14197 13855
rect 14231 13852 14243 13855
rect 14458 13852 14464 13864
rect 14231 13824 14464 13852
rect 14231 13821 14243 13824
rect 14185 13815 14243 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 15286 13852 15292 13864
rect 15247 13824 15292 13852
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15396 13852 15424 13892
rect 18782 13880 18788 13892
rect 18840 13880 18846 13932
rect 19242 13880 19248 13932
rect 19300 13920 19306 13932
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 19300 13892 20361 13920
rect 19300 13880 19306 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 15545 13855 15603 13861
rect 15545 13852 15557 13855
rect 15396 13824 15557 13852
rect 15545 13821 15557 13824
rect 15591 13821 15603 13855
rect 15545 13815 15603 13821
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 18693 13855 18751 13861
rect 18693 13852 18705 13855
rect 16356 13824 18705 13852
rect 16356 13812 16362 13824
rect 18693 13821 18705 13824
rect 18739 13821 18751 13855
rect 18693 13815 18751 13821
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19978 13852 19984 13864
rect 19576 13824 19984 13852
rect 19576 13812 19582 13824
rect 19978 13812 19984 13824
rect 20036 13852 20042 13864
rect 20257 13855 20315 13861
rect 20257 13852 20269 13855
rect 20036 13824 20269 13852
rect 20036 13812 20042 13824
rect 20257 13821 20269 13824
rect 20303 13821 20315 13855
rect 20257 13815 20315 13821
rect 18601 13787 18659 13793
rect 18601 13784 18613 13787
rect 9692 13756 18613 13784
rect 18601 13753 18613 13756
rect 18647 13753 18659 13787
rect 18601 13747 18659 13753
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 4985 13719 5043 13725
rect 4985 13716 4997 13719
rect 3844 13688 4997 13716
rect 3844 13676 3850 13688
rect 4985 13685 4997 13688
rect 5031 13685 5043 13719
rect 4985 13679 5043 13685
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 6546 13716 6552 13728
rect 5592 13688 6552 13716
rect 5592 13676 5598 13688
rect 6546 13676 6552 13688
rect 6604 13716 6610 13728
rect 8754 13716 8760 13728
rect 6604 13688 8760 13716
rect 6604 13676 6610 13688
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 9033 13719 9091 13725
rect 9033 13685 9045 13719
rect 9079 13716 9091 13719
rect 9306 13716 9312 13728
rect 9079 13688 9312 13716
rect 9079 13685 9091 13688
rect 9033 13679 9091 13685
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10870 13716 10876 13728
rect 10560 13688 10876 13716
rect 10560 13676 10566 13688
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11149 13719 11207 13725
rect 11149 13685 11161 13719
rect 11195 13716 11207 13719
rect 11330 13716 11336 13728
rect 11195 13688 11336 13716
rect 11195 13685 11207 13688
rect 11149 13679 11207 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 12437 13719 12495 13725
rect 12437 13685 12449 13719
rect 12483 13716 12495 13719
rect 12529 13719 12587 13725
rect 12529 13716 12541 13719
rect 12483 13688 12541 13716
rect 12483 13685 12495 13688
rect 12437 13679 12495 13685
rect 12529 13685 12541 13688
rect 12575 13685 12587 13719
rect 12894 13716 12900 13728
rect 12855 13688 12900 13716
rect 12529 13679 12587 13685
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 16298 13716 16304 13728
rect 15712 13688 16304 13716
rect 15712 13676 15718 13688
rect 16298 13676 16304 13688
rect 16356 13676 16362 13728
rect 18230 13716 18236 13728
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 19242 13676 19248 13728
rect 19300 13716 19306 13728
rect 20165 13719 20223 13725
rect 20165 13716 20177 13719
rect 19300 13688 20177 13716
rect 19300 13676 19306 13688
rect 20165 13685 20177 13688
rect 20211 13685 20223 13719
rect 20165 13679 20223 13685
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 1394 13512 1400 13524
rect 1355 13484 1400 13512
rect 1394 13472 1400 13484
rect 1452 13472 1458 13524
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 2866 13512 2872 13524
rect 2823 13484 2872 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 2866 13472 2872 13484
rect 2924 13512 2930 13524
rect 3050 13512 3056 13524
rect 2924 13484 3056 13512
rect 2924 13472 2930 13484
rect 3050 13472 3056 13484
rect 3108 13472 3114 13524
rect 8294 13512 8300 13524
rect 3988 13484 8300 13512
rect 2498 13404 2504 13456
rect 2556 13444 2562 13456
rect 3988 13444 4016 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 8478 13512 8484 13524
rect 8435 13484 8484 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 9677 13515 9735 13521
rect 9677 13481 9689 13515
rect 9723 13481 9735 13515
rect 9677 13475 9735 13481
rect 6454 13444 6460 13456
rect 2556 13416 4016 13444
rect 4080 13416 6460 13444
rect 2556 13404 2562 13416
rect 1762 13336 1768 13388
rect 1820 13376 1826 13388
rect 4080 13376 4108 13416
rect 6454 13404 6460 13416
rect 6512 13444 6518 13456
rect 6512 13416 7880 13444
rect 6512 13404 6518 13416
rect 1820 13348 4108 13376
rect 4157 13379 4215 13385
rect 1820 13336 1826 13348
rect 4157 13345 4169 13379
rect 4203 13376 4215 13379
rect 4246 13376 4252 13388
rect 4203 13348 4252 13376
rect 4203 13345 4215 13348
rect 4157 13339 4215 13345
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 5534 13376 5540 13388
rect 5491 13348 5540 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 5712 13379 5770 13385
rect 5712 13345 5724 13379
rect 5758 13376 5770 13379
rect 7742 13376 7748 13388
rect 5758 13348 7748 13376
rect 5758 13345 5770 13348
rect 5712 13339 5770 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 2774 13268 2780 13320
rect 2832 13308 2838 13320
rect 2869 13311 2927 13317
rect 2869 13308 2881 13311
rect 2832 13280 2881 13308
rect 2832 13268 2838 13280
rect 2869 13277 2881 13280
rect 2915 13277 2927 13311
rect 3050 13308 3056 13320
rect 3011 13280 3056 13308
rect 2869 13271 2927 13277
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13308 4491 13311
rect 5258 13308 5264 13320
rect 4479 13280 5264 13308
rect 4479 13277 4491 13280
rect 4433 13271 4491 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 7466 13308 7472 13320
rect 6840 13280 7472 13308
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 5166 13172 5172 13184
rect 2455 13144 5172 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5442 13132 5448 13184
rect 5500 13172 5506 13184
rect 6840 13181 6868 13280
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 7745 13243 7803 13249
rect 7745 13240 7757 13243
rect 7064 13212 7757 13240
rect 7064 13200 7070 13212
rect 7745 13209 7757 13212
rect 7791 13209 7803 13243
rect 7852 13240 7880 13416
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 9692 13444 9720 13475
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13481 10103 13515
rect 10045 13475 10103 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10318 13512 10324 13524
rect 10183 13484 10324 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10318 13472 10324 13484
rect 10376 13472 10382 13524
rect 11517 13515 11575 13521
rect 11517 13481 11529 13515
rect 11563 13512 11575 13515
rect 12618 13512 12624 13524
rect 11563 13484 12624 13512
rect 11563 13481 11575 13484
rect 11517 13475 11575 13481
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13481 13875 13515
rect 13817 13475 13875 13481
rect 14645 13515 14703 13521
rect 14645 13481 14657 13515
rect 14691 13512 14703 13515
rect 14734 13512 14740 13524
rect 14691 13484 14740 13512
rect 14691 13481 14703 13484
rect 14645 13475 14703 13481
rect 13630 13444 13636 13456
rect 9456 13416 9720 13444
rect 10704 13416 13636 13444
rect 9456 13404 9462 13416
rect 10704 13388 10732 13416
rect 13630 13404 13636 13416
rect 13688 13444 13694 13456
rect 13832 13444 13860 13475
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 18049 13515 18107 13521
rect 18049 13481 18061 13515
rect 18095 13512 18107 13515
rect 18230 13512 18236 13524
rect 18095 13484 18236 13512
rect 18095 13481 18107 13484
rect 18049 13475 18107 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19245 13515 19303 13521
rect 19245 13481 19257 13515
rect 19291 13512 19303 13515
rect 19702 13512 19708 13524
rect 19291 13484 19708 13512
rect 19291 13481 19303 13484
rect 19245 13475 19303 13481
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 13688 13416 13860 13444
rect 15749 13447 15807 13453
rect 13688 13404 13694 13416
rect 15749 13413 15761 13447
rect 15795 13444 15807 13447
rect 15838 13444 15844 13456
rect 15795 13416 15844 13444
rect 15795 13413 15807 13416
rect 15749 13407 15807 13413
rect 15838 13404 15844 13416
rect 15896 13404 15902 13456
rect 16022 13404 16028 13456
rect 16080 13444 16086 13456
rect 19334 13444 19340 13456
rect 16080 13416 19340 13444
rect 16080 13404 16086 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13376 7987 13379
rect 9030 13376 9036 13388
rect 7975 13348 9036 13376
rect 7975 13345 7987 13348
rect 7929 13339 7987 13345
rect 9030 13336 9036 13348
rect 9088 13336 9094 13388
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 10686 13376 10692 13388
rect 9640 13348 10692 13376
rect 9640 13336 9646 13348
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11790 13376 11796 13388
rect 11379 13348 11796 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12693 13379 12751 13385
rect 12693 13376 12705 13379
rect 12032 13348 12705 13376
rect 12032 13336 12038 13348
rect 12693 13345 12705 13348
rect 12739 13345 12751 13379
rect 12693 13339 12751 13345
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 14829 13379 14887 13385
rect 14829 13376 14841 13379
rect 14792 13348 14841 13376
rect 14792 13336 14798 13348
rect 14829 13345 14841 13348
rect 14875 13345 14887 13379
rect 15654 13376 15660 13388
rect 15615 13348 15660 13376
rect 14829 13339 14887 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 19518 13376 19524 13388
rect 16632 13348 19524 13376
rect 16632 13336 16638 13348
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 20530 13376 20536 13388
rect 19659 13348 20536 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13277 8539 13311
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8481 13271 8539 13277
rect 8496 13240 8524 13271
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9858 13308 9864 13320
rect 9732 13280 9864 13308
rect 9732 13268 9738 13280
rect 9858 13268 9864 13280
rect 9916 13308 9922 13320
rect 10229 13311 10287 13317
rect 10229 13308 10241 13311
rect 9916 13280 10241 13308
rect 9916 13268 9922 13280
rect 10229 13277 10241 13280
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12400 13280 12449 13308
rect 12400 13268 12406 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 15841 13311 15899 13317
rect 15841 13277 15853 13311
rect 15887 13277 15899 13311
rect 15841 13271 15899 13277
rect 9122 13240 9128 13252
rect 7852 13212 8156 13240
rect 8496 13212 9128 13240
rect 7745 13203 7803 13209
rect 6825 13175 6883 13181
rect 6825 13172 6837 13175
rect 5500 13144 6837 13172
rect 5500 13132 5506 13144
rect 6825 13141 6837 13144
rect 6871 13141 6883 13175
rect 8018 13172 8024 13184
rect 7979 13144 8024 13172
rect 6825 13135 6883 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8128 13172 8156 13212
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 13446 13200 13452 13252
rect 13504 13240 13510 13252
rect 15856 13240 15884 13271
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 18141 13311 18199 13317
rect 18141 13308 18153 13311
rect 16448 13280 18153 13308
rect 16448 13268 16454 13280
rect 18141 13277 18153 13280
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 18325 13311 18383 13317
rect 18325 13277 18337 13311
rect 18371 13308 18383 13311
rect 19334 13308 19340 13320
rect 18371 13280 19340 13308
rect 18371 13277 18383 13280
rect 18325 13271 18383 13277
rect 19334 13268 19340 13280
rect 19392 13268 19398 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19484 13280 19717 13308
rect 19484 13268 19490 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19886 13308 19892 13320
rect 19847 13280 19892 13308
rect 19705 13271 19763 13277
rect 19886 13268 19892 13280
rect 19944 13268 19950 13320
rect 13504 13212 15884 13240
rect 13504 13200 13510 13212
rect 16022 13200 16028 13252
rect 16080 13240 16086 13252
rect 17586 13240 17592 13252
rect 16080 13212 17592 13240
rect 16080 13200 16086 13212
rect 17586 13200 17592 13212
rect 17644 13200 17650 13252
rect 12158 13172 12164 13184
rect 8128 13144 12164 13172
rect 12158 13132 12164 13144
rect 12216 13132 12222 13184
rect 12618 13132 12624 13184
rect 12676 13172 12682 13184
rect 14090 13172 14096 13184
rect 12676 13144 14096 13172
rect 12676 13132 12682 13144
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 15194 13132 15200 13184
rect 15252 13172 15258 13184
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 15252 13144 15301 13172
rect 15252 13132 15258 13144
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 17494 13132 17500 13184
rect 17552 13172 17558 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17552 13144 17693 13172
rect 17552 13132 17558 13144
rect 17681 13141 17693 13144
rect 17727 13141 17739 13175
rect 17681 13135 17739 13141
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 6822 12968 6828 12980
rect 6783 12940 6828 12968
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7282 12968 7288 12980
rect 7156 12940 7288 12968
rect 7156 12928 7162 12940
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 12434 12968 12440 12980
rect 8076 12940 12440 12968
rect 8076 12928 8082 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12713 12971 12771 12977
rect 12713 12937 12725 12971
rect 12759 12968 12771 12971
rect 15013 12971 15071 12977
rect 12759 12940 14872 12968
rect 12759 12937 12771 12940
rect 12713 12931 12771 12937
rect 3878 12900 3884 12912
rect 3839 12872 3884 12900
rect 3878 12860 3884 12872
rect 3936 12900 3942 12912
rect 3936 12872 5304 12900
rect 3936 12860 3942 12872
rect 5166 12832 5172 12844
rect 5127 12804 5172 12832
rect 5166 12792 5172 12804
rect 5224 12792 5230 12844
rect 5276 12841 5304 12872
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 5718 12900 5724 12912
rect 5592 12872 5724 12900
rect 5592 12860 5598 12872
rect 5718 12860 5724 12872
rect 5776 12860 5782 12912
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 8389 12903 8447 12909
rect 8389 12900 8401 12903
rect 6788 12872 8401 12900
rect 6788 12860 6794 12872
rect 8389 12869 8401 12872
rect 8435 12869 8447 12903
rect 8389 12863 8447 12869
rect 10520 12872 10732 12900
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12801 5319 12835
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 5261 12795 5319 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 7800 12804 8953 12832
rect 7800 12792 7806 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 9306 12792 9312 12844
rect 9364 12832 9370 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 9364 12804 10425 12832
rect 9364 12792 9370 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 2768 12767 2826 12773
rect 2768 12733 2780 12767
rect 2814 12764 2826 12767
rect 3050 12764 3056 12776
rect 2814 12736 3056 12764
rect 2814 12733 2826 12736
rect 2768 12727 2826 12733
rect 2516 12696 2544 12727
rect 3050 12724 3056 12736
rect 3108 12764 3114 12776
rect 4522 12764 4528 12776
rect 3108 12736 4528 12764
rect 3108 12724 3114 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 6362 12724 6368 12776
rect 6420 12764 6426 12776
rect 10520 12764 10548 12872
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10704 12832 10732 12872
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 11698 12900 11704 12912
rect 11204 12872 11704 12900
rect 11204 12860 11210 12872
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 12342 12900 12348 12912
rect 12216 12872 12348 12900
rect 12216 12860 12222 12872
rect 12342 12860 12348 12872
rect 12400 12900 12406 12912
rect 14844 12900 14872 12940
rect 15013 12937 15025 12971
rect 15059 12968 15071 12971
rect 15102 12968 15108 12980
rect 15059 12940 15108 12968
rect 15059 12937 15071 12940
rect 15013 12931 15071 12937
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 19150 12968 19156 12980
rect 17604 12940 19156 12968
rect 17604 12900 17632 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 19334 12928 19340 12980
rect 19392 12968 19398 12980
rect 19702 12968 19708 12980
rect 19392 12940 19708 12968
rect 19392 12928 19398 12940
rect 19702 12928 19708 12940
rect 19760 12968 19766 12980
rect 20349 12971 20407 12977
rect 20349 12968 20361 12971
rect 19760 12940 20361 12968
rect 19760 12928 19766 12940
rect 20349 12937 20361 12940
rect 20395 12937 20407 12971
rect 20349 12931 20407 12937
rect 12400 12872 13676 12900
rect 14844 12872 17632 12900
rect 12400 12860 12406 12872
rect 12894 12832 12900 12844
rect 10704 12804 12900 12832
rect 10597 12795 10655 12801
rect 6420 12736 10548 12764
rect 6420 12724 6426 12736
rect 2682 12696 2688 12708
rect 2516 12668 2688 12696
rect 2682 12656 2688 12668
rect 2740 12656 2746 12708
rect 3234 12656 3240 12708
rect 3292 12696 3298 12708
rect 3602 12696 3608 12708
rect 3292 12668 3608 12696
rect 3292 12656 3298 12668
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 8110 12696 8116 12708
rect 3936 12668 8116 12696
rect 3936 12656 3942 12668
rect 8110 12656 8116 12668
rect 8168 12656 8174 12708
rect 8202 12656 8208 12708
rect 8260 12696 8266 12708
rect 9490 12696 9496 12708
rect 8260 12668 9496 12696
rect 8260 12656 8266 12668
rect 9490 12656 9496 12668
rect 9548 12696 9554 12708
rect 9548 12668 10456 12696
rect 9548 12656 9554 12668
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4709 12631 4767 12637
rect 4709 12628 4721 12631
rect 4212 12600 4721 12628
rect 4212 12588 4218 12600
rect 4709 12597 4721 12600
rect 4755 12597 4767 12631
rect 5074 12628 5080 12640
rect 5035 12600 5080 12628
rect 4709 12591 4767 12597
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7156 12600 7205 12628
rect 7156 12588 7162 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 7282 12588 7288 12640
rect 7340 12628 7346 12640
rect 7466 12628 7472 12640
rect 7340 12600 7472 12628
rect 7340 12588 7346 12600
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8754 12628 8760 12640
rect 8715 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 8849 12631 8907 12637
rect 8849 12597 8861 12631
rect 8895 12628 8907 12631
rect 9953 12631 10011 12637
rect 9953 12628 9965 12631
rect 8895 12600 9965 12628
rect 8895 12597 8907 12600
rect 8849 12591 8907 12597
rect 9953 12597 9965 12600
rect 9999 12597 10011 12631
rect 10318 12628 10324 12640
rect 10279 12600 10324 12628
rect 9953 12591 10011 12597
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10428 12628 10456 12668
rect 10612 12628 10640 12795
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13538 12832 13544 12844
rect 13412 12804 13544 12832
rect 13412 12792 13418 12804
rect 13538 12792 13544 12804
rect 13596 12792 13602 12844
rect 13648 12841 13676 12872
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 17037 12835 17095 12841
rect 13633 12795 13691 12801
rect 16592 12804 16988 12832
rect 12529 12767 12587 12773
rect 12529 12733 12541 12767
rect 12575 12764 12587 12767
rect 16592 12764 16620 12804
rect 16758 12764 16764 12776
rect 12575 12736 16620 12764
rect 16719 12736 16764 12764
rect 12575 12733 12587 12736
rect 12529 12727 12587 12733
rect 16758 12724 16764 12736
rect 16816 12724 16822 12776
rect 16960 12764 16988 12804
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 18782 12832 18788 12844
rect 17083 12804 18788 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 18782 12792 18788 12804
rect 18840 12832 18846 12844
rect 18840 12804 19104 12832
rect 18840 12792 18846 12804
rect 17310 12764 17316 12776
rect 16960 12736 17316 12764
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 17920 12736 18981 12764
rect 17920 12724 17926 12736
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 19076 12764 19104 12804
rect 19242 12773 19248 12776
rect 19225 12767 19248 12773
rect 19225 12764 19237 12767
rect 19076 12736 19237 12764
rect 18969 12727 19027 12733
rect 19225 12733 19237 12736
rect 19300 12764 19306 12776
rect 19300 12736 19373 12764
rect 19225 12727 19248 12733
rect 19242 12724 19248 12727
rect 19300 12724 19306 12736
rect 12894 12656 12900 12708
rect 12952 12696 12958 12708
rect 13262 12696 13268 12708
rect 12952 12668 13268 12696
rect 12952 12656 12958 12668
rect 13262 12656 13268 12668
rect 13320 12656 13326 12708
rect 13630 12656 13636 12708
rect 13688 12696 13694 12708
rect 13878 12699 13936 12705
rect 13878 12696 13890 12699
rect 13688 12668 13890 12696
rect 13688 12656 13694 12668
rect 13878 12665 13890 12668
rect 13924 12665 13936 12699
rect 13878 12659 13936 12665
rect 15562 12656 15568 12708
rect 15620 12696 15626 12708
rect 16114 12696 16120 12708
rect 15620 12668 16120 12696
rect 15620 12656 15626 12668
rect 16114 12656 16120 12668
rect 16172 12696 16178 12708
rect 18690 12696 18696 12708
rect 16172 12668 18696 12696
rect 16172 12656 16178 12668
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 10428 12600 10640 12628
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12526 12628 12532 12640
rect 11848 12600 12532 12628
rect 11848 12588 11854 12600
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 15286 12588 15292 12640
rect 15344 12628 15350 12640
rect 16853 12631 16911 12637
rect 16853 12628 16865 12631
rect 15344 12600 16865 12628
rect 15344 12588 15350 12600
rect 16853 12597 16865 12600
rect 16899 12597 16911 12631
rect 16853 12591 16911 12597
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17954 12628 17960 12640
rect 17460 12600 17960 12628
rect 17460 12588 17466 12600
rect 17954 12588 17960 12600
rect 18012 12588 18018 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4798 12424 4804 12436
rect 4295 12396 4804 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5442 12384 5448 12436
rect 5500 12424 5506 12436
rect 7650 12424 7656 12436
rect 5500 12396 7656 12424
rect 5500 12384 5506 12396
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 7800 12396 8125 12424
rect 7800 12384 7806 12396
rect 8113 12393 8125 12396
rect 8159 12393 8171 12427
rect 8113 12387 8171 12393
rect 10502 12384 10508 12436
rect 10560 12424 10566 12436
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 10560 12396 13645 12424
rect 10560 12384 10566 12396
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 14182 12384 14188 12436
rect 14240 12424 14246 12436
rect 15194 12424 15200 12436
rect 14240 12396 15200 12424
rect 14240 12384 14246 12396
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 15378 12424 15384 12436
rect 15335 12396 15384 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 18046 12424 18052 12436
rect 16715 12396 18052 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 4617 12359 4675 12365
rect 4617 12356 4629 12359
rect 1903 12328 4629 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 4617 12325 4629 12328
rect 4663 12325 4675 12359
rect 4617 12319 4675 12325
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 9953 12359 10011 12365
rect 4764 12328 8340 12356
rect 4764 12316 4770 12328
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 5442 12288 5448 12300
rect 2915 12260 5448 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 5442 12248 5448 12260
rect 5500 12248 5506 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6733 12291 6791 12297
rect 6733 12288 6745 12291
rect 5776 12260 6745 12288
rect 5776 12248 5782 12260
rect 6733 12257 6745 12260
rect 6779 12288 6791 12291
rect 6822 12288 6828 12300
rect 6779 12260 6828 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7000 12291 7058 12297
rect 7000 12257 7012 12291
rect 7046 12288 7058 12291
rect 8202 12288 8208 12300
rect 7046 12260 8208 12288
rect 7046 12257 7058 12260
rect 7000 12251 7058 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 8312 12220 8340 12328
rect 9953 12325 9965 12359
rect 9999 12356 10011 12359
rect 12158 12356 12164 12368
rect 9999 12328 10916 12356
rect 9999 12325 10011 12328
rect 9953 12319 10011 12325
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 8938 12288 8944 12300
rect 8720 12260 8944 12288
rect 8720 12248 8726 12260
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9122 12288 9128 12300
rect 9083 12260 9128 12288
rect 9122 12248 9128 12260
rect 9180 12248 9186 12300
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 9858 12288 9864 12300
rect 9723 12260 9864 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10686 12220 10692 12232
rect 8312 12192 10692 12220
rect 4801 12183 4859 12189
rect 3050 12152 3056 12164
rect 3011 12124 3056 12152
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 4522 12112 4528 12164
rect 4580 12152 4586 12164
rect 4816 12152 4844 12183
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10888 12220 10916 12328
rect 10980 12328 12164 12356
rect 10980 12297 11008 12328
rect 12158 12316 12164 12328
rect 12216 12316 12222 12368
rect 13722 12356 13728 12368
rect 12268 12328 13728 12356
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11232 12291 11290 12297
rect 11232 12257 11244 12291
rect 11278 12288 11290 12291
rect 12268 12288 12296 12328
rect 13722 12316 13728 12328
rect 13780 12316 13786 12368
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14366 12356 14372 12368
rect 13872 12328 14372 12356
rect 13872 12316 13878 12328
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 14642 12316 14648 12368
rect 14700 12356 14706 12368
rect 16316 12356 16344 12387
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 19242 12424 19248 12436
rect 19203 12396 19248 12424
rect 19242 12384 19248 12396
rect 19300 12384 19306 12436
rect 19426 12356 19432 12368
rect 14700 12328 15056 12356
rect 16316 12328 19432 12356
rect 14700 12316 14706 12328
rect 11278 12260 12296 12288
rect 11278 12257 11290 12260
rect 11232 12251 11290 12257
rect 12176 12232 12204 12260
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 13541 12291 13599 12297
rect 13541 12288 13553 12291
rect 13504 12260 13553 12288
rect 13504 12248 13510 12260
rect 13541 12257 13553 12260
rect 13587 12257 13599 12291
rect 13541 12251 13599 12257
rect 10888 12192 11008 12220
rect 5534 12152 5540 12164
rect 4580 12124 5540 12152
rect 4580 12112 4586 12124
rect 5534 12112 5540 12124
rect 5592 12112 5598 12164
rect 7742 12112 7748 12164
rect 7800 12152 7806 12164
rect 9858 12152 9864 12164
rect 7800 12124 9864 12152
rect 7800 12112 7806 12124
rect 9858 12112 9864 12124
rect 9916 12152 9922 12164
rect 10042 12152 10048 12164
rect 9916 12124 10048 12152
rect 9916 12112 9922 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 8662 12084 8668 12096
rect 5224 12056 8668 12084
rect 5224 12044 5230 12056
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9030 12084 9036 12096
rect 8987 12056 9036 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 10980 12084 11008 12192
rect 12158 12180 12164 12232
rect 12216 12180 12222 12232
rect 12618 12180 12624 12232
rect 12676 12220 12682 12232
rect 13740 12229 13768 12316
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 15028 12288 15056 12328
rect 19426 12316 19432 12328
rect 19484 12316 19490 12368
rect 17126 12288 17132 12300
rect 15028 12260 17132 12288
rect 14921 12251 14979 12257
rect 13725 12223 13783 12229
rect 12676 12192 13676 12220
rect 12676 12180 12682 12192
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12345 12155 12403 12161
rect 12345 12152 12357 12155
rect 12032 12124 12357 12152
rect 12032 12112 12038 12124
rect 12345 12121 12357 12124
rect 12391 12121 12403 12155
rect 12345 12115 12403 12121
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 13173 12155 13231 12161
rect 13173 12152 13185 12155
rect 12584 12124 13185 12152
rect 12584 12112 12590 12124
rect 13173 12121 13185 12124
rect 13219 12121 13231 12155
rect 13648 12152 13676 12192
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 14936 12152 14964 12251
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17862 12288 17868 12300
rect 17823 12260 17868 12288
rect 17862 12248 17868 12260
rect 17920 12248 17926 12300
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 18121 12291 18179 12297
rect 18121 12288 18133 12291
rect 18012 12260 18133 12288
rect 18012 12248 18018 12260
rect 18121 12257 18133 12260
rect 18167 12257 18179 12291
rect 18121 12251 18179 12257
rect 16574 12180 16580 12232
rect 16632 12220 16638 12232
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16632 12192 16773 12220
rect 16632 12180 16638 12192
rect 16761 12189 16773 12192
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 13648 12124 14964 12152
rect 13173 12115 13231 12121
rect 14274 12084 14280 12096
rect 10980 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 14734 12084 14740 12096
rect 14695 12056 14740 12084
rect 14734 12044 14740 12056
rect 14792 12044 14798 12096
rect 16960 12084 16988 12183
rect 18966 12112 18972 12164
rect 19024 12152 19030 12164
rect 20346 12152 20352 12164
rect 19024 12124 20352 12152
rect 19024 12112 19030 12124
rect 20346 12112 20352 12124
rect 20404 12112 20410 12164
rect 19794 12084 19800 12096
rect 16960 12056 19800 12084
rect 19794 12044 19800 12056
rect 19852 12084 19858 12096
rect 20622 12084 20628 12096
rect 19852 12056 20628 12084
rect 19852 12044 19858 12056
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 3513 11883 3571 11889
rect 3513 11849 3525 11883
rect 3559 11880 3571 11883
rect 4246 11880 4252 11892
rect 3559 11852 4252 11880
rect 3559 11849 3571 11852
rect 3513 11843 3571 11849
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5074 11880 5080 11892
rect 5035 11852 5080 11880
rect 5074 11840 5080 11852
rect 5132 11840 5138 11892
rect 8202 11880 8208 11892
rect 5552 11852 7788 11880
rect 8163 11852 8208 11880
rect 5552 11812 5580 11852
rect 1504 11784 5580 11812
rect 7760 11812 7788 11852
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8812 11852 9045 11880
rect 8812 11840 8818 11852
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 9033 11843 9091 11849
rect 9398 11840 9404 11892
rect 9456 11880 9462 11892
rect 9456 11852 10272 11880
rect 9456 11840 9462 11852
rect 8386 11812 8392 11824
rect 7760 11784 8392 11812
rect 1504 11753 1532 11784
rect 8386 11772 8392 11784
rect 8444 11772 8450 11824
rect 10042 11812 10048 11824
rect 8496 11784 10048 11812
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11744 2559 11747
rect 2958 11744 2964 11756
rect 2547 11716 2964 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 4062 11744 4068 11756
rect 4023 11716 4068 11744
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5592 11716 5641 11744
rect 5592 11704 5598 11716
rect 5629 11713 5641 11716
rect 5675 11713 5687 11747
rect 6822 11744 6828 11756
rect 6783 11716 6828 11744
rect 5629 11707 5687 11713
rect 6822 11704 6828 11716
rect 6880 11704 6886 11756
rect 8202 11704 8208 11756
rect 8260 11744 8266 11756
rect 8496 11744 8524 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10244 11812 10272 11852
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 10376 11852 10609 11880
rect 10376 11840 10382 11852
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 10597 11843 10655 11849
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 12802 11880 12808 11892
rect 10744 11852 12808 11880
rect 10744 11840 10750 11852
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 13173 11883 13231 11889
rect 13173 11880 13185 11883
rect 13044 11852 13185 11880
rect 13044 11840 13050 11852
rect 13173 11849 13185 11852
rect 13219 11849 13231 11883
rect 13173 11843 13231 11849
rect 14829 11883 14887 11889
rect 14829 11849 14841 11883
rect 14875 11880 14887 11883
rect 15102 11880 15108 11892
rect 14875 11852 15108 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 15102 11840 15108 11852
rect 15160 11840 15166 11892
rect 16393 11883 16451 11889
rect 16393 11880 16405 11883
rect 15304 11852 16405 11880
rect 10244 11784 11744 11812
rect 11716 11756 11744 11784
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 15304 11812 15332 11852
rect 16393 11849 16405 11852
rect 16439 11849 16451 11883
rect 16393 11843 16451 11849
rect 20622 11840 20628 11892
rect 20680 11880 20686 11892
rect 20809 11883 20867 11889
rect 20809 11880 20821 11883
rect 20680 11852 20821 11880
rect 20680 11840 20686 11852
rect 20809 11849 20821 11852
rect 20855 11849 20867 11883
rect 20809 11843 20867 11849
rect 17954 11812 17960 11824
rect 13872 11784 15332 11812
rect 15396 11784 17960 11812
rect 13872 11772 13878 11784
rect 8260 11716 8524 11744
rect 8260 11704 8266 11716
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9548 11716 9597 11744
rect 9548 11704 9554 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 10318 11704 10324 11756
rect 10376 11744 10382 11756
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10376 11716 11161 11744
rect 10376 11704 10382 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11698 11704 11704 11756
rect 11756 11704 11762 11756
rect 13722 11744 13728 11756
rect 13683 11716 13728 11744
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 15286 11744 15292 11756
rect 15247 11716 15292 11744
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15396 11753 15424 11784
rect 17954 11772 17960 11784
rect 18012 11772 18018 11824
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17126 11744 17132 11756
rect 17083 11716 17132 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 18322 11744 18328 11756
rect 18283 11716 18328 11744
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 3844 11648 3893 11676
rect 3844 11636 3850 11648
rect 3881 11645 3893 11648
rect 3927 11645 3939 11679
rect 3881 11639 3939 11645
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4154 11676 4160 11688
rect 4019 11648 4160 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 8754 11676 8760 11688
rect 4304 11648 8760 11676
rect 4304 11636 4310 11648
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 9306 11636 9312 11688
rect 9364 11676 9370 11688
rect 9364 11648 9536 11676
rect 9364 11636 9370 11648
rect 6638 11608 6644 11620
rect 5460 11580 6644 11608
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4798 11540 4804 11552
rect 4212 11512 4804 11540
rect 4212 11500 4218 11512
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5460 11549 5488 11580
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 7092 11611 7150 11617
rect 7092 11577 7104 11611
rect 7138 11608 7150 11611
rect 8478 11608 8484 11620
rect 7138 11580 8484 11608
rect 7138 11577 7150 11580
rect 7092 11571 7150 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 9508 11617 9536 11648
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10410 11676 10416 11688
rect 10100 11648 10416 11676
rect 10100 11636 10106 11648
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 11054 11676 11060 11688
rect 11015 11648 11060 11676
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 18138 11676 18144 11688
rect 11348 11648 17908 11676
rect 18099 11648 18144 11676
rect 9401 11611 9459 11617
rect 9401 11608 9413 11611
rect 8588 11580 9413 11608
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5132 11512 5457 11540
rect 5132 11500 5138 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5445 11503 5503 11509
rect 5537 11543 5595 11549
rect 5537 11509 5549 11543
rect 5583 11540 5595 11543
rect 5626 11540 5632 11552
rect 5583 11512 5632 11540
rect 5583 11509 5595 11512
rect 5537 11503 5595 11509
rect 5626 11500 5632 11512
rect 5684 11540 5690 11552
rect 8202 11540 8208 11552
rect 5684 11512 8208 11540
rect 5684 11500 5690 11512
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8588 11540 8616 11580
rect 9401 11577 9413 11580
rect 9447 11577 9459 11611
rect 9401 11571 9459 11577
rect 9493 11611 9551 11617
rect 9493 11577 9505 11611
rect 9539 11577 9551 11611
rect 9493 11571 9551 11577
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 10965 11611 11023 11617
rect 10965 11608 10977 11611
rect 10744 11580 10977 11608
rect 10744 11568 10750 11580
rect 10965 11577 10977 11580
rect 11011 11608 11023 11611
rect 11348 11608 11376 11648
rect 13541 11611 13599 11617
rect 13541 11608 13553 11611
rect 11011 11580 11376 11608
rect 12719 11580 13553 11608
rect 11011 11577 11023 11580
rect 10965 11571 11023 11577
rect 8352 11512 8616 11540
rect 8352 11500 8358 11512
rect 8754 11500 8760 11552
rect 8812 11540 8818 11552
rect 11882 11540 11888 11552
rect 8812 11512 11888 11540
rect 8812 11500 8818 11512
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 12719 11540 12747 11580
rect 13541 11577 13553 11580
rect 13587 11608 13599 11611
rect 16022 11608 16028 11620
rect 13587 11580 16028 11608
rect 13587 11577 13599 11580
rect 13541 11571 13599 11577
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 17770 11608 17776 11620
rect 16316 11580 17776 11608
rect 12584 11512 12747 11540
rect 12584 11500 12590 11512
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 13044 11512 13645 11540
rect 13044 11500 13050 11512
rect 13633 11509 13645 11512
rect 13679 11509 13691 11543
rect 13633 11503 13691 11509
rect 15197 11543 15255 11549
rect 15197 11509 15209 11543
rect 15243 11540 15255 11543
rect 16316 11540 16344 11580
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 17880 11608 17908 11648
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19702 11685 19708 11688
rect 19429 11679 19487 11685
rect 19429 11676 19441 11679
rect 19300 11648 19441 11676
rect 19300 11636 19306 11648
rect 19429 11645 19441 11648
rect 19475 11645 19487 11679
rect 19429 11639 19487 11645
rect 19696 11639 19708 11685
rect 19760 11676 19766 11688
rect 19760 11648 19796 11676
rect 19702 11636 19708 11639
rect 19760 11636 19766 11648
rect 18966 11608 18972 11620
rect 17880 11580 18972 11608
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 16758 11540 16764 11552
rect 15243 11512 16344 11540
rect 16719 11512 16764 11540
rect 15243 11509 15255 11512
rect 15197 11503 15255 11509
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 16853 11543 16911 11549
rect 16853 11509 16865 11543
rect 16899 11540 16911 11543
rect 17586 11540 17592 11552
rect 16899 11512 17592 11540
rect 16899 11509 16911 11512
rect 16853 11503 16911 11509
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 4246 11336 4252 11348
rect 1995 11308 4252 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 4246 11296 4252 11308
rect 4304 11296 4310 11348
rect 4430 11336 4436 11348
rect 4391 11308 4436 11336
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 6178 11336 6184 11348
rect 5583 11308 6184 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6457 11339 6515 11345
rect 6457 11336 6469 11339
rect 6328 11308 6469 11336
rect 6328 11296 6334 11308
rect 6457 11305 6469 11308
rect 6503 11305 6515 11339
rect 6457 11299 6515 11305
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 8386 11336 8392 11348
rect 6871 11308 8392 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9398 11336 9404 11348
rect 8536 11308 9404 11336
rect 8536 11296 8542 11308
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9861 11339 9919 11345
rect 9861 11305 9873 11339
rect 9907 11336 9919 11339
rect 10042 11336 10048 11348
rect 9907 11308 10048 11336
rect 9907 11305 9919 11308
rect 9861 11299 9919 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 11238 11336 11244 11348
rect 10152 11308 11244 11336
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 7190 11268 7196 11280
rect 3007 11240 7196 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 8128 11240 8524 11268
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11200 4307 11203
rect 5166 11200 5172 11212
rect 4295 11172 5172 11200
rect 4295 11169 4307 11172
rect 4249 11163 4307 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5399 11172 6776 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 5810 11132 5816 11144
rect 5316 11104 5816 11132
rect 5316 11092 5322 11104
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 6362 11064 6368 11076
rect 4948 11036 6368 11064
rect 4948 11024 4954 11036
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 6748 11064 6776 11172
rect 6914 11132 6920 11144
rect 6875 11104 6920 11132
rect 6914 11092 6920 11104
rect 6972 11092 6978 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 8128 11132 8156 11240
rect 8386 11200 8392 11212
rect 8347 11172 8392 11200
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8496 11200 8524 11240
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8938 11268 8944 11280
rect 8628 11240 8944 11268
rect 8628 11228 8634 11240
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 9582 11200 9588 11212
rect 8496 11172 9588 11200
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10152 11200 10180 11308
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 12032 11308 12173 11336
rect 12032 11296 12038 11308
rect 12161 11305 12173 11308
rect 12207 11336 12219 11339
rect 12618 11336 12624 11348
rect 12207 11308 12624 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12618 11296 12624 11308
rect 12676 11296 12682 11348
rect 13446 11336 13452 11348
rect 13407 11308 13452 11336
rect 13446 11296 13452 11308
rect 13504 11296 13510 11348
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14550 11336 14556 11348
rect 13955 11308 14556 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15381 11339 15439 11345
rect 15381 11305 15393 11339
rect 15427 11336 15439 11339
rect 16666 11336 16672 11348
rect 15427 11308 16672 11336
rect 15427 11305 15439 11308
rect 15381 11299 15439 11305
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 16776 11308 17356 11336
rect 10870 11268 10876 11280
rect 9732 11172 10180 11200
rect 10336 11240 10732 11268
rect 10831 11240 10876 11268
rect 9732 11160 9738 11172
rect 7147 11104 8156 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8481 11135 8539 11141
rect 8481 11132 8493 11135
rect 8260 11104 8493 11132
rect 8260 11092 8266 11104
rect 8481 11101 8493 11104
rect 8527 11132 8539 11135
rect 8570 11132 8576 11144
rect 8527 11104 8576 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8665 11135 8723 11141
rect 8665 11101 8677 11135
rect 8711 11132 8723 11135
rect 10336 11132 10364 11240
rect 10502 11160 10508 11212
rect 10560 11160 10566 11212
rect 10704 11200 10732 11240
rect 10870 11228 10876 11240
rect 10928 11228 10934 11280
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 11882 11268 11888 11280
rect 11664 11240 11888 11268
rect 11664 11228 11670 11240
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 13262 11228 13268 11280
rect 13320 11268 13326 11280
rect 16776 11268 16804 11308
rect 13320 11240 16804 11268
rect 13320 11228 13326 11240
rect 16850 11228 16856 11280
rect 16908 11268 16914 11280
rect 17190 11271 17248 11277
rect 17190 11268 17202 11271
rect 16908 11240 17202 11268
rect 16908 11228 16914 11240
rect 17190 11237 17202 11240
rect 17236 11237 17248 11271
rect 17328 11268 17356 11308
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 18012 11308 18337 11336
rect 18012 11296 18018 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 19518 11296 19524 11348
rect 19576 11336 19582 11348
rect 19705 11339 19763 11345
rect 19705 11336 19717 11339
rect 19576 11308 19717 11336
rect 19576 11296 19582 11308
rect 19705 11305 19717 11308
rect 19751 11305 19763 11339
rect 19705 11299 19763 11305
rect 19061 11271 19119 11277
rect 19061 11268 19073 11271
rect 17328 11240 19073 11268
rect 17190 11231 17248 11237
rect 19061 11237 19073 11240
rect 19107 11268 19119 11271
rect 19613 11271 19671 11277
rect 19613 11268 19625 11271
rect 19107 11240 19625 11268
rect 19107 11237 19119 11240
rect 19061 11231 19119 11237
rect 19613 11237 19625 11240
rect 19659 11237 19671 11271
rect 19613 11231 19671 11237
rect 11054 11200 11060 11212
rect 10704 11172 11060 11200
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 13817 11203 13875 11209
rect 13817 11169 13829 11203
rect 13863 11200 13875 11203
rect 14274 11200 14280 11212
rect 13863 11172 14280 11200
rect 13863 11169 13875 11172
rect 13817 11163 13875 11169
rect 14274 11160 14280 11172
rect 14332 11200 14338 11212
rect 15654 11200 15660 11212
rect 14332 11172 15660 11200
rect 14332 11160 14338 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 18138 11200 18144 11212
rect 15795 11172 18144 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 18138 11160 18144 11172
rect 18196 11160 18202 11212
rect 8711 11104 10364 11132
rect 8711 11101 8723 11104
rect 8665 11095 8723 11101
rect 7926 11064 7932 11076
rect 6748 11036 7932 11064
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 10520 11064 10548 11160
rect 11072 11132 11100 11160
rect 13722 11132 13728 11144
rect 11072 11104 13728 11132
rect 13722 11092 13728 11104
rect 13780 11132 13786 11144
rect 14001 11135 14059 11141
rect 14001 11132 14013 11135
rect 13780 11104 14013 11132
rect 13780 11092 13786 11104
rect 14001 11101 14013 11104
rect 14047 11101 14059 11135
rect 14001 11095 14059 11101
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15378 11132 15384 11144
rect 14424 11104 15384 11132
rect 14424 11092 14430 11104
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 15841 11135 15899 11141
rect 15841 11101 15853 11135
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 8067 11036 10548 11064
rect 15856 11064 15884 11095
rect 15930 11092 15936 11144
rect 15988 11132 15994 11144
rect 16942 11132 16948 11144
rect 15988 11104 16033 11132
rect 16903 11104 16948 11132
rect 15988 11092 15994 11104
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 18782 11132 18788 11144
rect 18104 11104 18788 11132
rect 18104 11092 18110 11104
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 19886 11132 19892 11144
rect 19847 11104 19892 11132
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 18690 11064 18696 11076
rect 15856 11036 16988 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 290 10956 296 11008
rect 348 10996 354 11008
rect 6914 10996 6920 11008
rect 348 10968 6920 10996
rect 348 10956 354 10968
rect 6914 10956 6920 10968
rect 6972 10996 6978 11008
rect 8202 10996 8208 11008
rect 6972 10968 8208 10996
rect 6972 10956 6978 10968
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 14182 10996 14188 11008
rect 10376 10968 14188 10996
rect 10376 10956 10382 10968
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 16960 10996 16988 11036
rect 17880 11036 18696 11064
rect 17880 10996 17908 11036
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 19245 11067 19303 11073
rect 19245 11033 19257 11067
rect 19291 11064 19303 11067
rect 19610 11064 19616 11076
rect 19291 11036 19616 11064
rect 19291 11033 19303 11036
rect 19245 11027 19303 11033
rect 19610 11024 19616 11036
rect 19668 11024 19674 11076
rect 16960 10968 17908 10996
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7248 10764 9260 10792
rect 7248 10752 7254 10764
rect 5810 10724 5816 10736
rect 5771 10696 5816 10724
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 9232 10724 9260 10764
rect 9398 10752 9404 10804
rect 9456 10792 9462 10804
rect 9493 10795 9551 10801
rect 9493 10792 9505 10795
rect 9456 10764 9505 10792
rect 9456 10752 9462 10764
rect 9493 10761 9505 10764
rect 9539 10761 9551 10795
rect 9493 10755 9551 10761
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 9999 10764 13676 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 10686 10724 10692 10736
rect 9232 10696 10692 10724
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 12158 10724 12164 10736
rect 12119 10696 12164 10724
rect 12158 10684 12164 10696
rect 12216 10684 12222 10736
rect 13648 10724 13676 10764
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 13780 10764 13829 10792
rect 13780 10752 13786 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 16850 10792 16856 10804
rect 13817 10755 13875 10761
rect 13924 10764 16436 10792
rect 16811 10764 16856 10792
rect 13924 10724 13952 10764
rect 13648 10696 13952 10724
rect 16408 10724 16436 10764
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 16942 10752 16948 10804
rect 17000 10792 17006 10804
rect 17681 10795 17739 10801
rect 17681 10792 17693 10795
rect 17000 10764 17693 10792
rect 17000 10752 17006 10764
rect 17681 10761 17693 10764
rect 17727 10761 17739 10795
rect 17681 10755 17739 10761
rect 18233 10795 18291 10801
rect 18233 10761 18245 10795
rect 18279 10792 18291 10795
rect 18874 10792 18880 10804
rect 18279 10764 18880 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 17402 10724 17408 10736
rect 16408 10696 17408 10724
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 3602 10656 3608 10668
rect 3563 10628 3608 10656
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 9214 10616 9220 10668
rect 9272 10656 9278 10668
rect 10597 10659 10655 10665
rect 9272 10628 10548 10656
rect 9272 10616 9278 10628
rect 2593 10591 2651 10597
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 3878 10588 3884 10600
rect 2639 10560 3884 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 4525 10523 4583 10529
rect 4525 10489 4537 10523
rect 4571 10520 4583 10523
rect 4614 10520 4620 10532
rect 4571 10492 4620 10520
rect 4571 10489 4583 10492
rect 4525 10483 4583 10489
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 5644 10452 5672 10551
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6788 10560 6837 10588
rect 6788 10548 6794 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 7098 10520 7104 10532
rect 7059 10492 7104 10520
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 7190 10452 7196 10464
rect 5644 10424 7196 10452
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 8128 10452 8156 10551
rect 8202 10548 8208 10600
rect 8260 10588 8266 10600
rect 10413 10591 10471 10597
rect 10413 10588 10425 10591
rect 8260 10560 10425 10588
rect 8260 10548 8266 10560
rect 10413 10557 10425 10560
rect 10459 10557 10471 10591
rect 10520 10588 10548 10628
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 17696 10656 17724 10755
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19334 10792 19340 10804
rect 19168 10764 19340 10792
rect 19168 10668 19196 10764
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 19150 10656 19156 10668
rect 10643 10628 10916 10656
rect 17696 10628 19156 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10520 10560 10793 10588
rect 10413 10551 10471 10557
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10888 10588 10916 10628
rect 19150 10616 19156 10628
rect 19208 10616 19214 10668
rect 12437 10591 12495 10597
rect 10888 10560 11376 10588
rect 10781 10551 10839 10557
rect 11348 10532 11376 10560
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 15286 10588 15292 10600
rect 12483 10560 15292 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 15286 10548 15292 10560
rect 15344 10588 15350 10600
rect 15473 10591 15531 10597
rect 15473 10588 15485 10591
rect 15344 10560 15485 10588
rect 15344 10548 15350 10560
rect 15473 10557 15485 10560
rect 15519 10557 15531 10591
rect 15473 10551 15531 10557
rect 15740 10591 15798 10597
rect 15740 10557 15752 10591
rect 15786 10588 15798 10591
rect 16482 10588 16488 10600
rect 15786 10560 16488 10588
rect 15786 10557 15798 10560
rect 15740 10551 15798 10557
rect 11054 10529 11060 10532
rect 8380 10523 8438 10529
rect 8380 10489 8392 10523
rect 8426 10520 8438 10523
rect 11048 10520 11060 10529
rect 8426 10492 10548 10520
rect 11015 10492 11060 10520
rect 8426 10489 8438 10492
rect 8380 10483 8438 10489
rect 9122 10452 9128 10464
rect 8128 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9950 10452 9956 10464
rect 9732 10424 9956 10452
rect 9732 10412 9738 10424
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 10318 10452 10324 10464
rect 10279 10424 10324 10452
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 10520 10452 10548 10492
rect 11048 10483 11060 10492
rect 11054 10480 11060 10483
rect 11112 10480 11118 10532
rect 11330 10480 11336 10532
rect 11388 10520 11394 10532
rect 12682 10523 12740 10529
rect 12682 10520 12694 10523
rect 11388 10492 12694 10520
rect 11388 10480 11394 10492
rect 12682 10489 12694 10492
rect 12728 10489 12740 10523
rect 15488 10520 15516 10551
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 17862 10588 17868 10600
rect 17823 10560 17868 10588
rect 17862 10548 17868 10560
rect 17920 10548 17926 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 16942 10520 16948 10532
rect 15488 10492 16948 10520
rect 12682 10483 12740 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 18064 10520 18092 10551
rect 17184 10492 18092 10520
rect 19420 10523 19478 10529
rect 17184 10480 17190 10492
rect 19420 10489 19432 10523
rect 19466 10520 19478 10523
rect 19886 10520 19892 10532
rect 19466 10492 19892 10520
rect 19466 10489 19478 10492
rect 19420 10483 19478 10489
rect 19886 10480 19892 10492
rect 19944 10520 19950 10532
rect 20438 10520 20444 10532
rect 19944 10492 20444 10520
rect 19944 10480 19950 10492
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 20162 10452 20168 10464
rect 10520 10424 20168 10452
rect 20162 10412 20168 10424
rect 20220 10452 20226 10464
rect 20533 10455 20591 10461
rect 20533 10452 20545 10455
rect 20220 10424 20545 10452
rect 20220 10412 20226 10424
rect 20533 10421 20545 10424
rect 20579 10421 20591 10455
rect 20533 10415 20591 10421
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4798 10248 4804 10260
rect 4755 10220 4804 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 5997 10251 6055 10257
rect 5997 10217 6009 10251
rect 6043 10248 6055 10251
rect 6822 10248 6828 10260
rect 6043 10220 6828 10248
rect 6043 10217 6055 10220
rect 5997 10211 6055 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8202 10248 8208 10260
rect 8067 10220 8208 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8478 10248 8484 10260
rect 8439 10220 8484 10248
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 10042 10248 10048 10260
rect 8628 10220 10048 10248
rect 8628 10208 8634 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10318 10208 10324 10260
rect 10376 10248 10382 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 10376 10220 12173 10248
rect 10376 10208 10382 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13909 10251 13967 10257
rect 13909 10248 13921 10251
rect 12768 10220 13921 10248
rect 12768 10208 12774 10220
rect 13909 10217 13921 10220
rect 13955 10217 13967 10251
rect 13909 10211 13967 10217
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 19518 10248 19524 10260
rect 16632 10220 19524 10248
rect 16632 10208 16638 10220
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 15556 10183 15614 10189
rect 7156 10152 15148 10180
rect 7156 10140 7162 10152
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10081 5871 10115
rect 5813 10075 5871 10081
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7558 10112 7564 10124
rect 6963 10084 7564 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 5828 10044 5856 10075
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10112 8447 10115
rect 10220 10115 10278 10121
rect 10220 10112 10232 10115
rect 8435 10084 8616 10112
rect 8435 10081 8447 10084
rect 8389 10075 8447 10081
rect 8478 10044 8484 10056
rect 5828 10016 8484 10044
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 8588 9976 8616 10084
rect 8680 10084 10232 10112
rect 8680 10053 8708 10084
rect 10220 10081 10232 10084
rect 10266 10112 10278 10115
rect 12526 10112 12532 10124
rect 10266 10084 11008 10112
rect 12487 10084 12532 10112
rect 10266 10081 10278 10084
rect 10220 10075 10278 10081
rect 10980 10056 11008 10084
rect 12526 10072 12532 10084
rect 12584 10072 12590 10124
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13412 10084 13737 10112
rect 13412 10072 13418 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 14734 10072 14740 10124
rect 14792 10112 14798 10124
rect 15013 10115 15071 10121
rect 15013 10112 15025 10115
rect 14792 10084 15025 10112
rect 14792 10072 14798 10084
rect 15013 10081 15025 10084
rect 15059 10081 15071 10115
rect 15120 10112 15148 10152
rect 15556 10149 15568 10183
rect 15602 10180 15614 10183
rect 15930 10180 15936 10192
rect 15602 10152 15936 10180
rect 15602 10149 15614 10152
rect 15556 10143 15614 10149
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 16390 10140 16396 10192
rect 16448 10180 16454 10192
rect 19153 10183 19211 10189
rect 19153 10180 19165 10183
rect 16448 10152 19165 10180
rect 16448 10140 16454 10152
rect 19153 10149 19165 10152
rect 19199 10149 19211 10183
rect 19153 10143 19211 10149
rect 17494 10112 17500 10124
rect 15120 10084 16795 10112
rect 17455 10084 17500 10112
rect 15013 10075 15071 10081
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9180 10016 9965 10044
rect 9180 10004 9186 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 10962 10004 10968 10056
rect 11020 10044 11026 10056
rect 11020 10016 11468 10044
rect 11020 10004 11026 10016
rect 9674 9976 9680 9988
rect 5408 9948 7227 9976
rect 8588 9948 9680 9976
rect 5408 9936 5414 9948
rect 7098 9908 7104 9920
rect 7059 9880 7104 9908
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 7199 9908 7227 9948
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 11330 9976 11336 9988
rect 11291 9948 11336 9976
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 11440 9976 11468 10016
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 12492 10016 12633 10044
rect 12492 10004 12498 10016
rect 12621 10013 12633 10016
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 12713 10007 12771 10013
rect 12728 9976 12756 10007
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 11440 9948 12756 9976
rect 16482 9936 16488 9988
rect 16540 9976 16546 9988
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 16540 9948 16681 9976
rect 16540 9936 16546 9948
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16767 9976 16795 10084
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 19168 10084 19257 10112
rect 17678 10044 17684 10056
rect 17639 10016 17684 10044
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 17954 9976 17960 9988
rect 16767 9948 17960 9976
rect 16669 9939 16727 9945
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 19168 9976 19196 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 19334 10044 19340 10056
rect 19295 10016 19340 10044
rect 19334 10004 19340 10016
rect 19392 10004 19398 10056
rect 19242 9976 19248 9988
rect 19168 9948 19248 9976
rect 19242 9936 19248 9948
rect 19300 9936 19306 9988
rect 12158 9908 12164 9920
rect 7199 9880 12164 9908
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 14829 9911 14887 9917
rect 14829 9877 14841 9911
rect 14875 9908 14887 9911
rect 17402 9908 17408 9920
rect 14875 9880 17408 9908
rect 14875 9877 14887 9880
rect 14829 9871 14887 9877
rect 17402 9868 17408 9880
rect 17460 9908 17466 9920
rect 17862 9908 17868 9920
rect 17460 9880 17868 9908
rect 17460 9868 17466 9880
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18782 9908 18788 9920
rect 18743 9880 18788 9908
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 3510 9664 3516 9716
rect 3568 9704 3574 9716
rect 10505 9707 10563 9713
rect 3568 9676 10456 9704
rect 3568 9664 3574 9676
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 8754 9636 8760 9648
rect 8536 9608 8760 9636
rect 8536 9596 8542 9608
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 5994 9568 6000 9580
rect 5767 9540 6000 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 5994 9528 6000 9540
rect 6052 9528 6058 9580
rect 10428 9568 10456 9676
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10962 9704 10968 9716
rect 10551 9676 10968 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 19334 9704 19340 9716
rect 11072 9676 19340 9704
rect 11072 9568 11100 9676
rect 19334 9664 19340 9676
rect 19392 9664 19398 9716
rect 12621 9639 12679 9645
rect 10428 9540 11100 9568
rect 11164 9608 12572 9636
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 6696 9472 6929 9500
rect 6696 9460 6702 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 8294 9500 8300 9512
rect 6917 9463 6975 9469
rect 8036 9472 8300 9500
rect 3605 9435 3663 9441
rect 3605 9401 3617 9435
rect 3651 9432 3663 9435
rect 3697 9435 3755 9441
rect 3697 9432 3709 9435
rect 3651 9404 3709 9432
rect 3651 9401 3663 9404
rect 3605 9395 3663 9401
rect 3697 9401 3709 9404
rect 3743 9432 3755 9435
rect 4798 9432 4804 9444
rect 3743 9404 4804 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4798 9392 4804 9404
rect 4856 9392 4862 9444
rect 7184 9435 7242 9441
rect 7184 9401 7196 9435
rect 7230 9432 7242 9435
rect 7742 9432 7748 9444
rect 7230 9404 7748 9432
rect 7230 9401 7242 9404
rect 7184 9395 7242 9401
rect 7742 9392 7748 9404
rect 7800 9392 7806 9444
rect 4709 9367 4767 9373
rect 4709 9333 4721 9367
rect 4755 9364 4767 9367
rect 8036 9364 8064 9472
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 9122 9500 9128 9512
rect 9083 9472 9128 9500
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 11164 9500 11192 9608
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 11974 9568 11980 9580
rect 11379 9540 11980 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12544 9568 12572 9608
rect 12621 9605 12633 9639
rect 12667 9636 12679 9639
rect 12894 9636 12900 9648
rect 12667 9608 12900 9636
rect 12667 9605 12679 9608
rect 12621 9599 12679 9605
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13044 9608 14872 9636
rect 13044 9596 13050 9608
rect 13262 9568 13268 9580
rect 12544 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14844 9568 14872 9608
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 16853 9639 16911 9645
rect 16853 9636 16865 9639
rect 15528 9608 16865 9636
rect 15528 9596 15534 9608
rect 16853 9605 16865 9608
rect 16899 9605 16911 9639
rect 16853 9599 16911 9605
rect 18509 9639 18567 9645
rect 18509 9605 18521 9639
rect 18555 9636 18567 9639
rect 18598 9636 18604 9648
rect 18555 9608 18604 9636
rect 18555 9605 18567 9608
rect 18509 9599 18567 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 20438 9596 20444 9648
rect 20496 9636 20502 9648
rect 20809 9639 20867 9645
rect 20809 9636 20821 9639
rect 20496 9608 20821 9636
rect 20496 9596 20502 9608
rect 20809 9605 20821 9608
rect 20855 9605 20867 9639
rect 20809 9599 20867 9605
rect 15746 9568 15752 9580
rect 14844 9540 15599 9568
rect 15707 9540 15752 9568
rect 12434 9500 12440 9512
rect 9272 9472 11192 9500
rect 12395 9472 12440 9500
rect 9272 9460 9278 9472
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13188 9472 14013 9500
rect 9392 9435 9450 9441
rect 9392 9401 9404 9435
rect 9438 9432 9450 9435
rect 9582 9432 9588 9444
rect 9438 9404 9588 9432
rect 9438 9401 9450 9404
rect 9392 9395 9450 9401
rect 9582 9392 9588 9404
rect 9640 9432 9646 9444
rect 9640 9404 10640 9432
rect 9640 9392 9646 9404
rect 8294 9364 8300 9376
rect 4755 9336 8064 9364
rect 8255 9336 8300 9364
rect 4755 9333 4767 9336
rect 4709 9327 4767 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9490 9364 9496 9376
rect 8904 9336 9496 9364
rect 8904 9324 8910 9336
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 10612 9364 10640 9404
rect 10686 9392 10692 9444
rect 10744 9432 10750 9444
rect 13188 9432 13216 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14734 9500 14740 9512
rect 14608 9472 14740 9500
rect 14608 9460 14614 9472
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 15571 9500 15599 9540
rect 15746 9528 15752 9540
rect 15804 9528 15810 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 19150 9568 19156 9580
rect 17736 9540 19156 9568
rect 17736 9528 17742 9540
rect 19150 9528 19156 9540
rect 19208 9568 19214 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19208 9540 19441 9568
rect 19208 9528 19214 9540
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 15571 9472 16681 9500
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18012 9472 18337 9500
rect 18012 9460 18018 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 10744 9404 13216 9432
rect 15473 9435 15531 9441
rect 10744 9392 10750 9404
rect 15473 9401 15485 9435
rect 15519 9401 15531 9435
rect 15473 9395 15531 9401
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 15654 9432 15660 9444
rect 15611 9404 15660 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 13446 9364 13452 9376
rect 10612 9336 13452 9364
rect 13446 9324 13452 9336
rect 13504 9324 13510 9376
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 13909 9367 13967 9373
rect 13596 9336 13641 9364
rect 13596 9324 13602 9336
rect 13909 9333 13921 9367
rect 13955 9364 13967 9367
rect 14090 9364 14096 9376
rect 13955 9336 14096 9364
rect 13955 9333 13967 9336
rect 13909 9327 13967 9333
rect 14090 9324 14096 9336
rect 14148 9364 14154 9376
rect 14550 9364 14556 9376
rect 14148 9336 14556 9364
rect 14148 9324 14154 9336
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15105 9367 15163 9373
rect 15105 9333 15117 9367
rect 15151 9364 15163 9367
rect 15286 9364 15292 9376
rect 15151 9336 15292 9364
rect 15151 9333 15163 9336
rect 15105 9327 15163 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15378 9324 15384 9376
rect 15436 9364 15442 9376
rect 15479 9364 15507 9395
rect 15654 9392 15660 9404
rect 15712 9392 15718 9444
rect 19696 9435 19754 9441
rect 19696 9401 19708 9435
rect 19742 9432 19754 9435
rect 19794 9432 19800 9444
rect 19742 9404 19800 9432
rect 19742 9401 19754 9404
rect 19696 9395 19754 9401
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 15436 9336 15507 9364
rect 15436 9324 15442 9336
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 4617 9163 4675 9169
rect 4617 9129 4629 9163
rect 4663 9160 4675 9163
rect 4890 9160 4896 9172
rect 4663 9132 4896 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 4890 9120 4896 9132
rect 4948 9120 4954 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7800 9132 8033 9160
rect 7800 9120 7806 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 8021 9123 8079 9129
rect 8202 9120 8208 9172
rect 8260 9160 8266 9172
rect 12986 9160 12992 9172
rect 8260 9132 12992 9160
rect 8260 9120 8266 9132
rect 12986 9120 12992 9132
rect 13044 9120 13050 9172
rect 13633 9163 13691 9169
rect 13633 9129 13645 9163
rect 13679 9160 13691 9163
rect 15378 9160 15384 9172
rect 13679 9132 15384 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 15378 9120 15384 9132
rect 15436 9120 15442 9172
rect 16390 9160 16396 9172
rect 16351 9132 16396 9160
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 16853 9163 16911 9169
rect 16853 9129 16865 9163
rect 16899 9160 16911 9163
rect 17770 9160 17776 9172
rect 16899 9132 17776 9160
rect 16899 9129 16911 9132
rect 16853 9123 16911 9129
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 19334 9160 19340 9172
rect 17972 9132 18184 9160
rect 19295 9132 19340 9160
rect 5629 9095 5687 9101
rect 5629 9061 5641 9095
rect 5675 9092 5687 9095
rect 16761 9095 16819 9101
rect 16761 9092 16773 9095
rect 5675 9064 16773 9092
rect 5675 9061 5687 9064
rect 5629 9055 5687 9061
rect 16761 9061 16773 9064
rect 16807 9061 16819 9095
rect 17034 9092 17040 9104
rect 16761 9055 16819 9061
rect 16960 9064 17040 9092
rect 6638 9024 6644 9036
rect 6599 8996 6644 9024
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 6908 9027 6966 9033
rect 6908 8993 6920 9027
rect 6954 9024 6966 9027
rect 7650 9024 7656 9036
rect 6954 8996 7656 9024
rect 6954 8993 6966 8996
rect 6908 8987 6966 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 9030 9024 9036 9036
rect 8991 8996 9036 9024
rect 9030 8984 9036 8996
rect 9088 8984 9094 9036
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 9180 8996 10701 9024
rect 9180 8984 9186 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 10956 9027 11014 9033
rect 10956 8993 10968 9027
rect 11002 9024 11014 9027
rect 11238 9024 11244 9036
rect 11002 8996 11244 9024
rect 11002 8993 11014 8996
rect 10956 8987 11014 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 13998 9024 14004 9036
rect 13959 8996 14004 9024
rect 13998 8984 14004 8996
rect 14056 8984 14062 9036
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 9024 14151 9027
rect 15289 9027 15347 9033
rect 14139 8996 15240 9024
rect 14139 8993 14151 8996
rect 14093 8987 14151 8993
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8956 9735 8959
rect 10134 8956 10140 8968
rect 9723 8928 10140 8956
rect 9723 8925 9735 8928
rect 9677 8919 9735 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 11698 8916 11704 8968
rect 11756 8956 11762 8968
rect 14108 8956 14136 8987
rect 11756 8928 14136 8956
rect 11756 8916 11762 8928
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 15212 8956 15240 8996
rect 15289 8993 15301 9027
rect 15335 9024 15347 9027
rect 16960 9024 16988 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 17972 9024 18000 9132
rect 15335 8996 16988 9024
rect 17052 8996 18000 9024
rect 18156 9024 18184 9132
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 18213 9027 18271 9033
rect 18213 9024 18225 9027
rect 18156 8996 18225 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 17052 8965 17080 8996
rect 18213 8993 18225 8996
rect 18259 9024 18271 9027
rect 19150 9024 19156 9036
rect 18259 8996 19156 9024
rect 18259 8993 18271 8996
rect 18213 8987 18271 8993
rect 19150 8984 19156 8996
rect 19208 8984 19214 9036
rect 17037 8959 17095 8965
rect 14240 8928 14285 8956
rect 15212 8928 16344 8956
rect 14240 8916 14246 8928
rect 10686 8888 10692 8900
rect 8496 8860 10692 8888
rect 2866 8780 2872 8832
rect 2924 8820 2930 8832
rect 8496 8820 8524 8860
rect 10686 8848 10692 8860
rect 10744 8848 10750 8900
rect 13814 8888 13820 8900
rect 11624 8860 13820 8888
rect 2924 8792 8524 8820
rect 2924 8780 2930 8792
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 8849 8823 8907 8829
rect 8849 8820 8861 8823
rect 8628 8792 8861 8820
rect 8628 8780 8634 8792
rect 8849 8789 8861 8792
rect 8895 8789 8907 8823
rect 8849 8783 8907 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 11624 8820 11652 8860
rect 13814 8848 13820 8860
rect 13872 8848 13878 8900
rect 13906 8848 13912 8900
rect 13964 8888 13970 8900
rect 15473 8891 15531 8897
rect 15473 8888 15485 8891
rect 13964 8860 15485 8888
rect 13964 8848 13970 8860
rect 15473 8857 15485 8860
rect 15519 8857 15531 8891
rect 16316 8888 16344 8928
rect 17037 8925 17049 8959
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 17678 8916 17684 8968
rect 17736 8956 17742 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17736 8928 17969 8956
rect 17736 8916 17742 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 17862 8888 17868 8900
rect 16316 8860 17868 8888
rect 15473 8851 15531 8857
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 12066 8820 12072 8832
rect 9916 8792 11652 8820
rect 12027 8792 12072 8820
rect 9916 8780 9922 8792
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 17770 8820 17776 8832
rect 14056 8792 17776 8820
rect 14056 8780 14062 8792
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 11425 8619 11483 8625
rect 11425 8585 11437 8619
rect 11471 8616 11483 8619
rect 15654 8616 15660 8628
rect 11471 8588 15660 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 16114 8616 16120 8628
rect 15804 8588 16120 8616
rect 15804 8576 15810 8588
rect 16114 8576 16120 8588
rect 16172 8616 16178 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16172 8588 16405 8616
rect 16172 8576 16178 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 7929 8551 7987 8557
rect 7929 8517 7941 8551
rect 7975 8548 7987 8551
rect 12342 8548 12348 8560
rect 7975 8520 12348 8548
rect 7975 8517 7987 8520
rect 7929 8511 7987 8517
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 14182 8548 14188 8560
rect 14095 8520 14188 8548
rect 14182 8508 14188 8520
rect 14240 8508 14246 8560
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17221 8551 17279 8557
rect 17221 8548 17233 8551
rect 16816 8520 17233 8548
rect 16816 8508 16822 8520
rect 17221 8517 17233 8520
rect 17267 8517 17279 8551
rect 17221 8511 17279 8517
rect 18230 8508 18236 8560
rect 18288 8548 18294 8560
rect 19518 8548 19524 8560
rect 18288 8520 19524 8548
rect 18288 8508 18294 8520
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 2406 8440 2412 8492
rect 2464 8480 2470 8492
rect 7006 8480 7012 8492
rect 2464 8452 7012 8480
rect 2464 8440 2470 8452
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 7742 8440 7748 8492
rect 7800 8480 7806 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 7800 8452 8493 8480
rect 7800 8440 7806 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 10045 8483 10103 8489
rect 10045 8480 10057 8483
rect 8481 8443 8539 8449
rect 8588 8452 10057 8480
rect 7650 8372 7656 8424
rect 7708 8412 7714 8424
rect 8588 8412 8616 8452
rect 10045 8449 10057 8452
rect 10091 8449 10103 8483
rect 14200 8480 14228 8508
rect 14200 8452 15148 8480
rect 10045 8443 10103 8449
rect 9858 8412 9864 8424
rect 7708 8384 8616 8412
rect 9819 8384 9864 8412
rect 7708 8372 7714 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 11241 8415 11299 8421
rect 11241 8412 11253 8415
rect 10376 8384 11253 8412
rect 10376 8372 10382 8384
rect 11241 8381 11253 8384
rect 11287 8412 11299 8415
rect 11882 8412 11888 8424
rect 11287 8384 11888 8412
rect 11287 8381 11299 8384
rect 11241 8375 11299 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 15013 8415 15071 8421
rect 15013 8412 15025 8415
rect 12851 8384 15025 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 15013 8381 15025 8384
rect 15059 8381 15071 8415
rect 15120 8412 15148 8452
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 18601 8483 18659 8489
rect 18601 8480 18613 8483
rect 16356 8452 18613 8480
rect 16356 8440 16362 8452
rect 18601 8449 18613 8452
rect 18647 8449 18659 8483
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 18601 8443 18659 8449
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 20622 8440 20628 8492
rect 20680 8480 20686 8492
rect 20680 8452 20725 8480
rect 20680 8440 20686 8452
rect 15269 8415 15327 8421
rect 15269 8412 15281 8415
rect 15120 8384 15281 8412
rect 15013 8375 15071 8381
rect 15269 8381 15281 8384
rect 15315 8381 15327 8415
rect 15269 8375 15327 8381
rect 4709 8347 4767 8353
rect 4709 8313 4721 8347
rect 4755 8344 4767 8347
rect 5626 8344 5632 8356
rect 4755 8316 5632 8344
rect 4755 8313 4767 8316
rect 4709 8307 4767 8313
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 8202 8344 8208 8356
rect 5767 8316 8208 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 8202 8304 8208 8316
rect 8260 8304 8266 8356
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 13050 8347 13108 8353
rect 13050 8344 13062 8347
rect 12124 8316 13062 8344
rect 12124 8304 12130 8316
rect 13050 8313 13062 8316
rect 13096 8313 13108 8347
rect 15028 8344 15056 8375
rect 15654 8372 15660 8424
rect 15712 8412 15718 8424
rect 17218 8412 17224 8424
rect 15712 8384 17224 8412
rect 15712 8372 15718 8384
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 17402 8412 17408 8424
rect 17363 8384 17408 8412
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 18138 8372 18144 8424
rect 18196 8412 18202 8424
rect 18417 8415 18475 8421
rect 18417 8412 18429 8415
rect 18196 8384 18429 8412
rect 18196 8372 18202 8384
rect 18417 8381 18429 8384
rect 18463 8381 18475 8415
rect 18417 8375 18475 8381
rect 16758 8344 16764 8356
rect 15028 8316 16764 8344
rect 13050 8307 13108 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 18509 8347 18567 8353
rect 18509 8313 18521 8347
rect 18555 8344 18567 8347
rect 18598 8344 18604 8356
rect 18555 8316 18604 8344
rect 18555 8313 18567 8316
rect 18509 8307 18567 8313
rect 18598 8304 18604 8316
rect 18656 8304 18662 8356
rect 19886 8344 19892 8356
rect 19847 8316 19892 8344
rect 19886 8304 19892 8316
rect 19944 8344 19950 8356
rect 20441 8347 20499 8353
rect 20441 8344 20453 8347
rect 19944 8316 20453 8344
rect 19944 8304 19950 8316
rect 20441 8313 20453 8316
rect 20487 8313 20499 8347
rect 20441 8307 20499 8313
rect 6914 8276 6920 8288
rect 6875 8248 6920 8276
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 8294 8276 8300 8288
rect 8255 8248 8300 8276
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 8389 8279 8447 8285
rect 8389 8245 8401 8279
rect 8435 8276 8447 8279
rect 9493 8279 9551 8285
rect 9493 8276 9505 8279
rect 8435 8248 9505 8276
rect 8435 8245 8447 8248
rect 8389 8239 8447 8245
rect 9493 8245 9505 8248
rect 9539 8245 9551 8279
rect 9493 8239 9551 8245
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10686 8276 10692 8288
rect 9999 8248 10692 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 17494 8276 17500 8288
rect 10836 8248 17500 8276
rect 10836 8236 10842 8248
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 18046 8276 18052 8288
rect 18007 8248 18052 8276
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 20070 8276 20076 8288
rect 20031 8248 20076 8276
rect 20070 8236 20076 8248
rect 20128 8236 20134 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 4430 8072 4436 8084
rect 4391 8044 4436 8072
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 6825 8075 6883 8081
rect 6825 8041 6837 8075
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 6638 8004 6644 8016
rect 5460 7976 6644 8004
rect 5460 7945 5488 7976
rect 6638 7964 6644 7976
rect 6696 7964 6702 8016
rect 6840 8004 6868 8035
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 6972 8044 8033 8072
rect 6972 8032 6978 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8478 8032 8484 8084
rect 8536 8072 8542 8084
rect 9030 8072 9036 8084
rect 8536 8044 9036 8072
rect 8536 8032 8542 8044
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 9180 8044 9229 8072
rect 9180 8032 9186 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10042 8072 10048 8084
rect 9916 8044 10048 8072
rect 9916 8032 9922 8044
rect 10042 8032 10048 8044
rect 10100 8032 10106 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 12483 8044 13553 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13909 8075 13967 8081
rect 13909 8041 13921 8075
rect 13955 8072 13967 8075
rect 18046 8072 18052 8084
rect 13955 8044 18052 8072
rect 13955 8041 13967 8044
rect 13909 8035 13967 8041
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19242 8072 19248 8084
rect 18831 8044 19248 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 6840 7976 7696 8004
rect 7668 7948 7696 7976
rect 8202 7964 8208 8016
rect 8260 8004 8266 8016
rect 15933 8007 15991 8013
rect 15933 8004 15945 8007
rect 8260 7976 15945 8004
rect 8260 7964 8266 7976
rect 15933 7973 15945 7976
rect 15979 7973 15991 8007
rect 15933 7967 15991 7973
rect 16022 7964 16028 8016
rect 16080 8004 16086 8016
rect 16080 7976 16125 8004
rect 16080 7964 16086 7976
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 19153 8007 19211 8013
rect 19153 8004 19165 8007
rect 18012 7976 19165 8004
rect 18012 7964 18018 7976
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5712 7939 5770 7945
rect 5712 7905 5724 7939
rect 5758 7936 5770 7939
rect 6914 7936 6920 7948
rect 5758 7908 6920 7936
rect 5758 7905 5770 7908
rect 5712 7899 5770 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7650 7896 7656 7948
rect 7708 7936 7714 7948
rect 7708 7908 8248 7936
rect 7708 7896 7714 7908
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 8220 7877 8248 7908
rect 8570 7896 8576 7948
rect 8628 7936 8634 7948
rect 10042 7945 10048 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 8628 7908 9413 7936
rect 8628 7896 8634 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 10036 7936 10048 7945
rect 10003 7908 10048 7936
rect 9401 7899 9459 7905
rect 10036 7899 10048 7908
rect 10042 7896 10048 7899
rect 10100 7896 10106 7948
rect 12342 7936 12348 7948
rect 12303 7908 12348 7936
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 17586 7936 17592 7948
rect 17499 7908 17592 7936
rect 17586 7896 17592 7908
rect 17644 7936 17650 7948
rect 18690 7936 18696 7948
rect 17644 7908 18696 7936
rect 17644 7896 17650 7908
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 8113 7871 8171 7877
rect 8113 7868 8125 7871
rect 7800 7840 8125 7868
rect 7800 7828 7806 7840
rect 8113 7837 8125 7840
rect 8159 7837 8171 7871
rect 8113 7831 8171 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 9122 7868 9128 7880
rect 8536 7840 9128 7868
rect 8536 7828 8542 7840
rect 9122 7828 9128 7840
rect 9180 7868 9186 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9180 7840 9781 7868
rect 9180 7828 9186 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12124 7840 12541 7868
rect 12124 7828 12130 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 14001 7871 14059 7877
rect 14001 7868 14013 7871
rect 13228 7840 14013 7868
rect 13228 7828 13234 7840
rect 14001 7837 14013 7840
rect 14047 7837 14059 7871
rect 14001 7831 14059 7837
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14148 7840 14193 7868
rect 14148 7828 14154 7840
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 17678 7868 17684 7880
rect 16172 7840 16217 7868
rect 17639 7840 17684 7868
rect 16172 7828 16178 7840
rect 17678 7828 17684 7840
rect 17736 7828 17742 7880
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 17828 7840 17873 7868
rect 17828 7828 17834 7840
rect 7653 7803 7711 7809
rect 7653 7769 7665 7803
rect 7699 7800 7711 7803
rect 8294 7800 8300 7812
rect 7699 7772 8300 7800
rect 7699 7769 7711 7772
rect 7653 7763 7711 7769
rect 8294 7760 8300 7772
rect 8352 7760 8358 7812
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 14642 7800 14648 7812
rect 11112 7772 14648 7800
rect 11112 7760 11118 7772
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 18322 7800 18328 7812
rect 15712 7772 18328 7800
rect 15712 7760 15718 7772
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 4338 7692 4344 7744
rect 4396 7732 4402 7744
rect 9398 7732 9404 7744
rect 4396 7704 9404 7732
rect 4396 7692 4402 7704
rect 9398 7692 9404 7704
rect 9456 7692 9462 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11238 7732 11244 7744
rect 11195 7704 11244 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11238 7692 11244 7704
rect 11296 7732 11302 7744
rect 11698 7732 11704 7744
rect 11296 7704 11704 7732
rect 11296 7692 11302 7704
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 11940 7704 11989 7732
rect 11940 7692 11946 7704
rect 11977 7701 11989 7704
rect 12023 7701 12035 7735
rect 11977 7695 12035 7701
rect 15565 7735 15623 7741
rect 15565 7701 15577 7735
rect 15611 7732 15623 7735
rect 15930 7732 15936 7744
rect 15611 7704 15936 7732
rect 15611 7701 15623 7704
rect 15565 7695 15623 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 17221 7735 17279 7741
rect 17221 7701 17233 7735
rect 17267 7732 17279 7735
rect 17954 7732 17960 7744
rect 17267 7704 17960 7732
rect 17267 7701 17279 7704
rect 17221 7695 17279 7701
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 19076 7732 19104 7976
rect 19153 7973 19165 7976
rect 19199 7973 19211 8007
rect 19153 7967 19211 7973
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19337 7871 19395 7877
rect 19337 7837 19349 7871
rect 19383 7837 19395 7871
rect 19337 7831 19395 7837
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 19352 7800 19380 7831
rect 19208 7772 19380 7800
rect 19208 7760 19214 7772
rect 19242 7732 19248 7744
rect 19076 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 5442 7528 5448 7540
rect 3200 7500 5448 7528
rect 3200 7488 3206 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 6457 7531 6515 7537
rect 6457 7497 6469 7531
rect 6503 7528 6515 7531
rect 6638 7528 6644 7540
rect 6503 7500 6644 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 12437 7531 12495 7537
rect 12437 7528 12449 7531
rect 12400 7500 12449 7528
rect 12400 7488 12406 7500
rect 12437 7497 12449 7500
rect 12483 7497 12495 7531
rect 12437 7491 12495 7497
rect 12986 7488 12992 7540
rect 13044 7528 13050 7540
rect 13044 7500 19104 7528
rect 13044 7488 13050 7500
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 9861 7463 9919 7469
rect 5684 7432 8524 7460
rect 5684 7420 5690 7432
rect 7006 7392 7012 7404
rect 6967 7364 7012 7392
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 8496 7392 8524 7432
rect 9861 7429 9873 7463
rect 9907 7460 9919 7463
rect 10042 7460 10048 7472
rect 9907 7432 10048 7460
rect 9907 7429 9919 7432
rect 9861 7423 9919 7429
rect 10042 7420 10048 7432
rect 10100 7460 10106 7472
rect 12618 7460 12624 7472
rect 10100 7432 12624 7460
rect 10100 7420 10106 7432
rect 12618 7420 12624 7432
rect 12676 7460 12682 7472
rect 16298 7460 16304 7472
rect 12676 7432 16304 7460
rect 12676 7420 12682 7432
rect 8496 7364 8616 7392
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 5166 7324 5172 7336
rect 3007 7296 3372 7324
rect 5127 7296 5172 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 3344 7268 3372 7296
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5442 7324 5448 7336
rect 5403 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7293 6699 7327
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6641 7287 6699 7293
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3206 7259 3264 7265
rect 3206 7256 3218 7259
rect 3108 7228 3218 7256
rect 3108 7216 3114 7228
rect 3206 7225 3218 7228
rect 3252 7225 3264 7259
rect 3206 7219 3264 7225
rect 3326 7216 3332 7268
rect 3384 7216 3390 7268
rect 6656 7256 6684 7287
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8588 7324 8616 7364
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11241 7395 11299 7401
rect 11241 7392 11253 7395
rect 11112 7364 11253 7392
rect 11112 7352 11118 7364
rect 11241 7361 11253 7364
rect 11287 7361 11299 7395
rect 11241 7355 11299 7361
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 11756 7364 13093 7392
rect 11756 7352 11762 7364
rect 13081 7361 13093 7364
rect 13127 7392 13139 7395
rect 14090 7392 14096 7404
rect 13127 7364 14096 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14660 7401 14688 7432
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 19076 7460 19104 7500
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19429 7531 19487 7537
rect 19429 7528 19441 7531
rect 19208 7500 19441 7528
rect 19208 7488 19214 7500
rect 19429 7497 19441 7500
rect 19475 7497 19487 7531
rect 19429 7491 19487 7497
rect 19334 7460 19340 7472
rect 19076 7432 19340 7460
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 14645 7395 14703 7401
rect 14645 7361 14657 7395
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15344 7364 16037 7392
rect 15344 7352 15350 7364
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 16482 7392 16488 7404
rect 16255 7364 16488 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 16482 7352 16488 7364
rect 16540 7352 16546 7404
rect 18046 7392 18052 7404
rect 18007 7364 18052 7392
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 12805 7327 12863 7333
rect 12805 7324 12817 7327
rect 8588 7296 12817 7324
rect 12805 7293 12817 7296
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 14056 7296 14381 7324
rect 14056 7284 14062 7296
rect 14369 7293 14381 7296
rect 14415 7293 14427 7327
rect 15930 7324 15936 7336
rect 15891 7296 15936 7324
rect 14369 7287 14427 7293
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20530 7324 20536 7336
rect 20036 7296 20536 7324
rect 20036 7284 20042 7296
rect 20530 7284 20536 7296
rect 20588 7284 20594 7336
rect 8570 7256 8576 7268
rect 4356 7228 6592 7256
rect 6656 7228 8576 7256
rect 4356 7197 4384 7228
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7157 4399 7191
rect 6564 7188 6592 7228
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 8754 7265 8760 7268
rect 8748 7219 8760 7265
rect 8812 7256 8818 7268
rect 11057 7259 11115 7265
rect 8812 7228 8848 7256
rect 8754 7216 8760 7219
rect 8812 7216 8818 7228
rect 11057 7225 11069 7259
rect 11103 7256 11115 7259
rect 17678 7256 17684 7268
rect 11103 7228 17684 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 17678 7216 17684 7228
rect 17736 7216 17742 7268
rect 18316 7259 18374 7265
rect 18316 7225 18328 7259
rect 18362 7256 18374 7259
rect 19058 7256 19064 7268
rect 18362 7228 19064 7256
rect 18362 7225 18374 7228
rect 18316 7219 18374 7225
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 6914 7188 6920 7200
rect 6564 7160 6920 7188
rect 4341 7151 4399 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 8720 7160 11161 7188
rect 8720 7148 8726 7160
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11149 7151 11207 7157
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 12802 7188 12808 7200
rect 11296 7160 12808 7188
rect 11296 7148 11302 7160
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 14001 7191 14059 7197
rect 14001 7188 14013 7191
rect 12943 7160 14013 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 14001 7157 14013 7160
rect 14047 7157 14059 7191
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 14001 7151 14059 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 21542 7188 21548 7200
rect 20763 7160 21548 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 21542 7148 21548 7160
rect 21600 7148 21606 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 5997 6987 6055 6993
rect 5997 6953 6009 6987
rect 6043 6984 6055 6987
rect 6822 6984 6828 6996
rect 6043 6956 6828 6984
rect 6043 6953 6055 6956
rect 5997 6947 6055 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 7742 6984 7748 6996
rect 7703 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 10873 6987 10931 6993
rect 10873 6953 10885 6987
rect 10919 6984 10931 6987
rect 11238 6984 11244 6996
rect 10919 6956 11244 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 13170 6984 13176 6996
rect 12115 6956 13176 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 14093 6987 14151 6993
rect 14093 6953 14105 6987
rect 14139 6984 14151 6987
rect 14274 6984 14280 6996
rect 14139 6956 14280 6984
rect 14139 6953 14151 6956
rect 14093 6947 14151 6953
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 7558 6876 7564 6928
rect 7616 6916 7622 6928
rect 8113 6919 8171 6925
rect 8113 6916 8125 6919
rect 7616 6888 8125 6916
rect 7616 6876 7622 6888
rect 8113 6885 8125 6888
rect 8159 6885 8171 6919
rect 11054 6916 11060 6928
rect 8113 6879 8171 6885
rect 8404 6888 11060 6916
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6848 5043 6851
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 5031 6820 6377 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 6365 6817 6377 6820
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 8404 6848 8432 6888
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 12342 6916 12348 6928
rect 11204 6888 12348 6916
rect 11204 6876 11210 6888
rect 12342 6876 12348 6888
rect 12400 6916 12406 6928
rect 12437 6919 12495 6925
rect 12437 6916 12449 6919
rect 12400 6888 12449 6916
rect 12400 6876 12406 6888
rect 12437 6885 12449 6888
rect 12483 6885 12495 6919
rect 12437 6879 12495 6885
rect 12802 6876 12808 6928
rect 12860 6916 12866 6928
rect 13078 6916 13084 6928
rect 12860 6888 13084 6916
rect 12860 6876 12866 6888
rect 13078 6876 13084 6888
rect 13136 6916 13142 6928
rect 13722 6916 13728 6928
rect 13136 6888 13728 6916
rect 13136 6876 13142 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 13998 6916 14004 6928
rect 13959 6888 14004 6916
rect 13998 6876 14004 6888
rect 14056 6876 14062 6928
rect 15556 6919 15614 6925
rect 15556 6885 15568 6919
rect 15602 6916 15614 6919
rect 16114 6916 16120 6928
rect 15602 6888 16120 6916
rect 15602 6885 15614 6888
rect 15556 6879 15614 6885
rect 16114 6876 16120 6888
rect 16172 6876 16178 6928
rect 18046 6916 18052 6928
rect 17696 6888 18052 6916
rect 6972 6820 8432 6848
rect 6972 6808 6978 6820
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 5776 6752 6469 6780
rect 5776 6740 5782 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6780 6699 6783
rect 7650 6780 7656 6792
rect 6687 6752 7656 6780
rect 6687 6749 6699 6752
rect 6641 6743 6699 6749
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 8404 6789 8432 6820
rect 10870 6808 10876 6860
rect 10928 6848 10934 6860
rect 10928 6820 13952 6848
rect 10928 6808 10934 6820
rect 8205 6783 8263 6789
rect 8205 6749 8217 6783
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8389 6783 8447 6789
rect 8389 6749 8401 6783
rect 8435 6749 8447 6783
rect 8389 6743 8447 6749
rect 1946 6672 1952 6724
rect 2004 6712 2010 6724
rect 2498 6712 2504 6724
rect 2004 6684 2504 6712
rect 2004 6672 2010 6684
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 8220 6712 8248 6743
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 11072 6789 11100 6820
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 8536 6752 10977 6780
rect 8536 6740 8542 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 10965 6743 11023 6749
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11146 6740 11152 6792
rect 11204 6780 11210 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 11204 6752 12541 6780
rect 11204 6740 11210 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 12618 6740 12624 6792
rect 12676 6780 12682 6792
rect 12676 6752 12721 6780
rect 12676 6740 12682 6752
rect 10502 6712 10508 6724
rect 2556 6684 8248 6712
rect 10463 6684 10508 6712
rect 2556 6672 2562 6684
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 12768 6684 13645 6712
rect 12768 6672 12774 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13924 6712 13952 6820
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 15252 6820 15301 6848
rect 15252 6808 15258 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 16758 6848 16764 6860
rect 15335 6820 16764 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 16758 6808 16764 6820
rect 16816 6808 16822 6860
rect 17696 6857 17724 6888
rect 18046 6876 18052 6888
rect 18104 6916 18110 6928
rect 18690 6916 18696 6928
rect 18104 6888 18696 6916
rect 18104 6876 18110 6888
rect 18690 6876 18696 6888
rect 18748 6876 18754 6928
rect 17681 6851 17739 6857
rect 17681 6817 17693 6851
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 17948 6851 18006 6857
rect 17948 6817 17960 6851
rect 17994 6848 18006 6851
rect 20622 6848 20628 6860
rect 17994 6820 20628 6848
rect 17994 6817 18006 6820
rect 17948 6811 18006 6817
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 14274 6780 14280 6792
rect 14235 6752 14280 6780
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14292 6712 14320 6740
rect 17126 6712 17132 6724
rect 13924 6684 14320 6712
rect 16408 6684 17132 6712
rect 13633 6675 13691 6681
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 3694 6644 3700 6656
rect 2740 6616 3700 6644
rect 2740 6604 2746 6616
rect 3694 6604 3700 6616
rect 3752 6644 3758 6656
rect 11146 6644 11152 6656
rect 3752 6616 11152 6644
rect 3752 6604 3758 6616
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 16408 6644 16436 6684
rect 17126 6672 17132 6684
rect 17184 6712 17190 6724
rect 17586 6712 17592 6724
rect 17184 6684 17592 6712
rect 17184 6672 17190 6684
rect 17586 6672 17592 6684
rect 17644 6672 17650 6724
rect 14240 6616 16436 6644
rect 14240 6604 14246 6616
rect 16482 6604 16488 6656
rect 16540 6644 16546 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16540 6616 16681 6644
rect 16540 6604 16546 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 19058 6644 19064 6656
rect 19019 6616 19064 6644
rect 16669 6607 16727 6613
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 5166 6440 5172 6452
rect 3835 6412 5172 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 14182 6440 14188 6452
rect 8996 6412 14188 6440
rect 8996 6400 9002 6412
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 14274 6400 14280 6452
rect 14332 6440 14338 6452
rect 16577 6443 16635 6449
rect 16577 6440 16589 6443
rect 14332 6412 16589 6440
rect 14332 6400 14338 6412
rect 16577 6409 16589 6412
rect 16623 6409 16635 6443
rect 16577 6403 16635 6409
rect 10689 6375 10747 6381
rect 10689 6341 10701 6375
rect 10735 6372 10747 6375
rect 12434 6372 12440 6384
rect 10735 6344 12440 6372
rect 10735 6341 10747 6344
rect 10689 6335 10747 6341
rect 12434 6332 12440 6344
rect 12492 6372 12498 6384
rect 12492 6344 13032 6372
rect 12492 6332 12498 6344
rect 4338 6304 4344 6316
rect 4299 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6638 6304 6644 6316
rect 6328 6276 6644 6304
rect 6328 6264 6334 6276
rect 6638 6264 6644 6276
rect 6696 6304 6702 6316
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6696 6276 6837 6304
rect 6696 6264 6702 6276
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 9180 6276 9321 6304
rect 9180 6264 9186 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 10502 6264 10508 6316
rect 10560 6304 10566 6316
rect 13004 6313 13032 6344
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 10560 6276 12909 6304
rect 10560 6264 10566 6276
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6273 13047 6307
rect 14458 6304 14464 6316
rect 12989 6267 13047 6273
rect 14016 6276 14464 6304
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 9214 6236 9220 6248
rect 2823 6208 6776 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 6748 6168 6776 6208
rect 7024 6208 9220 6236
rect 7024 6168 7052 6208
rect 9214 6196 9220 6208
rect 9272 6196 9278 6248
rect 9576 6239 9634 6245
rect 9576 6205 9588 6239
rect 9622 6236 9634 6239
rect 10870 6236 10876 6248
rect 9622 6208 10876 6236
rect 9622 6205 9634 6208
rect 9576 6199 9634 6205
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 14016 6236 14044 6276
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 15194 6304 15200 6316
rect 15155 6276 15200 6304
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 17586 6264 17592 6316
rect 17644 6304 17650 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 17644 6276 18613 6304
rect 17644 6264 17650 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6304 18843 6307
rect 19886 6304 19892 6316
rect 18831 6276 19892 6304
rect 18831 6273 18843 6276
rect 18785 6267 18843 6273
rect 19886 6264 19892 6276
rect 19944 6264 19950 6316
rect 20349 6307 20407 6313
rect 20349 6273 20361 6307
rect 20395 6304 20407 6307
rect 20622 6304 20628 6316
rect 20395 6276 20628 6304
rect 20395 6273 20407 6276
rect 20349 6267 20407 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 11164 6208 14044 6236
rect 14093 6239 14151 6245
rect 6748 6140 7052 6168
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 7650 6168 7656 6180
rect 7138 6140 7656 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 7650 6128 7656 6140
rect 7708 6128 7714 6180
rect 8294 6128 8300 6180
rect 8352 6168 8358 6180
rect 11164 6168 11192 6208
rect 14093 6205 14105 6239
rect 14139 6205 14151 6239
rect 14093 6199 14151 6205
rect 13906 6168 13912 6180
rect 8352 6140 11192 6168
rect 11256 6140 13912 6168
rect 8352 6128 8358 6140
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 4157 6103 4215 6109
rect 4157 6100 4169 6103
rect 3016 6072 4169 6100
rect 3016 6060 3022 6072
rect 4157 6069 4169 6072
rect 4203 6069 4215 6103
rect 4157 6063 4215 6069
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4798 6100 4804 6112
rect 4295 6072 4804 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 5721 6103 5779 6109
rect 5721 6069 5733 6103
rect 5767 6100 5779 6103
rect 7742 6100 7748 6112
rect 5767 6072 7748 6100
rect 5767 6069 5779 6072
rect 5721 6063 5779 6069
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 8202 6100 8208 6112
rect 8163 6072 8208 6100
rect 8202 6060 8208 6072
rect 8260 6060 8266 6112
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 11256 6100 11284 6140
rect 13906 6128 13912 6140
rect 13964 6128 13970 6180
rect 14108 6168 14136 6199
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 14366 6236 14372 6248
rect 14240 6208 14372 6236
rect 14240 6196 14246 6208
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 15464 6239 15522 6245
rect 15464 6205 15476 6239
rect 15510 6236 15522 6239
rect 16482 6236 16488 6248
rect 15510 6208 16488 6236
rect 15510 6205 15522 6208
rect 15464 6199 15522 6205
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 18509 6239 18567 6245
rect 18509 6236 18521 6239
rect 17552 6208 18521 6236
rect 17552 6196 17558 6208
rect 18509 6205 18521 6208
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 16850 6168 16856 6180
rect 14108 6140 16856 6168
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 20165 6171 20223 6177
rect 20165 6168 20177 6171
rect 18156 6140 20177 6168
rect 8444 6072 11284 6100
rect 8444 6060 8450 6072
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12124 6072 12449 6100
rect 12124 6060 12130 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 12802 6100 12808 6112
rect 12763 6072 12808 6100
rect 12437 6063 12495 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 16482 6100 16488 6112
rect 14323 6072 16488 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 18156 6109 18184 6140
rect 20165 6137 20177 6140
rect 20211 6137 20223 6171
rect 20165 6131 20223 6137
rect 18141 6103 18199 6109
rect 18141 6069 18153 6103
rect 18187 6069 18199 6103
rect 19702 6100 19708 6112
rect 19663 6072 19708 6100
rect 18141 6063 18199 6069
rect 19702 6060 19708 6072
rect 19760 6060 19766 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20073 6103 20131 6109
rect 20073 6100 20085 6103
rect 19852 6072 20085 6100
rect 19852 6060 19858 6072
rect 20073 6069 20085 6072
rect 20119 6069 20131 6103
rect 20073 6063 20131 6069
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2958 5896 2964 5908
rect 2919 5868 2964 5896
rect 2958 5856 2964 5868
rect 3016 5856 3022 5908
rect 7650 5896 7656 5908
rect 7611 5868 7656 5896
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 1949 5831 2007 5837
rect 1949 5828 1961 5831
rect 1903 5800 1961 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 1949 5797 1961 5800
rect 1995 5828 2007 5831
rect 1995 5800 5304 5828
rect 1995 5797 2007 5800
rect 1949 5791 2007 5797
rect 4338 5769 4344 5772
rect 4332 5760 4344 5769
rect 4299 5732 4344 5760
rect 4332 5723 4344 5732
rect 4338 5720 4344 5723
rect 4396 5720 4402 5772
rect 5276 5760 5304 5800
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 6518 5831 6576 5837
rect 6518 5828 6530 5831
rect 5500 5800 6530 5828
rect 5500 5788 5506 5800
rect 6518 5797 6530 5800
rect 6564 5797 6576 5831
rect 8680 5828 8708 5859
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 9272 5868 12265 5896
rect 9272 5856 9278 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 12345 5899 12403 5905
rect 12345 5865 12357 5899
rect 12391 5896 12403 5899
rect 12710 5896 12716 5908
rect 12391 5868 12716 5896
rect 12391 5865 12403 5868
rect 12345 5859 12403 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13449 5899 13507 5905
rect 13449 5896 13461 5899
rect 12860 5868 13461 5896
rect 12860 5856 12866 5868
rect 13449 5865 13461 5868
rect 13495 5865 13507 5899
rect 13449 5859 13507 5865
rect 13817 5899 13875 5905
rect 13817 5865 13829 5899
rect 13863 5896 13875 5899
rect 14734 5896 14740 5908
rect 13863 5868 14740 5896
rect 13863 5865 13875 5868
rect 13817 5859 13875 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 19794 5896 19800 5908
rect 19291 5868 19800 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 14366 5828 14372 5840
rect 8680 5800 14372 5828
rect 6518 5791 6576 5797
rect 14366 5788 14372 5800
rect 14424 5788 14430 5840
rect 17028 5831 17086 5837
rect 17028 5797 17040 5831
rect 17074 5828 17086 5831
rect 17770 5828 17776 5840
rect 17074 5800 17776 5828
rect 17074 5797 17086 5800
rect 17028 5791 17086 5797
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 18874 5788 18880 5840
rect 18932 5828 18938 5840
rect 19613 5831 19671 5837
rect 19613 5828 19625 5831
rect 18932 5800 19625 5828
rect 18932 5788 18938 5800
rect 19613 5797 19625 5800
rect 19659 5797 19671 5831
rect 19613 5791 19671 5797
rect 8294 5760 8300 5772
rect 5276 5732 8300 5760
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8478 5760 8484 5772
rect 8439 5732 8484 5760
rect 8478 5720 8484 5732
rect 8536 5720 8542 5772
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9674 5760 9680 5772
rect 9180 5732 9680 5760
rect 9180 5720 9186 5732
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 9990 5732 11192 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 6270 5692 6276 5704
rect 6231 5664 6276 5692
rect 4065 5655 4123 5661
rect 3142 5516 3148 5568
rect 3200 5556 3206 5568
rect 3326 5556 3332 5568
rect 3200 5528 3332 5556
rect 3200 5516 3206 5528
rect 3326 5516 3332 5528
rect 3384 5556 3390 5568
rect 4080 5556 4108 5655
rect 6270 5652 6276 5664
rect 6328 5652 6334 5704
rect 11164 5692 11192 5732
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 14608 5732 15669 5760
rect 14608 5720 14614 5732
rect 15657 5729 15669 5732
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 12434 5692 12440 5704
rect 11164 5664 12440 5692
rect 12434 5652 12440 5664
rect 12492 5692 12498 5704
rect 13906 5692 13912 5704
rect 12492 5664 12585 5692
rect 13867 5664 13912 5692
rect 12492 5652 12498 5664
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 14274 5692 14280 5704
rect 14139 5664 14280 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 16758 5652 16764 5704
rect 16816 5692 16822 5704
rect 16816 5664 16861 5692
rect 16816 5652 16822 5664
rect 18138 5652 18144 5704
rect 18196 5692 18202 5704
rect 19705 5695 19763 5701
rect 19705 5692 19717 5695
rect 18196 5664 19717 5692
rect 18196 5652 18202 5664
rect 19705 5661 19717 5664
rect 19751 5661 19763 5695
rect 19886 5692 19892 5704
rect 19847 5664 19892 5692
rect 19705 5655 19763 5661
rect 5442 5624 5448 5636
rect 5403 5596 5448 5624
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 19610 5624 19616 5636
rect 17972 5596 19616 5624
rect 6270 5556 6276 5568
rect 3384 5528 6276 5556
rect 3384 5516 3390 5528
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 11054 5556 11060 5568
rect 11015 5528 11060 5556
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11885 5559 11943 5565
rect 11885 5556 11897 5559
rect 11204 5528 11897 5556
rect 11204 5516 11210 5528
rect 11885 5525 11897 5528
rect 11931 5525 11943 5559
rect 11885 5519 11943 5525
rect 15841 5559 15899 5565
rect 15841 5525 15853 5559
rect 15887 5556 15899 5559
rect 17972 5556 18000 5596
rect 19610 5584 19616 5596
rect 19668 5584 19674 5636
rect 19720 5624 19748 5655
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 19978 5624 19984 5636
rect 19720 5596 19984 5624
rect 19978 5584 19984 5596
rect 20036 5584 20042 5636
rect 18138 5556 18144 5568
rect 15887 5528 18000 5556
rect 18099 5528 18144 5556
rect 15887 5525 15899 5528
rect 15841 5519 15899 5525
rect 18138 5516 18144 5528
rect 18196 5516 18202 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 4154 5352 4160 5364
rect 3384 5324 4160 5352
rect 3384 5312 3390 5324
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4338 5312 4344 5364
rect 4396 5352 4402 5364
rect 4525 5355 4583 5361
rect 4525 5352 4537 5355
rect 4396 5324 4537 5352
rect 4396 5312 4402 5324
rect 4525 5321 4537 5324
rect 4571 5321 4583 5355
rect 8754 5352 8760 5364
rect 8715 5324 8760 5352
rect 4525 5315 4583 5321
rect 8754 5312 8760 5324
rect 8812 5312 8818 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 18046 5352 18052 5364
rect 13964 5324 18052 5352
rect 13964 5312 13970 5324
rect 18046 5312 18052 5324
rect 18104 5312 18110 5364
rect 20438 5352 20444 5364
rect 19444 5324 20444 5352
rect 4890 5244 4896 5296
rect 4948 5284 4954 5296
rect 5350 5284 5356 5296
rect 4948 5256 5356 5284
rect 4948 5244 4954 5256
rect 5350 5244 5356 5256
rect 5408 5244 5414 5296
rect 12805 5287 12863 5293
rect 12805 5253 12817 5287
rect 12851 5284 12863 5287
rect 14550 5284 14556 5296
rect 12851 5256 14556 5284
rect 12851 5253 12863 5256
rect 12805 5247 12863 5253
rect 14550 5244 14556 5256
rect 14608 5244 14614 5296
rect 17037 5287 17095 5293
rect 17037 5253 17049 5287
rect 17083 5284 17095 5287
rect 19444 5284 19472 5324
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 20622 5312 20628 5364
rect 20680 5352 20686 5364
rect 20809 5355 20867 5361
rect 20809 5352 20821 5355
rect 20680 5324 20821 5352
rect 20680 5312 20686 5324
rect 20809 5321 20821 5324
rect 20855 5321 20867 5355
rect 20809 5315 20867 5321
rect 17083 5256 19472 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 3142 5216 3148 5228
rect 3103 5188 3148 5216
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6730 5216 6736 5228
rect 6328 5188 6736 5216
rect 6328 5176 6334 5188
rect 6730 5176 6736 5188
rect 6788 5216 6794 5228
rect 7377 5219 7435 5225
rect 7377 5216 7389 5219
rect 6788 5188 7389 5216
rect 6788 5176 6794 5188
rect 7377 5185 7389 5188
rect 7423 5185 7435 5219
rect 7377 5179 7435 5185
rect 8662 5176 8668 5228
rect 8720 5216 8726 5228
rect 9030 5216 9036 5228
rect 8720 5188 9036 5216
rect 8720 5176 8726 5188
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11112 5188 11345 5216
rect 11112 5176 11118 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 14182 5216 14188 5228
rect 14143 5188 14188 5216
rect 11333 5179 11391 5185
rect 14182 5176 14188 5188
rect 14240 5176 14246 5228
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 14332 5188 15853 5216
rect 14332 5176 14338 5188
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 18690 5176 18696 5228
rect 18748 5216 18754 5228
rect 19429 5219 19487 5225
rect 19429 5216 19441 5219
rect 18748 5188 19441 5216
rect 18748 5176 18754 5188
rect 19429 5185 19441 5188
rect 19475 5185 19487 5219
rect 19429 5179 19487 5185
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 5629 5111 5687 5117
rect 3412 5083 3470 5089
rect 3412 5049 3424 5083
rect 3458 5080 3470 5083
rect 4154 5080 4160 5092
rect 3458 5052 4160 5080
rect 3458 5049 3470 5052
rect 3412 5043 3470 5049
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 5644 5080 5672 5111
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7644 5151 7702 5157
rect 7644 5148 7656 5151
rect 7524 5120 7656 5148
rect 7524 5108 7530 5120
rect 7644 5117 7656 5120
rect 7690 5148 7702 5151
rect 8202 5148 8208 5160
rect 7690 5120 8208 5148
rect 7690 5117 7702 5120
rect 7644 5111 7702 5117
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 9677 5151 9735 5157
rect 9677 5148 9689 5151
rect 9456 5120 9689 5148
rect 9456 5108 9462 5120
rect 9677 5117 9689 5120
rect 9723 5148 9735 5151
rect 10778 5148 10784 5160
rect 9723 5120 10784 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 10778 5108 10784 5120
rect 10836 5108 10842 5160
rect 11146 5148 11152 5160
rect 11107 5120 11152 5148
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 11241 5151 11299 5157
rect 11241 5117 11253 5151
rect 11287 5148 11299 5151
rect 12066 5148 12072 5160
rect 11287 5120 12072 5148
rect 11287 5117 11299 5120
rect 11241 5111 11299 5117
rect 12066 5108 12072 5120
rect 12124 5108 12130 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 12986 5148 12992 5160
rect 12667 5120 12992 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 15654 5148 15660 5160
rect 13780 5120 15516 5148
rect 15615 5120 15660 5148
rect 13780 5108 13786 5120
rect 9030 5080 9036 5092
rect 5644 5052 9036 5080
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 15488 5080 15516 5120
rect 15654 5108 15660 5120
rect 15712 5108 15718 5160
rect 16853 5151 16911 5157
rect 16853 5148 16865 5151
rect 15764 5120 16865 5148
rect 15764 5080 15792 5120
rect 16853 5117 16865 5120
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 18325 5151 18383 5157
rect 18325 5117 18337 5151
rect 18371 5117 18383 5151
rect 18325 5111 18383 5117
rect 10796 5052 11652 5080
rect 15488 5052 15792 5080
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 8202 5012 8208 5024
rect 5859 4984 8208 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 9861 5015 9919 5021
rect 9861 4981 9873 5015
rect 9907 5012 9919 5015
rect 10686 5012 10692 5024
rect 9907 4984 10692 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10796 5021 10824 5052
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 4981 10839 5015
rect 11624 5012 11652 5052
rect 16206 5040 16212 5092
rect 16264 5080 16270 5092
rect 18340 5080 18368 5111
rect 16264 5052 18368 5080
rect 19696 5083 19754 5089
rect 16264 5040 16270 5052
rect 19696 5049 19708 5083
rect 19742 5080 19754 5083
rect 19886 5080 19892 5092
rect 19742 5052 19892 5080
rect 19742 5049 19754 5052
rect 19696 5043 19754 5049
rect 19886 5040 19892 5052
rect 19944 5040 19950 5092
rect 12618 5012 12624 5024
rect 11624 4984 12624 5012
rect 10781 4975 10839 4981
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13906 5012 13912 5024
rect 13771 4984 13912 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 13998 4972 14004 5024
rect 14056 5012 14062 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 14056 4984 14105 5012
rect 14056 4972 14062 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 14332 4984 15301 5012
rect 14332 4972 14338 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 18046 5012 18052 5024
rect 15804 4984 18052 5012
rect 15804 4972 15810 4984
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 5012 18567 5015
rect 20254 5012 20260 5024
rect 18555 4984 20260 5012
rect 18555 4981 18567 4984
rect 18509 4975 18567 4981
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 4798 4808 4804 4820
rect 2455 4780 4804 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 4798 4768 4804 4780
rect 4856 4768 4862 4820
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 5718 4808 5724 4820
rect 4939 4780 5724 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6457 4811 6515 4817
rect 6457 4777 6469 4811
rect 6503 4808 6515 4811
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 6503 4780 8493 4808
rect 6503 4777 6515 4780
rect 6457 4771 6515 4777
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 9030 4768 9036 4820
rect 9088 4808 9094 4820
rect 12253 4811 12311 4817
rect 9088 4780 11284 4808
rect 9088 4768 9094 4780
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 6362 4740 6368 4752
rect 2188 4712 6368 4740
rect 2188 4700 2194 4712
rect 6362 4700 6368 4712
rect 6420 4700 6426 4752
rect 6546 4700 6552 4752
rect 6604 4740 6610 4752
rect 6917 4743 6975 4749
rect 6917 4740 6929 4743
rect 6604 4712 6929 4740
rect 6604 4700 6610 4712
rect 6917 4709 6929 4712
rect 6963 4709 6975 4743
rect 6917 4703 6975 4709
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 8389 4743 8447 4749
rect 8389 4740 8401 4743
rect 7800 4712 8401 4740
rect 7800 4700 7806 4712
rect 8389 4709 8401 4712
rect 8435 4709 8447 4743
rect 8389 4703 8447 4709
rect 11054 4700 11060 4752
rect 11112 4749 11118 4752
rect 11112 4743 11176 4749
rect 11112 4709 11130 4743
rect 11164 4709 11176 4743
rect 11256 4740 11284 4780
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12526 4808 12532 4820
rect 12299 4780 12532 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 15289 4811 15347 4817
rect 15289 4808 15301 4811
rect 14139 4780 15301 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 15289 4777 15301 4780
rect 15335 4777 15347 4811
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15289 4771 15347 4777
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 17313 4811 17371 4817
rect 17313 4808 17325 4811
rect 16264 4780 17325 4808
rect 16264 4768 16270 4780
rect 17313 4777 17325 4780
rect 17359 4777 17371 4811
rect 17313 4771 17371 4777
rect 13814 4740 13820 4752
rect 11256 4712 13820 4740
rect 11112 4703 11176 4709
rect 11112 4700 11118 4703
rect 13814 4700 13820 4712
rect 13872 4700 13878 4752
rect 14001 4743 14059 4749
rect 14001 4709 14013 4743
rect 14047 4740 14059 4743
rect 14274 4740 14280 4752
rect 14047 4712 14280 4740
rect 14047 4709 14059 4712
rect 14001 4703 14059 4709
rect 14274 4700 14280 4712
rect 14332 4700 14338 4752
rect 17405 4743 17463 4749
rect 17405 4740 17417 4743
rect 14936 4712 17417 4740
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 2832 4644 2877 4672
rect 2832 4632 2838 4644
rect 4246 4632 4252 4684
rect 4304 4672 4310 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 4304 4644 5273 4672
rect 4304 4632 4310 4644
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 5261 4635 5319 4641
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 6825 4675 6883 4681
rect 6825 4672 6837 4675
rect 5592 4644 6837 4672
rect 5592 4632 5598 4644
rect 6825 4641 6837 4644
rect 6871 4641 6883 4675
rect 9769 4675 9827 4681
rect 9769 4672 9781 4675
rect 6825 4635 6883 4641
rect 7944 4644 9781 4672
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 4154 4604 4160 4616
rect 3099 4576 4160 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 2884 4536 2912 4567
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 4890 4536 4896 4548
rect 2884 4508 4896 4536
rect 4890 4496 4896 4508
rect 4948 4496 4954 4548
rect 5368 4536 5396 4567
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 7101 4607 7159 4613
rect 5500 4576 5545 4604
rect 5500 4564 5506 4576
rect 7101 4573 7113 4607
rect 7147 4604 7159 4607
rect 7466 4604 7472 4616
rect 7147 4576 7472 4604
rect 7147 4573 7159 4576
rect 7101 4567 7159 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 6914 4536 6920 4548
rect 5368 4508 6920 4536
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 7944 4468 7972 4644
rect 9769 4641 9781 4644
rect 9815 4672 9827 4675
rect 14936 4672 14964 4712
rect 17405 4709 17417 4712
rect 17451 4709 17463 4743
rect 17405 4703 17463 4709
rect 18138 4700 18144 4752
rect 18196 4740 18202 4752
rect 18598 4740 18604 4752
rect 18196 4712 18604 4740
rect 18196 4700 18202 4712
rect 18598 4700 18604 4712
rect 18656 4740 18662 4752
rect 18754 4743 18812 4749
rect 18754 4740 18766 4743
rect 18656 4712 18766 4740
rect 18656 4700 18662 4712
rect 18754 4709 18766 4712
rect 18800 4709 18812 4743
rect 18754 4703 18812 4709
rect 9815 4644 14964 4672
rect 15657 4675 15715 4681
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 15657 4641 15669 4675
rect 15703 4672 15715 4675
rect 20530 4672 20536 4684
rect 15703 4644 20536 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 20530 4632 20536 4644
rect 20588 4632 20594 4684
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 8754 4604 8760 4616
rect 8711 4576 8760 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10873 4607 10931 4613
rect 10873 4604 10885 4607
rect 9732 4576 10885 4604
rect 9732 4564 9738 4576
rect 10873 4573 10885 4576
rect 10919 4573 10931 4607
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 10873 4567 10931 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 15841 4607 15899 4613
rect 15841 4573 15853 4607
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17770 4604 17776 4616
rect 17635 4576 17776 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 8021 4539 8079 4545
rect 8021 4505 8033 4539
rect 8067 4536 8079 4539
rect 9766 4536 9772 4548
rect 8067 4508 9772 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 12526 4496 12532 4548
rect 12584 4536 12590 4548
rect 14182 4536 14188 4548
rect 12584 4508 14188 4536
rect 12584 4496 12590 4508
rect 14182 4496 14188 4508
rect 14240 4536 14246 4548
rect 15856 4536 15884 4567
rect 17770 4564 17776 4576
rect 17828 4564 17834 4616
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 14240 4508 15884 4536
rect 14240 4496 14246 4508
rect 5040 4440 7972 4468
rect 5040 4428 5046 4440
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 9858 4468 9864 4480
rect 8536 4440 9864 4468
rect 8536 4428 8542 4440
rect 9858 4428 9864 4440
rect 9916 4428 9922 4480
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 11146 4468 11152 4480
rect 9999 4440 11152 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 13633 4471 13691 4477
rect 13633 4437 13645 4471
rect 13679 4468 13691 4471
rect 14090 4468 14096 4480
rect 13679 4440 14096 4468
rect 13679 4437 13691 4440
rect 13633 4431 13691 4437
rect 14090 4428 14096 4440
rect 14148 4428 14154 4480
rect 16945 4471 17003 4477
rect 16945 4437 16957 4471
rect 16991 4468 17003 4471
rect 18138 4468 18144 4480
rect 16991 4440 18144 4468
rect 16991 4437 17003 4440
rect 16945 4431 17003 4437
rect 18138 4428 18144 4440
rect 18196 4428 18202 4480
rect 19702 4428 19708 4480
rect 19760 4468 19766 4480
rect 19889 4471 19947 4477
rect 19889 4468 19901 4471
rect 19760 4440 19901 4468
rect 19760 4428 19766 4440
rect 19889 4437 19901 4440
rect 19935 4437 19947 4471
rect 19889 4431 19947 4437
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 3142 4264 3148 4276
rect 2792 4236 3148 4264
rect 2792 4137 2820 4236
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 4154 4264 4160 4276
rect 4115 4236 4160 4264
rect 4154 4224 4160 4236
rect 4212 4224 4218 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6420 4236 15056 4264
rect 6420 4224 6426 4236
rect 7009 4199 7067 4205
rect 7009 4165 7021 4199
rect 7055 4196 7067 4199
rect 10594 4196 10600 4208
rect 7055 4168 7788 4196
rect 7055 4165 7067 4168
rect 7009 4159 7067 4165
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4097 2835 4131
rect 2777 4091 2835 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4097 5779 4131
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 5721 4091 5779 4097
rect 3044 4063 3102 4069
rect 3044 4029 3056 4063
rect 3090 4060 3102 4063
rect 5736 4060 5764 4091
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7760 4128 7788 4168
rect 9600 4168 10600 4196
rect 8478 4128 8484 4140
rect 7760 4100 8484 4128
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 5810 4060 5816 4072
rect 3090 4032 5816 4060
rect 3090 4029 3102 4032
rect 3044 4023 3102 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 8573 4063 8631 4069
rect 7524 4032 7569 4060
rect 7524 4020 7530 4032
rect 8573 4029 8585 4063
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 8840 4063 8898 4069
rect 8840 4029 8852 4063
rect 8886 4060 8898 4063
rect 9600 4060 9628 4168
rect 10594 4156 10600 4168
rect 10652 4156 10658 4208
rect 13817 4199 13875 4205
rect 13817 4165 13829 4199
rect 13863 4196 13875 4199
rect 14274 4196 14280 4208
rect 13863 4168 14280 4196
rect 13863 4165 13875 4168
rect 13817 4159 13875 4165
rect 14274 4156 14280 4168
rect 14332 4196 14338 4208
rect 14734 4196 14740 4208
rect 14332 4168 14740 4196
rect 14332 4156 14338 4168
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 13964 4100 14504 4128
rect 13964 4088 13970 4100
rect 8886 4032 9628 4060
rect 8886 4029 8898 4032
rect 8840 4023 8898 4029
rect 842 3952 848 4004
rect 900 3992 906 4004
rect 3234 3992 3240 4004
rect 900 3964 3240 3992
rect 900 3952 906 3964
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 5537 3995 5595 4001
rect 5537 3992 5549 3995
rect 3344 3964 5549 3992
rect 1765 3927 1823 3933
rect 1765 3893 1777 3927
rect 1811 3924 1823 3927
rect 3344 3924 3372 3964
rect 5537 3961 5549 3964
rect 5583 3961 5595 3995
rect 5537 3955 5595 3961
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 8588 3992 8616 4023
rect 9674 4020 9680 4072
rect 9732 4060 9738 4072
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 9732 4032 10793 4060
rect 9732 4020 9738 4032
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10870 4020 10876 4072
rect 10928 4060 10934 4072
rect 11974 4060 11980 4072
rect 10928 4032 11980 4060
rect 10928 4020 10934 4032
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 12437 4063 12495 4069
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12437 4023 12495 4029
rect 9490 3992 9496 4004
rect 5776 3964 6776 3992
rect 8588 3964 9496 3992
rect 5776 3952 5782 3964
rect 5166 3924 5172 3936
rect 1811 3896 3372 3924
rect 5127 3896 5172 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5408 3896 5641 3924
rect 5408 3884 5414 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 6638 3924 6644 3936
rect 5960 3896 6644 3924
rect 5960 3884 5966 3896
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 6748 3924 6776 3964
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 10594 3992 10600 4004
rect 9784 3964 10600 3992
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 6748 3896 7389 3924
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 9784 3924 9812 3964
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10686 3952 10692 4004
rect 10744 3992 10750 4004
rect 11057 3995 11115 4001
rect 11057 3992 11069 3995
rect 10744 3964 11069 3992
rect 10744 3952 10750 3964
rect 11057 3961 11069 3964
rect 11103 3961 11115 3995
rect 12452 3992 12480 4023
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12693 4063 12751 4069
rect 12693 4060 12705 4063
rect 12584 4032 12705 4060
rect 12584 4020 12590 4032
rect 12693 4029 12705 4032
rect 12739 4029 12751 4063
rect 14274 4060 14280 4072
rect 12693 4023 12751 4029
rect 12820 4032 14280 4060
rect 12820 3992 12848 4032
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 12452 3964 12848 3992
rect 14476 3992 14504 4100
rect 15028 4069 15056 4236
rect 17052 4168 19472 4196
rect 17052 4137 17080 4168
rect 15197 4131 15255 4137
rect 15197 4097 15209 4131
rect 15243 4097 15255 4131
rect 15197 4091 15255 4097
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4097 17095 4131
rect 19444 4128 19472 4168
rect 17037 4091 17095 4097
rect 17144 4100 18828 4128
rect 19444 4100 19564 4128
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 15105 3995 15163 4001
rect 15105 3992 15117 3995
rect 14476 3964 15117 3992
rect 11057 3955 11115 3961
rect 15105 3961 15117 3964
rect 15151 3961 15163 3995
rect 15105 3955 15163 3961
rect 9950 3924 9956 3936
rect 7800 3896 9812 3924
rect 9911 3896 9956 3924
rect 7800 3884 7806 3896
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 11238 3924 11244 3936
rect 10284 3896 11244 3924
rect 10284 3884 10290 3896
rect 11238 3884 11244 3896
rect 11296 3884 11302 3936
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14056 3896 14657 3924
rect 14056 3884 14062 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 14645 3887 14703 3893
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 15212 3924 15240 4091
rect 15746 4020 15752 4072
rect 15804 4060 15810 4072
rect 16758 4060 16764 4072
rect 15804 4032 16764 4060
rect 15804 4020 15810 4032
rect 16758 4020 16764 4032
rect 16816 4060 16822 4072
rect 17144 4060 17172 4100
rect 16816 4032 17172 4060
rect 16816 4020 16822 4032
rect 17494 4020 17500 4072
rect 17552 4060 17558 4072
rect 18325 4063 18383 4069
rect 18325 4060 18337 4063
rect 17552 4032 18337 4060
rect 17552 4020 17558 4032
rect 18325 4029 18337 4032
rect 18371 4029 18383 4063
rect 18800 4060 18828 4100
rect 19429 4063 19487 4069
rect 19429 4060 19441 4063
rect 18800 4032 19441 4060
rect 18325 4023 18383 4029
rect 19429 4029 19441 4032
rect 19475 4029 19487 4063
rect 19536 4060 19564 4100
rect 19702 4069 19708 4072
rect 19685 4063 19708 4069
rect 19685 4060 19697 4063
rect 19536 4032 19697 4060
rect 19429 4023 19487 4029
rect 19685 4029 19697 4032
rect 19760 4060 19766 4072
rect 19760 4032 19833 4060
rect 19685 4023 19708 4029
rect 19702 4020 19708 4023
rect 19760 4020 19766 4032
rect 22646 3992 22652 4004
rect 18524 3964 22652 3992
rect 14792 3896 15240 3924
rect 16393 3927 16451 3933
rect 14792 3884 14798 3896
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 16574 3924 16580 3936
rect 16439 3896 16580 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16758 3924 16764 3936
rect 16719 3896 16764 3924
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 18046 3924 18052 3936
rect 16899 3896 18052 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18524 3933 18552 3964
rect 22646 3952 22652 3964
rect 22704 3952 22710 4004
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3893 18567 3927
rect 18509 3887 18567 3893
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 20809 3927 20867 3933
rect 20809 3924 20821 3927
rect 19944 3896 20821 3924
rect 19944 3884 19950 3896
rect 20809 3893 20821 3896
rect 20855 3893 20867 3927
rect 20809 3887 20867 3893
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1780 3692 3188 3720
rect 1780 3593 1808 3692
rect 3160 3652 3188 3692
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 5534 3720 5540 3732
rect 3292 3692 5540 3720
rect 3292 3680 3298 3692
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5810 3720 5816 3732
rect 5771 3692 5816 3720
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 5902 3680 5908 3732
rect 5960 3720 5966 3732
rect 9582 3720 9588 3732
rect 5960 3692 9588 3720
rect 5960 3680 5966 3692
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 9824 3692 11069 3720
rect 9824 3680 9830 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 11057 3683 11115 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14090 3680 14096 3732
rect 14148 3720 14154 3732
rect 14148 3692 14193 3720
rect 14148 3680 14154 3692
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 15378 3720 15384 3732
rect 14424 3692 15384 3720
rect 14424 3680 14430 3692
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15528 3692 16160 3720
rect 15528 3680 15534 3692
rect 3160 3624 10732 3652
rect 1765 3587 1823 3593
rect 1765 3553 1777 3587
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 2682 3544 2688 3596
rect 2740 3584 2746 3596
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 2740 3556 2881 3584
rect 2740 3544 2746 3556
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 4700 3587 4758 3593
rect 4700 3553 4712 3587
rect 4746 3584 4758 3587
rect 5442 3584 5448 3596
rect 4746 3556 5448 3584
rect 4746 3553 4758 3556
rect 4700 3547 4758 3553
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 7000 3587 7058 3593
rect 7000 3553 7012 3587
rect 7046 3584 7058 3587
rect 9766 3584 9772 3596
rect 7046 3556 9772 3584
rect 7046 3553 7058 3556
rect 7000 3547 7058 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9950 3593 9956 3596
rect 9944 3584 9956 3593
rect 9863 3556 9956 3584
rect 9944 3547 9956 3556
rect 10008 3584 10014 3596
rect 10318 3584 10324 3596
rect 10008 3556 10324 3584
rect 9950 3544 9956 3547
rect 10008 3544 10014 3556
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 290 3476 296 3528
rect 348 3516 354 3528
rect 348 3488 4384 3516
rect 348 3476 354 3488
rect 1394 3408 1400 3460
rect 1452 3448 1458 3460
rect 4246 3448 4252 3460
rect 1452 3420 4252 3448
rect 1452 3408 1458 3420
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2866 3380 2872 3392
rect 1995 3352 2872 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 3050 3380 3056 3392
rect 3011 3352 3056 3380
rect 3050 3340 3056 3352
rect 3108 3340 3114 3392
rect 4356 3380 4384 3488
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 4488 3488 4533 3516
rect 4488 3476 4494 3488
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 6840 3516 6868 3544
rect 5868 3488 6868 3516
rect 5868 3476 5874 3488
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 9306 3516 9312 3528
rect 8352 3488 9312 3516
rect 8352 3476 8358 3488
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9548 3488 9689 3516
rect 9548 3476 9554 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 10704 3516 10732 3624
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 16132 3652 16160 3692
rect 16758 3680 16764 3732
rect 16816 3720 16822 3732
rect 17957 3723 18015 3729
rect 17957 3720 17969 3723
rect 16816 3692 17969 3720
rect 16816 3680 16822 3692
rect 17957 3689 17969 3692
rect 18003 3689 18015 3723
rect 17957 3683 18015 3689
rect 18417 3723 18475 3729
rect 18417 3689 18429 3723
rect 18463 3720 18475 3723
rect 19242 3720 19248 3732
rect 18463 3692 19248 3720
rect 18463 3689 18475 3692
rect 18417 3683 18475 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 17773 3655 17831 3661
rect 17773 3652 17785 3655
rect 11204 3624 14044 3652
rect 16132 3624 17785 3652
rect 11204 3612 11210 3624
rect 14016 3596 14044 3624
rect 17773 3621 17785 3624
rect 17819 3652 17831 3655
rect 18325 3655 18383 3661
rect 18325 3652 18337 3655
rect 17819 3624 18337 3652
rect 17819 3621 17831 3624
rect 17773 3615 17831 3621
rect 18325 3621 18337 3624
rect 18371 3621 18383 3655
rect 18325 3615 18383 3621
rect 11882 3584 11888 3596
rect 11843 3556 11888 3584
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 13906 3584 13912 3596
rect 12176 3556 13912 3584
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 10704 3488 12081 3516
rect 9677 3479 9735 3485
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 12069 3479 12127 3485
rect 7668 3420 8248 3448
rect 7668 3380 7696 3420
rect 4356 3352 7696 3380
rect 7742 3340 7748 3392
rect 7800 3380 7806 3392
rect 8113 3383 8171 3389
rect 8113 3380 8125 3383
rect 7800 3352 8125 3380
rect 7800 3340 7806 3352
rect 8113 3349 8125 3352
rect 8159 3349 8171 3383
rect 8220 3380 8248 3420
rect 12176 3380 12204 3556
rect 13906 3544 13912 3556
rect 13964 3544 13970 3596
rect 13998 3544 14004 3596
rect 14056 3544 14062 3596
rect 15654 3584 15660 3596
rect 14292 3556 15660 3584
rect 14292 3525 14320 3556
rect 15654 3544 15660 3556
rect 15712 3584 15718 3596
rect 16005 3587 16063 3593
rect 16005 3584 16017 3587
rect 15712 3556 16017 3584
rect 15712 3544 15718 3556
rect 16005 3553 16017 3556
rect 16051 3553 16063 3587
rect 16005 3547 16063 3553
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 18690 3584 18696 3596
rect 16448 3556 18696 3584
rect 16448 3544 16454 3556
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 18782 3544 18788 3596
rect 18840 3584 18846 3596
rect 19521 3587 19579 3593
rect 19521 3584 19533 3587
rect 18840 3556 19533 3584
rect 18840 3544 18846 3556
rect 19521 3553 19533 3556
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 20254 3544 20260 3596
rect 20312 3584 20318 3596
rect 22094 3584 22100 3596
rect 20312 3556 22100 3584
rect 20312 3544 20318 3556
rect 22094 3544 22100 3556
rect 22152 3544 22158 3596
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14458 3476 14464 3528
rect 14516 3516 14522 3528
rect 15470 3516 15476 3528
rect 14516 3488 15476 3516
rect 14516 3476 14522 3488
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15746 3516 15752 3528
rect 15707 3488 15752 3516
rect 15746 3476 15752 3488
rect 15804 3476 15810 3528
rect 17770 3516 17776 3528
rect 17144 3488 17776 3516
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 15764 3448 15792 3476
rect 17144 3457 17172 3488
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3485 19763 3519
rect 19705 3479 19763 3485
rect 14884 3420 15792 3448
rect 17129 3451 17187 3457
rect 14884 3408 14890 3420
rect 17129 3417 17141 3451
rect 17175 3417 17187 3451
rect 17129 3411 17187 3417
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 19720 3448 19748 3479
rect 17920 3420 19748 3448
rect 17920 3408 17926 3420
rect 8220 3352 12204 3380
rect 13633 3383 13691 3389
rect 8113 3343 8171 3349
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13906 3380 13912 3392
rect 13679 3352 13912 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 17034 3380 17040 3392
rect 14056 3352 17040 3380
rect 14056 3340 14062 3352
rect 17034 3340 17040 3352
rect 17092 3340 17098 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 5442 3176 5448 3188
rect 2792 3148 5304 3176
rect 5403 3148 5448 3176
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2792 2972 2820 3148
rect 3145 3111 3203 3117
rect 3145 3077 3157 3111
rect 3191 3077 3203 3111
rect 5276 3108 5304 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 6840 3148 7972 3176
rect 6840 3108 6868 3148
rect 5276 3080 6868 3108
rect 3145 3071 3203 3077
rect 3160 3040 3188 3071
rect 3160 3012 4200 3040
rect 2958 2972 2964 2984
rect 1903 2944 2820 2972
rect 2919 2944 2964 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 4062 2972 4068 2984
rect 3200 2944 4068 2972
rect 3200 2932 3206 2944
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4172 2972 4200 3012
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6788 3012 6837 3040
rect 6788 3000 6794 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 5902 2972 5908 2984
rect 4172 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 4332 2907 4390 2913
rect 4332 2873 4344 2907
rect 4378 2904 4390 2907
rect 6914 2904 6920 2916
rect 4378 2876 6920 2904
rect 4378 2873 4390 2876
rect 4332 2867 4390 2873
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 7092 2907 7150 2913
rect 7092 2873 7104 2907
rect 7138 2904 7150 2907
rect 7374 2904 7380 2916
rect 7138 2876 7380 2904
rect 7138 2873 7150 2876
rect 7092 2867 7150 2873
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 7944 2904 7972 3148
rect 8110 3136 8116 3188
rect 8168 3176 8174 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 8168 3148 8217 3176
rect 8168 3136 8174 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 8205 3139 8263 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 10870 3176 10876 3188
rect 10284 3148 10876 3176
rect 10284 3136 10290 3148
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11425 3179 11483 3185
rect 11425 3145 11437 3179
rect 11471 3176 11483 3179
rect 11471 3148 15608 3176
rect 11471 3145 11483 3148
rect 11425 3139 11483 3145
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 12526 3108 12532 3120
rect 8352 3080 12532 3108
rect 8352 3068 8358 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 15580 3108 15608 3148
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15712 3148 15761 3176
rect 15712 3136 15718 3148
rect 15749 3145 15761 3148
rect 15795 3145 15807 3179
rect 18046 3176 18052 3188
rect 18007 3148 18052 3176
rect 15749 3139 15807 3145
rect 18046 3136 18052 3148
rect 18104 3136 18110 3188
rect 19334 3108 19340 3120
rect 15580 3080 19340 3108
rect 19334 3068 19340 3080
rect 19392 3068 19398 3120
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 9824 3012 10241 3040
rect 9824 3000 9830 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 14274 3040 14280 3052
rect 10229 3003 10287 3009
rect 10336 3012 14280 3040
rect 8202 2932 8208 2984
rect 8260 2972 8266 2984
rect 10336 2972 10364 3012
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14366 3000 14372 3052
rect 14424 3040 14430 3052
rect 16850 3040 16856 3052
rect 14424 3012 14469 3040
rect 16811 3012 16856 3040
rect 14424 3000 14430 3012
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 19116 3012 20177 3040
rect 19116 3000 19122 3012
rect 20165 3009 20177 3012
rect 20211 3009 20223 3043
rect 20165 3003 20223 3009
rect 8260 2944 10364 2972
rect 11241 2975 11299 2981
rect 8260 2932 8266 2944
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 12342 2972 12348 2984
rect 11287 2944 12348 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12713 2975 12771 2981
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 15562 2972 15568 2984
rect 12759 2944 13216 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 12989 2907 13047 2913
rect 12989 2904 13001 2907
rect 7944 2876 13001 2904
rect 12989 2873 13001 2876
rect 13035 2873 13047 2907
rect 13188 2904 13216 2944
rect 14476 2944 15568 2972
rect 14476 2904 14504 2944
rect 15562 2932 15568 2944
rect 15620 2932 15626 2984
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16632 2944 16681 2972
rect 16632 2932 16638 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 18138 2932 18144 2984
rect 18196 2972 18202 2984
rect 18509 2975 18567 2981
rect 18509 2972 18521 2975
rect 18196 2944 18521 2972
rect 18196 2932 18202 2944
rect 18509 2941 18521 2944
rect 18555 2941 18567 2975
rect 18509 2935 18567 2941
rect 19981 2975 20039 2981
rect 19981 2941 19993 2975
rect 20027 2972 20039 2975
rect 20070 2972 20076 2984
rect 20027 2944 20076 2972
rect 20027 2941 20039 2944
rect 19981 2935 20039 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 13188 2876 14504 2904
rect 14636 2907 14694 2913
rect 12989 2867 13047 2873
rect 14636 2873 14648 2907
rect 14682 2904 14694 2907
rect 14734 2904 14740 2916
rect 14682 2876 14740 2904
rect 14682 2873 14694 2876
rect 14636 2867 14694 2873
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 18417 2907 18475 2913
rect 18417 2904 18429 2907
rect 18012 2876 18429 2904
rect 18012 2864 18018 2876
rect 18417 2873 18429 2876
rect 18463 2873 18475 2907
rect 18417 2867 18475 2873
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10137 2839 10195 2845
rect 10137 2805 10149 2839
rect 10183 2836 10195 2839
rect 10502 2836 10508 2848
rect 10183 2808 10508 2836
rect 10183 2805 10195 2808
rect 10137 2799 10195 2805
rect 10502 2796 10508 2808
rect 10560 2796 10566 2848
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 13722 2836 13728 2848
rect 10652 2808 13728 2836
rect 10652 2796 10658 2808
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 14550 2796 14556 2848
rect 14608 2836 14614 2848
rect 18138 2836 18144 2848
rect 14608 2808 18144 2836
rect 14608 2796 14614 2808
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 19610 2836 19616 2848
rect 19571 2808 19616 2836
rect 19610 2796 19616 2808
rect 19668 2796 19674 2848
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 20073 2839 20131 2845
rect 20073 2836 20085 2839
rect 19852 2808 20085 2836
rect 19852 2796 19858 2808
rect 20073 2805 20085 2808
rect 20119 2805 20131 2839
rect 20073 2799 20131 2805
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5350 2632 5356 2644
rect 4939 2604 5356 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 7193 2635 7251 2641
rect 7193 2601 7205 2635
rect 7239 2632 7251 2635
rect 7466 2632 7472 2644
rect 7239 2604 7472 2632
rect 7239 2601 7251 2604
rect 7193 2595 7251 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7653 2635 7711 2641
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 9674 2632 9680 2644
rect 7699 2604 9680 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 10502 2632 10508 2644
rect 9815 2604 10508 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 11609 2635 11667 2641
rect 11609 2601 11621 2635
rect 11655 2632 11667 2635
rect 18782 2632 18788 2644
rect 11655 2604 18788 2632
rect 11655 2601 11667 2604
rect 11609 2595 11667 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 2884 2536 10548 2564
rect 2884 2505 2912 2536
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 5261 2499 5319 2505
rect 5261 2496 5273 2499
rect 4856 2468 5273 2496
rect 4856 2456 4862 2468
rect 5261 2465 5273 2468
rect 5307 2465 5319 2499
rect 5261 2459 5319 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7561 2499 7619 2505
rect 7561 2496 7573 2499
rect 7064 2468 7573 2496
rect 7064 2456 7070 2468
rect 7561 2465 7573 2468
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 9214 2456 9220 2508
rect 9272 2496 9278 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9272 2468 10149 2496
rect 9272 2456 9278 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10229 2499 10287 2505
rect 10229 2465 10241 2499
rect 10275 2496 10287 2499
rect 10410 2496 10416 2508
rect 10275 2468 10416 2496
rect 10275 2465 10287 2468
rect 10229 2459 10287 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 1872 2360 1900 2391
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5132 2400 5365 2428
rect 5132 2388 5138 2400
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 7742 2428 7748 2440
rect 5500 2400 5545 2428
rect 7703 2400 7748 2428
rect 5500 2388 5506 2400
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10520 2428 10548 2536
rect 11440 2536 13768 2564
rect 11440 2505 11468 2536
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2465 11483 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 11425 2459 11483 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 10376 2400 10421 2428
rect 10520 2400 12817 2428
rect 10376 2388 10382 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 13740 2428 13768 2536
rect 13814 2524 13820 2576
rect 13872 2564 13878 2576
rect 14185 2567 14243 2573
rect 14185 2564 14197 2567
rect 13872 2536 14197 2564
rect 13872 2524 13878 2536
rect 14185 2533 14197 2536
rect 14231 2533 14243 2567
rect 17862 2564 17868 2576
rect 14185 2527 14243 2533
rect 16040 2536 17868 2564
rect 13906 2496 13912 2508
rect 13867 2468 13912 2496
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 16040 2505 16068 2536
rect 17862 2524 17868 2536
rect 17920 2524 17926 2576
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2465 16083 2499
rect 17126 2496 17132 2508
rect 17087 2468 17132 2496
rect 16025 2459 16083 2465
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 18969 2499 19027 2505
rect 18969 2465 18981 2499
rect 19015 2496 19027 2499
rect 19610 2496 19616 2508
rect 19015 2468 19616 2496
rect 19015 2465 19027 2468
rect 18969 2459 19027 2465
rect 19610 2456 19616 2468
rect 19668 2456 19674 2508
rect 19153 2431 19211 2437
rect 19153 2428 19165 2431
rect 13740 2400 19165 2428
rect 12805 2391 12863 2397
rect 19153 2397 19165 2400
rect 19199 2397 19211 2431
rect 19153 2391 19211 2397
rect 5718 2360 5724 2372
rect 1872 2332 5724 2360
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 7190 2320 7196 2372
rect 7248 2360 7254 2372
rect 8110 2360 8116 2372
rect 7248 2332 8116 2360
rect 7248 2320 7254 2332
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 9766 2320 9772 2372
rect 9824 2360 9830 2372
rect 10134 2360 10140 2372
rect 9824 2332 10140 2360
rect 9824 2320 9830 2332
rect 10134 2320 10140 2332
rect 10192 2320 10198 2372
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 11790 2360 11796 2372
rect 10928 2332 11796 2360
rect 10928 2320 10934 2332
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 16209 2363 16267 2369
rect 16209 2329 16221 2363
rect 16255 2360 16267 2363
rect 20990 2360 20996 2372
rect 16255 2332 20996 2360
rect 16255 2329 16267 2332
rect 16209 2323 16267 2329
rect 20990 2320 20996 2332
rect 21048 2320 21054 2372
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 17313 2295 17371 2301
rect 17313 2261 17325 2295
rect 17359 2292 17371 2295
rect 17678 2292 17684 2304
rect 17359 2264 17684 2292
rect 17359 2261 17371 2264
rect 17313 2255 17371 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3050 2048 3056 2100
rect 3108 2088 3114 2100
rect 13170 2088 13176 2100
rect 3108 2060 13176 2088
rect 3108 2048 3114 2060
rect 13170 2048 13176 2060
rect 13228 2048 13234 2100
rect 5074 1980 5080 2032
rect 5132 2020 5138 2032
rect 17954 2020 17960 2032
rect 5132 1992 17960 2020
rect 5132 1980 5138 1992
rect 17954 1980 17960 1992
rect 18012 1980 18018 2032
rect 10778 1912 10784 1964
rect 10836 1952 10842 1964
rect 15930 1952 15936 1964
rect 10836 1924 15936 1952
rect 10836 1912 10842 1924
rect 15930 1912 15936 1924
rect 15988 1912 15994 1964
rect 9398 1300 9404 1352
rect 9456 1340 9462 1352
rect 18138 1340 18144 1352
rect 9456 1312 18144 1340
rect 9456 1300 9462 1312
rect 18138 1300 18144 1312
rect 18196 1300 18202 1352
rect 10410 1232 10416 1284
rect 10468 1272 10474 1284
rect 18046 1272 18052 1284
rect 10468 1244 18052 1272
rect 10468 1232 10474 1244
rect 18046 1232 18052 1244
rect 18104 1232 18110 1284
rect 9674 1164 9680 1216
rect 9732 1204 9738 1216
rect 10962 1204 10968 1216
rect 9732 1176 10968 1204
rect 9732 1164 9738 1176
rect 10962 1164 10968 1176
rect 11020 1204 11026 1216
rect 17954 1204 17960 1216
rect 11020 1176 17960 1204
rect 11020 1164 11026 1176
rect 17954 1164 17960 1176
rect 18012 1164 18018 1216
<< via1 >>
rect 10232 21088 10284 21140
rect 18328 21088 18380 21140
rect 3148 20952 3200 21004
rect 18696 20952 18748 21004
rect 2872 20884 2924 20936
rect 17960 20884 18012 20936
rect 2228 20816 2280 20868
rect 18052 20816 18104 20868
rect 1952 20748 2004 20800
rect 18144 20748 18196 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 1952 20587 2004 20596
rect 1952 20553 1961 20587
rect 1961 20553 1995 20587
rect 1995 20553 2004 20587
rect 1952 20544 2004 20553
rect 3148 20544 3200 20596
rect 3240 20544 3292 20596
rect 18144 20544 18196 20596
rect 5448 20476 5500 20528
rect 6920 20519 6972 20528
rect 6920 20485 6929 20519
rect 6929 20485 6963 20519
rect 6963 20485 6972 20519
rect 6920 20476 6972 20485
rect 7564 20476 7616 20528
rect 11060 20476 11112 20528
rect 11152 20476 11204 20528
rect 3148 20340 3200 20392
rect 4804 20408 4856 20460
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 6828 20408 6880 20460
rect 8484 20408 8536 20460
rect 5724 20340 5776 20392
rect 6184 20340 6236 20392
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 10324 20340 10376 20392
rect 20352 20476 20404 20528
rect 14188 20408 14240 20460
rect 14740 20408 14792 20460
rect 19616 20408 19668 20460
rect 6736 20272 6788 20324
rect 2504 20204 2556 20256
rect 2872 20204 2924 20256
rect 5080 20204 5132 20256
rect 5264 20204 5316 20256
rect 6368 20204 6420 20256
rect 9864 20272 9916 20324
rect 10140 20272 10192 20324
rect 10600 20204 10652 20256
rect 11796 20272 11848 20324
rect 14004 20272 14056 20324
rect 14372 20272 14424 20324
rect 12256 20204 12308 20256
rect 13268 20204 13320 20256
rect 13820 20204 13872 20256
rect 17224 20340 17276 20392
rect 19708 20383 19760 20392
rect 19708 20349 19717 20383
rect 19717 20349 19751 20383
rect 19751 20349 19760 20383
rect 19708 20340 19760 20349
rect 15568 20272 15620 20324
rect 15660 20204 15712 20256
rect 16212 20204 16264 20256
rect 17776 20204 17828 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2228 20000 2280 20052
rect 4804 19932 4856 19984
rect 5172 19932 5224 19984
rect 9680 20000 9732 20052
rect 11704 20000 11756 20052
rect 13268 20000 13320 20052
rect 17868 20000 17920 20052
rect 9772 19932 9824 19984
rect 9956 19975 10008 19984
rect 9956 19941 9990 19975
rect 9990 19941 10008 19975
rect 9956 19932 10008 19941
rect 6644 19864 6696 19916
rect 6828 19864 6880 19916
rect 7472 19864 7524 19916
rect 13360 19864 13412 19916
rect 4252 19839 4304 19848
rect 4252 19805 4261 19839
rect 4261 19805 4295 19839
rect 4295 19805 4304 19839
rect 4252 19796 4304 19805
rect 5632 19703 5684 19712
rect 5632 19669 5641 19703
rect 5641 19669 5675 19703
rect 5675 19669 5684 19703
rect 9680 19839 9732 19848
rect 9680 19805 9696 19839
rect 9696 19805 9730 19839
rect 9730 19805 9732 19839
rect 9680 19796 9732 19805
rect 11060 19796 11112 19848
rect 11888 19796 11940 19848
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 13636 19796 13688 19848
rect 16028 19864 16080 19916
rect 18052 19864 18104 19916
rect 19524 19907 19576 19916
rect 19524 19873 19533 19907
rect 19533 19873 19567 19907
rect 19567 19873 19576 19907
rect 19524 19864 19576 19873
rect 8024 19728 8076 19780
rect 16120 19796 16172 19848
rect 17132 19796 17184 19848
rect 5632 19660 5684 19669
rect 8116 19660 8168 19712
rect 8392 19660 8444 19712
rect 15844 19728 15896 19780
rect 17316 19728 17368 19780
rect 10968 19660 11020 19712
rect 14188 19660 14240 19712
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1400 19456 1452 19508
rect 4804 19431 4856 19440
rect 4804 19397 4813 19431
rect 4813 19397 4847 19431
rect 4847 19397 4856 19431
rect 4804 19388 4856 19397
rect 7564 19388 7616 19440
rect 8024 19388 8076 19440
rect 9956 19456 10008 19508
rect 10140 19456 10192 19508
rect 10600 19456 10652 19508
rect 13084 19456 13136 19508
rect 17132 19456 17184 19508
rect 19524 19456 19576 19508
rect 3332 19320 3384 19372
rect 2412 19252 2464 19304
rect 2596 19252 2648 19304
rect 7472 19320 7524 19372
rect 848 19184 900 19236
rect 2872 19184 2924 19236
rect 2504 19159 2556 19168
rect 2504 19125 2513 19159
rect 2513 19125 2547 19159
rect 2547 19125 2556 19159
rect 2504 19116 2556 19125
rect 5908 19252 5960 19304
rect 6092 19252 6144 19304
rect 8116 19295 8168 19304
rect 8116 19261 8125 19295
rect 8125 19261 8159 19295
rect 8159 19261 8168 19295
rect 8116 19252 8168 19261
rect 8392 19295 8444 19304
rect 8392 19261 8426 19295
rect 8426 19261 8444 19295
rect 8392 19252 8444 19261
rect 8668 19252 8720 19304
rect 4160 19184 4212 19236
rect 6644 19184 6696 19236
rect 8300 19184 8352 19236
rect 9680 19320 9732 19372
rect 10416 19320 10468 19372
rect 10968 19363 11020 19372
rect 9220 19252 9272 19304
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 20168 19363 20220 19372
rect 20168 19329 20177 19363
rect 20177 19329 20211 19363
rect 20211 19329 20220 19363
rect 20168 19320 20220 19329
rect 12624 19252 12676 19304
rect 12900 19252 12952 19304
rect 13268 19252 13320 19304
rect 15108 19252 15160 19304
rect 16120 19252 16172 19304
rect 16948 19252 17000 19304
rect 13452 19227 13504 19236
rect 13452 19193 13486 19227
rect 13486 19193 13504 19227
rect 13452 19184 13504 19193
rect 4344 19116 4396 19168
rect 5540 19116 5592 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 6460 19116 6512 19168
rect 9312 19116 9364 19168
rect 9496 19159 9548 19168
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 10324 19159 10376 19168
rect 10324 19125 10333 19159
rect 10333 19125 10367 19159
rect 10367 19125 10376 19159
rect 10324 19116 10376 19125
rect 10876 19116 10928 19168
rect 14372 19116 14424 19168
rect 15844 19184 15896 19236
rect 17132 19184 17184 19236
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 16764 19159 16816 19168
rect 16764 19125 16773 19159
rect 16773 19125 16807 19159
rect 16807 19125 16816 19159
rect 16764 19116 16816 19125
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 3240 18912 3292 18964
rect 5816 18912 5868 18964
rect 13268 18912 13320 18964
rect 13452 18912 13504 18964
rect 15476 18912 15528 18964
rect 17224 18912 17276 18964
rect 2596 18776 2648 18828
rect 4068 18776 4120 18828
rect 5172 18844 5224 18896
rect 5632 18844 5684 18896
rect 6000 18844 6052 18896
rect 6644 18844 6696 18896
rect 7012 18844 7064 18896
rect 5540 18776 5592 18828
rect 10416 18844 10468 18896
rect 10968 18844 11020 18896
rect 11060 18844 11112 18896
rect 11980 18844 12032 18896
rect 12072 18844 12124 18896
rect 16764 18844 16816 18896
rect 5356 18708 5408 18760
rect 6644 18708 6696 18760
rect 7012 18708 7064 18760
rect 8668 18776 8720 18828
rect 8944 18776 8996 18828
rect 12348 18776 12400 18828
rect 12624 18776 12676 18828
rect 13084 18776 13136 18828
rect 17960 18776 18012 18828
rect 5264 18640 5316 18692
rect 6828 18683 6880 18692
rect 6828 18649 6837 18683
rect 6837 18649 6871 18683
rect 6871 18649 6880 18683
rect 6828 18640 6880 18649
rect 1492 18572 1544 18624
rect 2964 18572 3016 18624
rect 3792 18572 3844 18624
rect 7196 18640 7248 18692
rect 9680 18708 9732 18760
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 16120 18708 16172 18760
rect 20996 18844 21048 18896
rect 18144 18776 18196 18828
rect 18972 18751 19024 18760
rect 8760 18640 8812 18692
rect 11336 18640 11388 18692
rect 13544 18640 13596 18692
rect 9128 18572 9180 18624
rect 9312 18572 9364 18624
rect 13176 18572 13228 18624
rect 13268 18572 13320 18624
rect 14648 18572 14700 18624
rect 18972 18717 18981 18751
rect 18981 18717 19015 18751
rect 19015 18717 19024 18751
rect 18972 18708 19024 18717
rect 19156 18751 19208 18760
rect 19156 18717 19165 18751
rect 19165 18717 19199 18751
rect 19199 18717 19208 18751
rect 19156 18708 19208 18717
rect 17592 18572 17644 18624
rect 18144 18572 18196 18624
rect 18788 18572 18840 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 5172 18368 5224 18420
rect 6644 18368 6696 18420
rect 6736 18368 6788 18420
rect 8208 18368 8260 18420
rect 10692 18368 10744 18420
rect 16028 18368 16080 18420
rect 5356 18300 5408 18352
rect 5816 18232 5868 18284
rect 6736 18232 6788 18284
rect 9128 18275 9180 18284
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 2504 18207 2556 18216
rect 2504 18173 2513 18207
rect 2513 18173 2547 18207
rect 2547 18173 2556 18207
rect 2504 18164 2556 18173
rect 2596 18164 2648 18216
rect 5540 18207 5592 18216
rect 3516 18096 3568 18148
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 6000 18164 6052 18216
rect 7288 18164 7340 18216
rect 8484 18096 8536 18148
rect 8852 18164 8904 18216
rect 9496 18232 9548 18284
rect 9588 18232 9640 18284
rect 11060 18232 11112 18284
rect 11888 18232 11940 18284
rect 14004 18232 14056 18284
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 16764 18232 16816 18284
rect 20352 18232 20404 18284
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 11796 18164 11848 18216
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 12440 18164 12492 18173
rect 10876 18096 10928 18148
rect 13084 18164 13136 18216
rect 15292 18164 15344 18216
rect 15844 18164 15896 18216
rect 17500 18164 17552 18216
rect 19156 18164 19208 18216
rect 20260 18207 20312 18216
rect 20260 18173 20269 18207
rect 20269 18173 20303 18207
rect 20303 18173 20312 18207
rect 20260 18164 20312 18173
rect 13544 18096 13596 18148
rect 14096 18139 14148 18148
rect 14096 18105 14105 18139
rect 14105 18105 14139 18139
rect 14139 18105 14148 18139
rect 14096 18096 14148 18105
rect 3792 18028 3844 18080
rect 4160 18028 4212 18080
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 5356 18028 5408 18080
rect 7012 18028 7064 18080
rect 7104 18028 7156 18080
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 9128 18028 9180 18080
rect 12164 18028 12216 18080
rect 12532 18028 12584 18080
rect 13728 18028 13780 18080
rect 15476 18096 15528 18148
rect 15568 18096 15620 18148
rect 19524 18096 19576 18148
rect 18144 18028 18196 18080
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 2780 17824 2832 17876
rect 4344 17824 4396 17876
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 6276 17824 6328 17876
rect 2596 17620 2648 17672
rect 3332 17620 3384 17672
rect 5540 17756 5592 17808
rect 5632 17756 5684 17808
rect 6736 17756 6788 17808
rect 7012 17756 7064 17808
rect 12624 17824 12676 17876
rect 18788 17867 18840 17876
rect 15200 17756 15252 17808
rect 18788 17833 18797 17867
rect 18797 17833 18831 17867
rect 18831 17833 18840 17867
rect 18788 17824 18840 17833
rect 19708 17756 19760 17808
rect 6460 17688 6512 17740
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 3516 17552 3568 17604
rect 4804 17552 4856 17604
rect 5448 17620 5500 17672
rect 7472 17688 7524 17740
rect 10140 17688 10192 17740
rect 11244 17731 11296 17740
rect 11244 17697 11278 17731
rect 11278 17697 11296 17731
rect 11244 17688 11296 17697
rect 14188 17688 14240 17740
rect 7380 17620 7432 17672
rect 10968 17663 11020 17672
rect 5264 17552 5316 17604
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 16028 17620 16080 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 18880 17663 18932 17672
rect 16120 17620 16172 17629
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 19432 17688 19484 17740
rect 18604 17552 18656 17604
rect 3700 17484 3752 17536
rect 4896 17484 4948 17536
rect 7656 17484 7708 17536
rect 8208 17484 8260 17536
rect 12808 17484 12860 17536
rect 16488 17484 16540 17536
rect 17224 17484 17276 17536
rect 17684 17484 17736 17536
rect 19800 17484 19852 17536
rect 20444 17484 20496 17536
rect 20812 17484 20864 17536
rect 22100 17484 22152 17536
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 3516 17280 3568 17332
rect 3792 17280 3844 17332
rect 6276 17280 6328 17332
rect 6460 17280 6512 17332
rect 3332 17212 3384 17264
rect 6644 17212 6696 17264
rect 10048 17280 10100 17332
rect 10692 17280 10744 17332
rect 11244 17212 11296 17264
rect 11796 17212 11848 17264
rect 14096 17280 14148 17332
rect 18880 17280 18932 17332
rect 20996 17280 21048 17332
rect 22652 17280 22704 17332
rect 4160 17144 4212 17196
rect 5816 17144 5868 17196
rect 7748 17144 7800 17196
rect 8300 17144 8352 17196
rect 12624 17144 12676 17196
rect 2596 17119 2648 17128
rect 2596 17085 2630 17119
rect 2630 17085 2648 17119
rect 4896 17119 4948 17128
rect 2596 17076 2648 17085
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 2504 17008 2556 17060
rect 2872 17008 2924 17060
rect 7104 17076 7156 17128
rect 8484 17076 8536 17128
rect 12808 17119 12860 17128
rect 1584 16940 1636 16992
rect 5448 17008 5500 17060
rect 8852 17051 8904 17060
rect 8852 17017 8886 17051
rect 8886 17017 8904 17051
rect 8852 17008 8904 17017
rect 12808 17085 12817 17119
rect 12817 17085 12851 17119
rect 12851 17085 12860 17119
rect 12808 17076 12860 17085
rect 14004 17119 14056 17128
rect 14004 17085 14013 17119
rect 14013 17085 14047 17119
rect 14047 17085 14056 17119
rect 14004 17076 14056 17085
rect 17868 17212 17920 17264
rect 14556 17144 14608 17196
rect 18604 17187 18656 17196
rect 14464 17076 14516 17128
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 16488 17076 16540 17128
rect 19340 17212 19392 17264
rect 20444 17212 20496 17264
rect 19156 17144 19208 17196
rect 4160 16940 4212 16992
rect 4896 16940 4948 16992
rect 6276 16940 6328 16992
rect 7012 16940 7064 16992
rect 10416 16940 10468 16992
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 17040 17008 17092 17060
rect 17592 17008 17644 17060
rect 20352 17008 20404 17060
rect 11244 16940 11296 16949
rect 13360 16940 13412 16992
rect 14372 16940 14424 16992
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 18052 16983 18104 16992
rect 15568 16940 15620 16949
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 11244 16779 11296 16788
rect 3792 16668 3844 16720
rect 2504 16600 2556 16652
rect 3700 16600 3752 16652
rect 11244 16745 11253 16779
rect 11253 16745 11287 16779
rect 11287 16745 11296 16779
rect 11244 16736 11296 16745
rect 11704 16779 11756 16788
rect 11704 16745 11713 16779
rect 11713 16745 11747 16779
rect 11747 16745 11756 16779
rect 11704 16736 11756 16745
rect 11888 16736 11940 16788
rect 18052 16736 18104 16788
rect 5172 16668 5224 16720
rect 6828 16668 6880 16720
rect 7012 16668 7064 16720
rect 15568 16668 15620 16720
rect 18604 16668 18656 16720
rect 7288 16600 7340 16652
rect 7840 16600 7892 16652
rect 8208 16600 8260 16652
rect 8392 16600 8444 16652
rect 11152 16600 11204 16652
rect 11244 16600 11296 16652
rect 11704 16600 11756 16652
rect 12900 16600 12952 16652
rect 4804 16575 4856 16584
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 5632 16532 5684 16584
rect 8852 16532 8904 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 15200 16600 15252 16652
rect 14740 16532 14792 16584
rect 4896 16464 4948 16516
rect 18052 16600 18104 16652
rect 16120 16532 16172 16584
rect 16488 16575 16540 16584
rect 16488 16541 16497 16575
rect 16497 16541 16531 16575
rect 16531 16541 16540 16575
rect 16488 16532 16540 16541
rect 20260 16600 20312 16652
rect 19156 16575 19208 16584
rect 19156 16541 19165 16575
rect 19165 16541 19199 16575
rect 19199 16541 19208 16575
rect 19156 16532 19208 16541
rect 1768 16396 1820 16448
rect 7748 16396 7800 16448
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 9864 16396 9916 16448
rect 11244 16396 11296 16448
rect 16856 16396 16908 16448
rect 17776 16396 17828 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 4988 16192 5040 16244
rect 6000 16192 6052 16244
rect 6368 16192 6420 16244
rect 6460 16192 6512 16244
rect 7012 16192 7064 16244
rect 2964 16056 3016 16108
rect 5264 16056 5316 16108
rect 5816 16099 5868 16108
rect 5816 16065 5825 16099
rect 5825 16065 5859 16099
rect 5859 16065 5868 16099
rect 5816 16056 5868 16065
rect 6184 16056 6236 16108
rect 8668 16056 8720 16108
rect 9956 16056 10008 16108
rect 3608 15988 3660 16040
rect 3976 16031 4028 16040
rect 3976 15997 3985 16031
rect 3985 15997 4019 16031
rect 4019 15997 4028 16031
rect 3976 15988 4028 15997
rect 5724 15988 5776 16040
rect 6368 15988 6420 16040
rect 6920 15988 6972 16040
rect 9680 15988 9732 16040
rect 14372 16192 14424 16244
rect 14832 16192 14884 16244
rect 16488 16192 16540 16244
rect 17500 16192 17552 16244
rect 19156 16192 19208 16244
rect 19984 16192 20036 16244
rect 12900 16124 12952 16176
rect 10876 16056 10928 16108
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 13728 16056 13780 16108
rect 15292 16124 15344 16176
rect 20168 16124 20220 16176
rect 16488 16056 16540 16108
rect 18604 16099 18656 16108
rect 18604 16065 18613 16099
rect 18613 16065 18647 16099
rect 18647 16065 18656 16099
rect 18604 16056 18656 16065
rect 2596 15963 2648 15972
rect 2596 15929 2605 15963
rect 2605 15929 2639 15963
rect 2639 15929 2648 15963
rect 2596 15920 2648 15929
rect 11704 15920 11756 15972
rect 6460 15852 6512 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 8300 15852 8352 15904
rect 9220 15852 9272 15904
rect 9956 15852 10008 15904
rect 10508 15852 10560 15904
rect 10600 15852 10652 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 11428 15852 11480 15904
rect 12624 15852 12676 15904
rect 14004 15852 14056 15904
rect 14464 15963 14516 15972
rect 14464 15929 14498 15963
rect 14498 15929 14516 15963
rect 16764 15988 16816 16040
rect 17408 15988 17460 16040
rect 19248 15988 19300 16040
rect 14464 15920 14516 15929
rect 19340 15920 19392 15972
rect 15568 15852 15620 15904
rect 16672 15852 16724 15904
rect 16856 15852 16908 15904
rect 20260 15895 20312 15904
rect 20260 15861 20269 15895
rect 20269 15861 20303 15895
rect 20303 15861 20312 15895
rect 20260 15852 20312 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 6828 15648 6880 15700
rect 7104 15648 7156 15700
rect 7288 15691 7340 15700
rect 7288 15657 7297 15691
rect 7297 15657 7331 15691
rect 7331 15657 7340 15691
rect 7288 15648 7340 15657
rect 7564 15648 7616 15700
rect 10600 15691 10652 15700
rect 10600 15657 10609 15691
rect 10609 15657 10643 15691
rect 10643 15657 10652 15691
rect 10600 15648 10652 15657
rect 15200 15648 15252 15700
rect 16856 15648 16908 15700
rect 17868 15648 17920 15700
rect 19616 15648 19668 15700
rect 3332 15580 3384 15632
rect 5540 15580 5592 15632
rect 6184 15623 6236 15632
rect 6184 15589 6218 15623
rect 6218 15589 6236 15623
rect 8576 15623 8628 15632
rect 6184 15580 6236 15589
rect 8576 15589 8585 15623
rect 8585 15589 8619 15623
rect 8619 15589 8628 15623
rect 8576 15580 8628 15589
rect 8668 15580 8720 15632
rect 15844 15580 15896 15632
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 4160 15512 4212 15564
rect 5356 15512 5408 15564
rect 8208 15512 8260 15564
rect 10508 15555 10560 15564
rect 5264 15444 5316 15496
rect 2964 15376 3016 15428
rect 5448 15376 5500 15428
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 11888 15512 11940 15564
rect 14280 15512 14332 15564
rect 14464 15512 14516 15564
rect 15292 15512 15344 15564
rect 15384 15512 15436 15564
rect 17408 15580 17460 15632
rect 17776 15555 17828 15564
rect 17776 15521 17810 15555
rect 17810 15521 17828 15555
rect 17776 15512 17828 15521
rect 10600 15444 10652 15496
rect 11796 15487 11848 15496
rect 11796 15453 11805 15487
rect 11805 15453 11839 15487
rect 11839 15453 11848 15487
rect 11796 15444 11848 15453
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 16488 15487 16540 15496
rect 16488 15453 16497 15487
rect 16497 15453 16531 15487
rect 16531 15453 16540 15487
rect 17500 15487 17552 15496
rect 16488 15444 16540 15453
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 6828 15308 6880 15360
rect 7288 15308 7340 15360
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 13176 15308 13228 15317
rect 15660 15308 15712 15360
rect 16580 15308 16632 15360
rect 18788 15308 18840 15360
rect 19248 15308 19300 15360
rect 19892 15351 19944 15360
rect 19892 15317 19901 15351
rect 19901 15317 19935 15351
rect 19935 15317 19944 15351
rect 19892 15308 19944 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 5264 15104 5316 15156
rect 5724 15104 5776 15156
rect 6460 15104 6512 15156
rect 7288 15104 7340 15156
rect 11244 15104 11296 15156
rect 12624 15104 12676 15156
rect 15200 15104 15252 15156
rect 16948 15104 17000 15156
rect 20168 15104 20220 15156
rect 10600 15079 10652 15088
rect 10600 15045 10609 15079
rect 10609 15045 10643 15079
rect 10643 15045 10652 15079
rect 10600 15036 10652 15045
rect 3424 14900 3476 14952
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 7196 14968 7248 15020
rect 15292 15011 15344 15020
rect 6920 14900 6972 14952
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 9312 14900 9364 14952
rect 4068 14832 4120 14884
rect 7196 14832 7248 14884
rect 7748 14832 7800 14884
rect 10784 14900 10836 14952
rect 12348 14900 12400 14952
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 16856 15011 16908 15020
rect 16856 14977 16865 15011
rect 16865 14977 16899 15011
rect 16899 14977 16908 15011
rect 16856 14968 16908 14977
rect 4896 14764 4948 14816
rect 6460 14764 6512 14816
rect 6552 14764 6604 14816
rect 8852 14764 8904 14816
rect 9588 14832 9640 14884
rect 13176 14832 13228 14884
rect 13452 14900 13504 14952
rect 16580 14943 16632 14952
rect 16580 14909 16589 14943
rect 16589 14909 16623 14943
rect 16623 14909 16632 14943
rect 16580 14900 16632 14909
rect 17500 14900 17552 14952
rect 17868 14900 17920 14952
rect 19248 14900 19300 14952
rect 14464 14832 14516 14884
rect 14648 14832 14700 14884
rect 10876 14764 10928 14816
rect 11796 14764 11848 14816
rect 12348 14764 12400 14816
rect 12624 14764 12676 14816
rect 18696 14764 18748 14816
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 4896 14560 4948 14612
rect 5264 14560 5316 14612
rect 7104 14560 7156 14612
rect 6460 14492 6512 14544
rect 7656 14492 7708 14544
rect 7840 14492 7892 14544
rect 8484 14560 8536 14612
rect 10508 14560 10560 14612
rect 14188 14560 14240 14612
rect 15292 14560 15344 14612
rect 15844 14560 15896 14612
rect 9956 14492 10008 14544
rect 12072 14492 12124 14544
rect 12992 14492 13044 14544
rect 13176 14492 13228 14544
rect 16028 14492 16080 14544
rect 16396 14492 16448 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 4804 14399 4856 14408
rect 4804 14365 4813 14399
rect 4813 14365 4847 14399
rect 4847 14365 4856 14399
rect 4804 14356 4856 14365
rect 7288 14424 7340 14476
rect 10324 14424 10376 14476
rect 7656 14399 7708 14408
rect 7656 14365 7665 14399
rect 7665 14365 7699 14399
rect 7699 14365 7708 14399
rect 7656 14356 7708 14365
rect 7748 14356 7800 14408
rect 9864 14356 9916 14408
rect 10232 14356 10284 14408
rect 10876 14424 10928 14476
rect 11888 14424 11940 14476
rect 12808 14424 12860 14476
rect 13820 14424 13872 14476
rect 14464 14424 14516 14476
rect 14740 14424 14792 14476
rect 15292 14424 15344 14476
rect 17868 14424 17920 14476
rect 19616 14467 19668 14476
rect 19616 14433 19625 14467
rect 19625 14433 19659 14467
rect 19659 14433 19668 14467
rect 19616 14424 19668 14433
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12900 14356 12952 14408
rect 13452 14356 13504 14408
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 20168 14356 20220 14408
rect 2044 14220 2096 14272
rect 3700 14220 3752 14272
rect 10968 14288 11020 14340
rect 11060 14288 11112 14340
rect 11980 14288 12032 14340
rect 12164 14288 12216 14340
rect 15292 14288 15344 14340
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 9680 14220 9732 14272
rect 10232 14220 10284 14272
rect 10324 14220 10376 14272
rect 17132 14220 17184 14272
rect 18144 14220 18196 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 3700 14016 3752 14068
rect 1860 13991 1912 14000
rect 1860 13957 1869 13991
rect 1869 13957 1903 13991
rect 1903 13957 1912 13991
rect 1860 13948 1912 13957
rect 4068 13948 4120 14000
rect 7288 13991 7340 14000
rect 7288 13957 7297 13991
rect 7297 13957 7331 13991
rect 7331 13957 7340 13991
rect 7288 13948 7340 13957
rect 1676 13855 1728 13864
rect 1676 13821 1685 13855
rect 1685 13821 1719 13855
rect 1719 13821 1728 13855
rect 1676 13812 1728 13821
rect 2688 13812 2740 13864
rect 2872 13812 2924 13864
rect 3884 13744 3936 13796
rect 6184 13880 6236 13932
rect 8208 13948 8260 14000
rect 9036 13880 9088 13932
rect 6828 13812 6880 13864
rect 6920 13812 6972 13864
rect 9864 14016 9916 14068
rect 12072 14016 12124 14068
rect 18788 14016 18840 14068
rect 20076 14016 20128 14068
rect 12900 13948 12952 14000
rect 16396 13948 16448 14000
rect 10692 13880 10744 13932
rect 13728 13880 13780 13932
rect 14556 13880 14608 13932
rect 15200 13880 15252 13932
rect 18788 13923 18840 13932
rect 4804 13744 4856 13796
rect 7840 13744 7892 13796
rect 8852 13744 8904 13796
rect 9588 13744 9640 13796
rect 10416 13812 10468 13864
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 11704 13812 11756 13864
rect 12992 13855 13044 13864
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 14464 13812 14516 13864
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 18788 13889 18797 13923
rect 18797 13889 18831 13923
rect 18831 13889 18840 13923
rect 18788 13880 18840 13889
rect 19248 13880 19300 13932
rect 16304 13812 16356 13864
rect 19524 13812 19576 13864
rect 19984 13812 20036 13864
rect 3792 13676 3844 13728
rect 5540 13676 5592 13728
rect 6552 13676 6604 13728
rect 8760 13676 8812 13728
rect 9312 13676 9364 13728
rect 10508 13676 10560 13728
rect 10876 13676 10928 13728
rect 11336 13676 11388 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 15660 13676 15712 13728
rect 16304 13676 16356 13728
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 19248 13676 19300 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 1400 13515 1452 13524
rect 1400 13481 1409 13515
rect 1409 13481 1443 13515
rect 1443 13481 1452 13515
rect 1400 13472 1452 13481
rect 2872 13472 2924 13524
rect 3056 13472 3108 13524
rect 2504 13404 2556 13456
rect 8300 13472 8352 13524
rect 8484 13472 8536 13524
rect 1768 13336 1820 13388
rect 6460 13404 6512 13456
rect 4252 13336 4304 13388
rect 5540 13336 5592 13388
rect 7748 13336 7800 13388
rect 2780 13268 2832 13320
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 5264 13268 5316 13320
rect 5172 13132 5224 13184
rect 5448 13132 5500 13184
rect 7472 13268 7524 13320
rect 7012 13200 7064 13252
rect 9404 13404 9456 13456
rect 9956 13472 10008 13524
rect 10324 13472 10376 13524
rect 12624 13472 12676 13524
rect 13636 13404 13688 13456
rect 14740 13472 14792 13524
rect 18236 13472 18288 13524
rect 19708 13472 19760 13524
rect 15844 13404 15896 13456
rect 16028 13404 16080 13456
rect 19340 13404 19392 13456
rect 9036 13336 9088 13388
rect 9588 13336 9640 13388
rect 10692 13336 10744 13388
rect 11796 13336 11848 13388
rect 11980 13336 12032 13388
rect 14740 13336 14792 13388
rect 15660 13379 15712 13388
rect 15660 13345 15669 13379
rect 15669 13345 15703 13379
rect 15703 13345 15712 13379
rect 15660 13336 15712 13345
rect 16580 13336 16632 13388
rect 19524 13336 19576 13388
rect 20536 13336 20588 13388
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 9680 13268 9732 13320
rect 9864 13268 9916 13320
rect 12348 13268 12400 13320
rect 8024 13175 8076 13184
rect 8024 13141 8033 13175
rect 8033 13141 8067 13175
rect 8067 13141 8076 13175
rect 8024 13132 8076 13141
rect 9128 13200 9180 13252
rect 13452 13200 13504 13252
rect 16396 13268 16448 13320
rect 19340 13268 19392 13320
rect 19432 13268 19484 13320
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 16028 13200 16080 13252
rect 17592 13200 17644 13252
rect 12164 13132 12216 13184
rect 12624 13132 12676 13184
rect 14096 13132 14148 13184
rect 15200 13132 15252 13184
rect 17500 13132 17552 13184
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 6828 12971 6880 12980
rect 6828 12937 6837 12971
rect 6837 12937 6871 12971
rect 6871 12937 6880 12971
rect 6828 12928 6880 12937
rect 7104 12928 7156 12980
rect 7288 12928 7340 12980
rect 8024 12928 8076 12980
rect 12440 12928 12492 12980
rect 3884 12903 3936 12912
rect 3884 12869 3893 12903
rect 3893 12869 3927 12903
rect 3927 12869 3936 12903
rect 3884 12860 3936 12869
rect 5172 12835 5224 12844
rect 5172 12801 5181 12835
rect 5181 12801 5215 12835
rect 5215 12801 5224 12835
rect 5172 12792 5224 12801
rect 5540 12860 5592 12912
rect 5724 12860 5776 12912
rect 6736 12860 6788 12912
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 7748 12792 7800 12844
rect 9312 12792 9364 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 3056 12724 3108 12776
rect 4528 12724 4580 12776
rect 6368 12724 6420 12776
rect 11152 12860 11204 12912
rect 11704 12860 11756 12912
rect 12164 12860 12216 12912
rect 12348 12860 12400 12912
rect 15108 12928 15160 12980
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 19156 12928 19208 12980
rect 19340 12928 19392 12980
rect 19708 12928 19760 12980
rect 2688 12656 2740 12708
rect 3240 12656 3292 12708
rect 3608 12656 3660 12708
rect 3884 12656 3936 12708
rect 8116 12656 8168 12708
rect 8208 12656 8260 12708
rect 9496 12656 9548 12708
rect 4160 12588 4212 12640
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 7104 12588 7156 12640
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 7472 12588 7524 12640
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 8760 12588 8812 12597
rect 10324 12631 10376 12640
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 12900 12792 12952 12844
rect 13360 12792 13412 12844
rect 13544 12792 13596 12844
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 18788 12792 18840 12844
rect 17316 12724 17368 12776
rect 17868 12724 17920 12776
rect 19248 12767 19300 12776
rect 19248 12733 19271 12767
rect 19271 12733 19300 12767
rect 19248 12724 19300 12733
rect 12900 12656 12952 12708
rect 13268 12656 13320 12708
rect 13636 12656 13688 12708
rect 15568 12656 15620 12708
rect 16120 12656 16172 12708
rect 18696 12656 18748 12708
rect 11796 12588 11848 12640
rect 12532 12588 12584 12640
rect 15292 12588 15344 12640
rect 17408 12588 17460 12640
rect 17960 12588 18012 12640
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 4804 12384 4856 12436
rect 5448 12384 5500 12436
rect 7656 12384 7708 12436
rect 7748 12384 7800 12436
rect 10508 12384 10560 12436
rect 14188 12384 14240 12436
rect 15200 12384 15252 12436
rect 15384 12384 15436 12436
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 5448 12248 5500 12300
rect 5724 12248 5776 12300
rect 6828 12248 6880 12300
rect 8208 12248 8260 12300
rect 8668 12248 8720 12300
rect 8944 12248 8996 12300
rect 9128 12291 9180 12300
rect 9128 12257 9137 12291
rect 9137 12257 9171 12291
rect 9171 12257 9180 12291
rect 9128 12248 9180 12257
rect 9864 12248 9916 12300
rect 3056 12155 3108 12164
rect 3056 12121 3065 12155
rect 3065 12121 3099 12155
rect 3099 12121 3108 12155
rect 3056 12112 3108 12121
rect 4528 12112 4580 12164
rect 10692 12180 10744 12232
rect 12164 12316 12216 12368
rect 13728 12316 13780 12368
rect 13820 12316 13872 12368
rect 14372 12316 14424 12368
rect 14648 12316 14700 12368
rect 18052 12384 18104 12436
rect 19248 12427 19300 12436
rect 19248 12393 19257 12427
rect 19257 12393 19291 12427
rect 19291 12393 19300 12427
rect 19248 12384 19300 12393
rect 13452 12248 13504 12300
rect 5540 12112 5592 12164
rect 7748 12112 7800 12164
rect 9864 12112 9916 12164
rect 10048 12112 10100 12164
rect 5172 12044 5224 12096
rect 8668 12044 8720 12096
rect 9036 12044 9088 12096
rect 12164 12180 12216 12232
rect 12624 12180 12676 12232
rect 19432 12316 19484 12368
rect 11980 12112 12032 12164
rect 12532 12112 12584 12164
rect 17132 12248 17184 12300
rect 17868 12291 17920 12300
rect 17868 12257 17877 12291
rect 17877 12257 17911 12291
rect 17911 12257 17920 12291
rect 17868 12248 17920 12257
rect 17960 12248 18012 12300
rect 16580 12180 16632 12232
rect 14280 12044 14332 12096
rect 14740 12087 14792 12096
rect 14740 12053 14749 12087
rect 14749 12053 14783 12087
rect 14783 12053 14792 12087
rect 14740 12044 14792 12053
rect 18972 12112 19024 12164
rect 20352 12112 20404 12164
rect 19800 12044 19852 12096
rect 20628 12044 20680 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 4252 11840 4304 11892
rect 5080 11883 5132 11892
rect 5080 11849 5089 11883
rect 5089 11849 5123 11883
rect 5123 11849 5132 11883
rect 5080 11840 5132 11849
rect 8208 11883 8260 11892
rect 8208 11849 8217 11883
rect 8217 11849 8251 11883
rect 8251 11849 8260 11883
rect 8208 11840 8260 11849
rect 8760 11840 8812 11892
rect 9404 11840 9456 11892
rect 8392 11772 8444 11824
rect 2964 11704 3016 11756
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 5540 11704 5592 11756
rect 6828 11747 6880 11756
rect 6828 11713 6837 11747
rect 6837 11713 6871 11747
rect 6871 11713 6880 11747
rect 6828 11704 6880 11713
rect 8208 11704 8260 11756
rect 10048 11772 10100 11824
rect 10324 11840 10376 11892
rect 10692 11840 10744 11892
rect 12808 11840 12860 11892
rect 12992 11840 13044 11892
rect 15108 11840 15160 11892
rect 13820 11772 13872 11824
rect 20628 11840 20680 11892
rect 9496 11704 9548 11756
rect 10324 11704 10376 11756
rect 11704 11704 11756 11756
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 17960 11772 18012 11824
rect 17132 11704 17184 11756
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 3792 11636 3844 11688
rect 4160 11636 4212 11688
rect 4252 11636 4304 11688
rect 8760 11636 8812 11688
rect 9312 11636 9364 11688
rect 4160 11500 4212 11552
rect 4804 11500 4856 11552
rect 5080 11500 5132 11552
rect 6644 11568 6696 11620
rect 8484 11568 8536 11620
rect 10048 11636 10100 11688
rect 10416 11636 10468 11688
rect 11060 11679 11112 11688
rect 11060 11645 11069 11679
rect 11069 11645 11103 11679
rect 11103 11645 11112 11679
rect 11060 11636 11112 11645
rect 18144 11679 18196 11688
rect 5632 11500 5684 11552
rect 8208 11500 8260 11552
rect 8300 11500 8352 11552
rect 10692 11568 10744 11620
rect 8760 11500 8812 11552
rect 11888 11500 11940 11552
rect 12532 11500 12584 11552
rect 16028 11568 16080 11620
rect 12992 11500 13044 11552
rect 17776 11568 17828 11620
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 19248 11636 19300 11688
rect 19708 11679 19760 11688
rect 19708 11645 19742 11679
rect 19742 11645 19760 11679
rect 19708 11636 19760 11645
rect 18972 11568 19024 11620
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 17592 11500 17644 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 4252 11296 4304 11348
rect 4436 11339 4488 11348
rect 4436 11305 4445 11339
rect 4445 11305 4479 11339
rect 4479 11305 4488 11339
rect 4436 11296 4488 11305
rect 6184 11296 6236 11348
rect 6276 11296 6328 11348
rect 8392 11296 8444 11348
rect 8484 11296 8536 11348
rect 9404 11296 9456 11348
rect 10048 11296 10100 11348
rect 7196 11228 7248 11280
rect 5172 11160 5224 11212
rect 5264 11092 5316 11144
rect 5816 11092 5868 11144
rect 4896 11024 4948 11076
rect 6368 11024 6420 11076
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 8576 11228 8628 11280
rect 8944 11228 8996 11280
rect 9588 11160 9640 11212
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 11244 11296 11296 11348
rect 11980 11296 12032 11348
rect 12624 11296 12676 11348
rect 13452 11339 13504 11348
rect 13452 11305 13461 11339
rect 13461 11305 13495 11339
rect 13495 11305 13504 11339
rect 13452 11296 13504 11305
rect 14556 11296 14608 11348
rect 16672 11296 16724 11348
rect 10876 11271 10928 11280
rect 9680 11160 9732 11169
rect 8208 11092 8260 11144
rect 8576 11092 8628 11144
rect 10508 11160 10560 11212
rect 10876 11237 10885 11271
rect 10885 11237 10919 11271
rect 10919 11237 10928 11271
rect 10876 11228 10928 11237
rect 11612 11228 11664 11280
rect 11888 11228 11940 11280
rect 13268 11228 13320 11280
rect 16856 11228 16908 11280
rect 17960 11296 18012 11348
rect 19524 11296 19576 11348
rect 11060 11160 11112 11212
rect 14280 11160 14332 11212
rect 15660 11160 15712 11212
rect 18144 11160 18196 11212
rect 7932 11024 7984 11076
rect 13728 11092 13780 11144
rect 14372 11092 14424 11144
rect 15384 11092 15436 11144
rect 15936 11135 15988 11144
rect 15936 11101 15945 11135
rect 15945 11101 15979 11135
rect 15979 11101 15988 11135
rect 16948 11135 17000 11144
rect 15936 11092 15988 11101
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 18052 11092 18104 11144
rect 18788 11092 18840 11144
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 296 10956 348 11008
rect 6920 10956 6972 11008
rect 8208 10956 8260 11008
rect 10324 10956 10376 11008
rect 14188 10956 14240 11008
rect 18696 11024 18748 11076
rect 19616 11024 19668 11076
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 7196 10752 7248 10804
rect 5816 10727 5868 10736
rect 5816 10693 5825 10727
rect 5825 10693 5859 10727
rect 5859 10693 5868 10727
rect 5816 10684 5868 10693
rect 9404 10752 9456 10804
rect 10692 10684 10744 10736
rect 12164 10727 12216 10736
rect 12164 10693 12173 10727
rect 12173 10693 12207 10727
rect 12207 10693 12216 10727
rect 12164 10684 12216 10693
rect 13728 10752 13780 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 16948 10752 17000 10804
rect 17408 10684 17460 10736
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 9220 10616 9272 10668
rect 3884 10548 3936 10600
rect 4620 10523 4672 10532
rect 4620 10489 4629 10523
rect 4629 10489 4663 10523
rect 4663 10489 4672 10523
rect 4620 10480 4672 10489
rect 6736 10548 6788 10600
rect 7104 10523 7156 10532
rect 7104 10489 7113 10523
rect 7113 10489 7147 10523
rect 7147 10489 7156 10523
rect 7104 10480 7156 10489
rect 7196 10412 7248 10464
rect 8208 10548 8260 10600
rect 18880 10752 18932 10804
rect 19340 10752 19392 10804
rect 19156 10659 19208 10668
rect 19156 10625 19165 10659
rect 19165 10625 19199 10659
rect 19199 10625 19208 10659
rect 19156 10616 19208 10625
rect 15292 10548 15344 10600
rect 11060 10523 11112 10532
rect 9128 10412 9180 10464
rect 9680 10412 9732 10464
rect 9956 10412 10008 10464
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 11060 10489 11094 10523
rect 11094 10489 11112 10523
rect 11060 10480 11112 10489
rect 11336 10480 11388 10532
rect 16488 10548 16540 10600
rect 17868 10591 17920 10600
rect 17868 10557 17877 10591
rect 17877 10557 17911 10591
rect 17911 10557 17920 10591
rect 17868 10548 17920 10557
rect 16948 10480 17000 10532
rect 17132 10480 17184 10532
rect 19892 10480 19944 10532
rect 20444 10480 20496 10532
rect 20168 10412 20220 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 4804 10251 4856 10260
rect 4804 10217 4813 10251
rect 4813 10217 4847 10251
rect 4847 10217 4856 10251
rect 4804 10208 4856 10217
rect 6828 10208 6880 10260
rect 8208 10208 8260 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 8576 10208 8628 10260
rect 10048 10208 10100 10260
rect 10324 10208 10376 10260
rect 12716 10208 12768 10260
rect 16580 10208 16632 10260
rect 19524 10208 19576 10260
rect 7104 10140 7156 10192
rect 7564 10072 7616 10124
rect 8484 10004 8536 10056
rect 5356 9936 5408 9988
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 13360 10072 13412 10124
rect 14740 10072 14792 10124
rect 15936 10140 15988 10192
rect 16396 10140 16448 10192
rect 17500 10115 17552 10124
rect 9128 10004 9180 10056
rect 10968 10004 11020 10056
rect 7104 9911 7156 9920
rect 7104 9877 7113 9911
rect 7113 9877 7147 9911
rect 7147 9877 7156 9911
rect 7104 9868 7156 9877
rect 9680 9936 9732 9988
rect 11336 9979 11388 9988
rect 11336 9945 11345 9979
rect 11345 9945 11379 9979
rect 11379 9945 11388 9979
rect 11336 9936 11388 9945
rect 12440 10004 12492 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 16488 9936 16540 9988
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 17960 9936 18012 9988
rect 19340 10047 19392 10056
rect 19340 10013 19349 10047
rect 19349 10013 19383 10047
rect 19383 10013 19392 10047
rect 19340 10004 19392 10013
rect 19248 9936 19300 9988
rect 12164 9868 12216 9920
rect 17408 9868 17460 9920
rect 17868 9868 17920 9920
rect 18788 9911 18840 9920
rect 18788 9877 18797 9911
rect 18797 9877 18831 9911
rect 18831 9877 18840 9911
rect 18788 9868 18840 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 3516 9664 3568 9716
rect 8484 9596 8536 9648
rect 8760 9596 8812 9648
rect 6000 9528 6052 9580
rect 10968 9664 11020 9716
rect 19340 9664 19392 9716
rect 6644 9460 6696 9512
rect 4804 9392 4856 9444
rect 7748 9392 7800 9444
rect 8300 9460 8352 9512
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 9220 9460 9272 9512
rect 11980 9528 12032 9580
rect 12900 9596 12952 9648
rect 12992 9596 13044 9648
rect 13268 9528 13320 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 15476 9596 15528 9648
rect 18604 9596 18656 9648
rect 20444 9596 20496 9648
rect 15752 9571 15804 9580
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 9588 9392 9640 9444
rect 8300 9367 8352 9376
rect 8300 9333 8309 9367
rect 8309 9333 8343 9367
rect 8343 9333 8352 9367
rect 8300 9324 8352 9333
rect 8852 9324 8904 9376
rect 9496 9324 9548 9376
rect 10692 9392 10744 9444
rect 14556 9460 14608 9512
rect 14740 9460 14792 9512
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 17684 9528 17736 9580
rect 19156 9528 19208 9580
rect 17960 9460 18012 9512
rect 13452 9324 13504 9376
rect 13544 9367 13596 9376
rect 13544 9333 13553 9367
rect 13553 9333 13587 9367
rect 13587 9333 13596 9367
rect 13544 9324 13596 9333
rect 14096 9324 14148 9376
rect 14556 9324 14608 9376
rect 15292 9324 15344 9376
rect 15384 9324 15436 9376
rect 15660 9392 15712 9444
rect 19800 9392 19852 9444
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 4896 9120 4948 9172
rect 7748 9120 7800 9172
rect 8208 9120 8260 9172
rect 12992 9120 13044 9172
rect 15384 9120 15436 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 17776 9120 17828 9172
rect 19340 9163 19392 9172
rect 6644 9027 6696 9036
rect 6644 8993 6653 9027
rect 6653 8993 6687 9027
rect 6687 8993 6696 9027
rect 6644 8984 6696 8993
rect 7656 8984 7708 9036
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 9128 8984 9180 9036
rect 11244 8984 11296 9036
rect 14004 9027 14056 9036
rect 14004 8993 14013 9027
rect 14013 8993 14047 9027
rect 14047 8993 14056 9027
rect 14004 8984 14056 8993
rect 10140 8916 10192 8968
rect 11704 8916 11756 8968
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 17040 9052 17092 9104
rect 19340 9129 19349 9163
rect 19349 9129 19383 9163
rect 19383 9129 19392 9163
rect 19340 9120 19392 9129
rect 19156 8984 19208 9036
rect 14188 8916 14240 8925
rect 2872 8780 2924 8832
rect 10692 8848 10744 8900
rect 8576 8780 8628 8832
rect 9864 8780 9916 8832
rect 13820 8848 13872 8900
rect 13912 8848 13964 8900
rect 17684 8916 17736 8968
rect 17868 8848 17920 8900
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 14004 8780 14056 8832
rect 17776 8780 17828 8832
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 15660 8576 15712 8628
rect 15752 8576 15804 8628
rect 16120 8576 16172 8628
rect 12348 8508 12400 8560
rect 14188 8551 14240 8560
rect 14188 8517 14197 8551
rect 14197 8517 14231 8551
rect 14231 8517 14240 8551
rect 14188 8508 14240 8517
rect 16764 8508 16816 8560
rect 18236 8508 18288 8560
rect 19524 8508 19576 8560
rect 2412 8440 2464 8492
rect 7012 8440 7064 8492
rect 7748 8440 7800 8492
rect 7656 8372 7708 8424
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 10324 8372 10376 8424
rect 11888 8372 11940 8424
rect 16304 8440 16356 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20628 8483 20680 8492
rect 20628 8449 20637 8483
rect 20637 8449 20671 8483
rect 20671 8449 20680 8483
rect 20628 8440 20680 8449
rect 5632 8304 5684 8356
rect 8208 8304 8260 8356
rect 12072 8304 12124 8356
rect 15660 8372 15712 8424
rect 17224 8372 17276 8424
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 18144 8372 18196 8424
rect 16764 8304 16816 8356
rect 18604 8304 18656 8356
rect 19892 8347 19944 8356
rect 19892 8313 19901 8347
rect 19901 8313 19935 8347
rect 19935 8313 19944 8347
rect 19892 8304 19944 8313
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 8300 8279 8352 8288
rect 8300 8245 8309 8279
rect 8309 8245 8343 8279
rect 8343 8245 8352 8279
rect 8300 8236 8352 8245
rect 10692 8236 10744 8288
rect 10784 8236 10836 8288
rect 17500 8236 17552 8288
rect 18052 8279 18104 8288
rect 18052 8245 18061 8279
rect 18061 8245 18095 8279
rect 18095 8245 18104 8279
rect 18052 8236 18104 8245
rect 20076 8279 20128 8288
rect 20076 8245 20085 8279
rect 20085 8245 20119 8279
rect 20119 8245 20128 8279
rect 20076 8236 20128 8245
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 4436 8075 4488 8084
rect 4436 8041 4445 8075
rect 4445 8041 4479 8075
rect 4479 8041 4488 8075
rect 4436 8032 4488 8041
rect 6644 7964 6696 8016
rect 6920 8032 6972 8084
rect 8484 8032 8536 8084
rect 9036 8032 9088 8084
rect 9128 8032 9180 8084
rect 9864 8032 9916 8084
rect 10048 8032 10100 8084
rect 18052 8032 18104 8084
rect 19248 8032 19300 8084
rect 8208 7964 8260 8016
rect 16028 8007 16080 8016
rect 16028 7973 16037 8007
rect 16037 7973 16071 8007
rect 16071 7973 16080 8007
rect 16028 7964 16080 7973
rect 17960 7964 18012 8016
rect 6920 7896 6972 7948
rect 7656 7896 7708 7948
rect 7748 7828 7800 7880
rect 8576 7896 8628 7948
rect 10048 7939 10100 7948
rect 10048 7905 10082 7939
rect 10082 7905 10100 7939
rect 10048 7896 10100 7905
rect 12348 7939 12400 7948
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 18696 7896 18748 7948
rect 8484 7828 8536 7880
rect 9128 7828 9180 7880
rect 12072 7828 12124 7880
rect 13176 7828 13228 7880
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 17684 7871 17736 7880
rect 16120 7828 16172 7837
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 8300 7760 8352 7812
rect 11060 7760 11112 7812
rect 14648 7760 14700 7812
rect 15660 7760 15712 7812
rect 18328 7760 18380 7812
rect 4344 7692 4396 7744
rect 9404 7692 9456 7744
rect 11244 7692 11296 7744
rect 11704 7692 11756 7744
rect 11888 7692 11940 7744
rect 15936 7692 15988 7744
rect 17960 7692 18012 7744
rect 19248 7871 19300 7880
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 19156 7760 19208 7812
rect 19248 7692 19300 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 3148 7488 3200 7540
rect 5448 7488 5500 7540
rect 6644 7488 6696 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 12348 7488 12400 7540
rect 12992 7488 13044 7540
rect 5632 7420 5684 7472
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 10048 7420 10100 7472
rect 12624 7420 12676 7472
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 5448 7327 5500 7336
rect 5448 7293 5457 7327
rect 5457 7293 5491 7327
rect 5491 7293 5500 7327
rect 5448 7284 5500 7293
rect 6828 7327 6880 7336
rect 3056 7216 3108 7268
rect 3332 7216 3384 7268
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 11060 7352 11112 7404
rect 11704 7352 11756 7404
rect 14096 7352 14148 7404
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 16304 7420 16356 7472
rect 19156 7488 19208 7540
rect 19340 7420 19392 7472
rect 15292 7352 15344 7404
rect 16488 7352 16540 7404
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 14004 7284 14056 7336
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 19984 7284 20036 7336
rect 20536 7327 20588 7336
rect 20536 7293 20545 7327
rect 20545 7293 20579 7327
rect 20579 7293 20588 7327
rect 20536 7284 20588 7293
rect 8576 7216 8628 7268
rect 8760 7259 8812 7268
rect 8760 7225 8794 7259
rect 8794 7225 8812 7259
rect 8760 7216 8812 7225
rect 17684 7216 17736 7268
rect 19064 7216 19116 7268
rect 6920 7148 6972 7200
rect 8668 7148 8720 7200
rect 11244 7148 11296 7200
rect 12808 7148 12860 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 21548 7148 21600 7200
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 6828 6944 6880 6996
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 11244 6944 11296 6996
rect 13176 6944 13228 6996
rect 14280 6944 14332 6996
rect 7564 6876 7616 6928
rect 6920 6808 6972 6860
rect 11060 6876 11112 6928
rect 11152 6876 11204 6928
rect 12348 6876 12400 6928
rect 12808 6876 12860 6928
rect 13084 6876 13136 6928
rect 13728 6876 13780 6928
rect 14004 6919 14056 6928
rect 14004 6885 14013 6919
rect 14013 6885 14047 6919
rect 14047 6885 14056 6919
rect 14004 6876 14056 6885
rect 16120 6876 16172 6928
rect 5724 6740 5776 6792
rect 7656 6740 7708 6792
rect 10876 6808 10928 6860
rect 1952 6672 2004 6724
rect 2504 6672 2556 6724
rect 8484 6740 8536 6792
rect 11152 6740 11204 6792
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 10508 6715 10560 6724
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 12716 6672 12768 6724
rect 15200 6808 15252 6860
rect 16764 6808 16816 6860
rect 18052 6876 18104 6928
rect 18696 6876 18748 6928
rect 20628 6808 20680 6860
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 2688 6604 2740 6656
rect 3700 6604 3752 6656
rect 11152 6604 11204 6656
rect 14188 6604 14240 6656
rect 17132 6672 17184 6724
rect 17592 6672 17644 6724
rect 16488 6604 16540 6656
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 5172 6400 5224 6452
rect 8944 6400 8996 6452
rect 14188 6400 14240 6452
rect 14280 6400 14332 6452
rect 12440 6332 12492 6384
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 6276 6264 6328 6316
rect 6644 6264 6696 6316
rect 9128 6264 9180 6316
rect 10508 6264 10560 6316
rect 9220 6196 9272 6248
rect 10876 6196 10928 6248
rect 14464 6264 14516 6316
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 17592 6264 17644 6316
rect 19892 6264 19944 6316
rect 20628 6264 20680 6316
rect 7656 6128 7708 6180
rect 8300 6128 8352 6180
rect 2964 6060 3016 6112
rect 4804 6060 4856 6112
rect 7748 6060 7800 6112
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8392 6060 8444 6112
rect 13912 6128 13964 6180
rect 14188 6196 14240 6248
rect 14372 6196 14424 6248
rect 16488 6196 16540 6248
rect 17500 6196 17552 6248
rect 16856 6128 16908 6180
rect 12072 6060 12124 6112
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 16488 6060 16540 6112
rect 19708 6103 19760 6112
rect 19708 6069 19717 6103
rect 19717 6069 19751 6103
rect 19751 6069 19760 6103
rect 19708 6060 19760 6069
rect 19800 6060 19852 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2964 5899 3016 5908
rect 2964 5865 2973 5899
rect 2973 5865 3007 5899
rect 3007 5865 3016 5899
rect 2964 5856 3016 5865
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 4344 5763 4396 5772
rect 4344 5729 4378 5763
rect 4378 5729 4396 5763
rect 4344 5720 4396 5729
rect 5448 5788 5500 5840
rect 9220 5856 9272 5908
rect 12716 5856 12768 5908
rect 12808 5856 12860 5908
rect 14740 5856 14792 5908
rect 19800 5856 19852 5908
rect 14372 5788 14424 5840
rect 17776 5788 17828 5840
rect 18880 5788 18932 5840
rect 8300 5720 8352 5772
rect 8484 5763 8536 5772
rect 8484 5729 8493 5763
rect 8493 5729 8527 5763
rect 8527 5729 8536 5763
rect 8484 5720 8536 5729
rect 9128 5720 9180 5772
rect 9680 5763 9732 5772
rect 9680 5729 9689 5763
rect 9689 5729 9723 5763
rect 9723 5729 9732 5763
rect 9680 5720 9732 5729
rect 6276 5695 6328 5704
rect 3148 5516 3200 5568
rect 3332 5516 3384 5568
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 14556 5720 14608 5772
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 13912 5695 13964 5704
rect 12440 5652 12492 5661
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 14280 5652 14332 5704
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 18144 5652 18196 5704
rect 19892 5695 19944 5704
rect 5448 5627 5500 5636
rect 5448 5593 5457 5627
rect 5457 5593 5491 5627
rect 5491 5593 5500 5627
rect 5448 5584 5500 5593
rect 6276 5516 6328 5568
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 11152 5516 11204 5568
rect 19616 5584 19668 5636
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 19984 5584 20036 5636
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18144 5516 18196 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 3332 5312 3384 5364
rect 4160 5312 4212 5364
rect 4344 5312 4396 5364
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 13912 5312 13964 5364
rect 18052 5312 18104 5364
rect 4896 5244 4948 5296
rect 5356 5244 5408 5296
rect 14556 5244 14608 5296
rect 20444 5312 20496 5364
rect 20628 5312 20680 5364
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 6276 5176 6328 5228
rect 6736 5176 6788 5228
rect 8668 5176 8720 5228
rect 9036 5176 9088 5228
rect 11060 5176 11112 5228
rect 14188 5219 14240 5228
rect 14188 5185 14197 5219
rect 14197 5185 14231 5219
rect 14231 5185 14240 5219
rect 14188 5176 14240 5185
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 18696 5176 18748 5228
rect 4160 5040 4212 5092
rect 7472 5108 7524 5160
rect 8208 5108 8260 5160
rect 9404 5108 9456 5160
rect 10784 5108 10836 5160
rect 11152 5151 11204 5160
rect 11152 5117 11161 5151
rect 11161 5117 11195 5151
rect 11195 5117 11204 5151
rect 11152 5108 11204 5117
rect 12072 5108 12124 5160
rect 12992 5108 13044 5160
rect 13728 5108 13780 5160
rect 15660 5151 15712 5160
rect 9036 5040 9088 5092
rect 15660 5117 15669 5151
rect 15669 5117 15703 5151
rect 15703 5117 15712 5151
rect 15660 5108 15712 5117
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 8208 4972 8260 5024
rect 10692 4972 10744 5024
rect 16212 5040 16264 5092
rect 19892 5040 19944 5092
rect 12624 4972 12676 5024
rect 13912 4972 13964 5024
rect 14004 4972 14056 5024
rect 14280 4972 14332 5024
rect 15752 5015 15804 5024
rect 15752 4981 15761 5015
rect 15761 4981 15795 5015
rect 15795 4981 15804 5015
rect 15752 4972 15804 4981
rect 18052 4972 18104 5024
rect 20260 4972 20312 5024
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 4804 4768 4856 4820
rect 5724 4768 5776 4820
rect 9036 4768 9088 4820
rect 2136 4700 2188 4752
rect 6368 4700 6420 4752
rect 6552 4700 6604 4752
rect 7748 4700 7800 4752
rect 11060 4700 11112 4752
rect 12532 4768 12584 4820
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 16212 4768 16264 4820
rect 13820 4700 13872 4752
rect 14280 4700 14332 4752
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 4252 4632 4304 4684
rect 5540 4632 5592 4684
rect 4160 4564 4212 4616
rect 4896 4496 4948 4548
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 7472 4564 7524 4616
rect 6920 4496 6972 4548
rect 4988 4428 5040 4480
rect 18144 4700 18196 4752
rect 18604 4700 18656 4752
rect 20536 4632 20588 4684
rect 8760 4564 8812 4616
rect 9680 4564 9732 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 9772 4496 9824 4548
rect 12532 4496 12584 4548
rect 14188 4496 14240 4548
rect 17776 4564 17828 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 8484 4428 8536 4480
rect 9864 4428 9916 4480
rect 11152 4428 11204 4480
rect 14096 4428 14148 4480
rect 18144 4428 18196 4480
rect 19708 4428 19760 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 3148 4224 3200 4276
rect 4160 4267 4212 4276
rect 4160 4233 4169 4267
rect 4169 4233 4203 4267
rect 4203 4233 4212 4267
rect 4160 4224 4212 4233
rect 6368 4224 6420 4276
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 8484 4088 8536 4140
rect 5816 4020 5868 4072
rect 7472 4063 7524 4072
rect 7472 4029 7481 4063
rect 7481 4029 7515 4063
rect 7515 4029 7524 4063
rect 7472 4020 7524 4029
rect 10600 4156 10652 4208
rect 14280 4156 14332 4208
rect 14740 4156 14792 4208
rect 13912 4088 13964 4140
rect 848 3952 900 4004
rect 3240 3952 3292 4004
rect 5724 3952 5776 4004
rect 9680 4020 9732 4072
rect 10876 4020 10928 4072
rect 11980 4020 12032 4072
rect 5172 3927 5224 3936
rect 5172 3893 5181 3927
rect 5181 3893 5215 3927
rect 5215 3893 5224 3927
rect 5172 3884 5224 3893
rect 5356 3884 5408 3936
rect 5908 3884 5960 3936
rect 6644 3884 6696 3936
rect 9496 3952 9548 4004
rect 7748 3884 7800 3936
rect 10600 3952 10652 4004
rect 10692 3952 10744 4004
rect 12532 4020 12584 4072
rect 14280 4020 14332 4072
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10232 3884 10284 3936
rect 11244 3884 11296 3936
rect 14004 3884 14056 3936
rect 14740 3884 14792 3936
rect 15752 4020 15804 4072
rect 16764 4020 16816 4072
rect 17500 4020 17552 4072
rect 19708 4063 19760 4072
rect 19708 4029 19731 4063
rect 19731 4029 19760 4063
rect 19708 4020 19760 4029
rect 16580 3884 16632 3936
rect 16764 3927 16816 3936
rect 16764 3893 16773 3927
rect 16773 3893 16807 3927
rect 16807 3893 16816 3927
rect 16764 3884 16816 3893
rect 18052 3884 18104 3936
rect 22652 3952 22704 4004
rect 19892 3884 19944 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 3240 3680 3292 3732
rect 5540 3680 5592 3732
rect 5816 3723 5868 3732
rect 5816 3689 5825 3723
rect 5825 3689 5859 3723
rect 5859 3689 5868 3723
rect 5816 3680 5868 3689
rect 5908 3680 5960 3732
rect 9588 3680 9640 3732
rect 9772 3680 9824 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 14372 3680 14424 3732
rect 15384 3680 15436 3732
rect 15476 3680 15528 3732
rect 2688 3544 2740 3596
rect 5448 3544 5500 3596
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 6828 3544 6880 3596
rect 9772 3544 9824 3596
rect 9956 3587 10008 3596
rect 9956 3553 9990 3587
rect 9990 3553 10008 3587
rect 9956 3544 10008 3553
rect 10324 3544 10376 3596
rect 296 3476 348 3528
rect 1400 3408 1452 3460
rect 4252 3408 4304 3460
rect 2872 3340 2924 3392
rect 3056 3383 3108 3392
rect 3056 3349 3065 3383
rect 3065 3349 3099 3383
rect 3099 3349 3108 3383
rect 3056 3340 3108 3349
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 5816 3476 5868 3528
rect 8300 3476 8352 3528
rect 9312 3476 9364 3528
rect 9496 3476 9548 3528
rect 11152 3612 11204 3664
rect 16764 3680 16816 3732
rect 19248 3680 19300 3732
rect 11888 3587 11940 3596
rect 11888 3553 11897 3587
rect 11897 3553 11931 3587
rect 11931 3553 11940 3587
rect 11888 3544 11940 3553
rect 7748 3340 7800 3392
rect 13912 3544 13964 3596
rect 14004 3544 14056 3596
rect 15660 3544 15712 3596
rect 16396 3544 16448 3596
rect 18696 3544 18748 3596
rect 18788 3544 18840 3596
rect 20260 3544 20312 3596
rect 22100 3544 22152 3596
rect 14464 3476 14516 3528
rect 15476 3476 15528 3528
rect 15752 3519 15804 3528
rect 15752 3485 15761 3519
rect 15761 3485 15795 3519
rect 15795 3485 15804 3519
rect 15752 3476 15804 3485
rect 14832 3408 14884 3460
rect 17776 3476 17828 3528
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 17868 3408 17920 3460
rect 13912 3340 13964 3392
rect 14004 3340 14056 3392
rect 17040 3340 17092 3392
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 5448 3179 5500 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 5448 3145 5457 3179
rect 5457 3145 5491 3179
rect 5491 3145 5500 3179
rect 5448 3136 5500 3145
rect 2964 2975 3016 2984
rect 2964 2941 2973 2975
rect 2973 2941 3007 2975
rect 3007 2941 3016 2975
rect 2964 2932 3016 2941
rect 3148 2932 3200 2984
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 6736 3000 6788 3052
rect 5908 2932 5960 2984
rect 6920 2864 6972 2916
rect 7380 2864 7432 2916
rect 8116 3136 8168 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 10232 3136 10284 3188
rect 10876 3136 10928 3188
rect 8300 3068 8352 3120
rect 12532 3068 12584 3120
rect 15660 3136 15712 3188
rect 18052 3179 18104 3188
rect 18052 3145 18061 3179
rect 18061 3145 18095 3179
rect 18095 3145 18104 3179
rect 18052 3136 18104 3145
rect 19340 3068 19392 3120
rect 9772 3000 9824 3052
rect 8208 2932 8260 2984
rect 14280 3000 14332 3052
rect 14372 3043 14424 3052
rect 14372 3009 14381 3043
rect 14381 3009 14415 3043
rect 14415 3009 14424 3043
rect 16856 3043 16908 3052
rect 14372 3000 14424 3009
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 19064 3000 19116 3052
rect 12348 2932 12400 2984
rect 15568 2932 15620 2984
rect 16580 2932 16632 2984
rect 18144 2932 18196 2984
rect 20076 2932 20128 2984
rect 14740 2864 14792 2916
rect 17960 2864 18012 2916
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 10508 2796 10560 2848
rect 10600 2796 10652 2848
rect 13728 2796 13780 2848
rect 14556 2796 14608 2848
rect 18144 2796 18196 2848
rect 19616 2839 19668 2848
rect 19616 2805 19625 2839
rect 19625 2805 19659 2839
rect 19659 2805 19668 2839
rect 19616 2796 19668 2805
rect 19800 2796 19852 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 5356 2592 5408 2644
rect 7472 2592 7524 2644
rect 9680 2592 9732 2644
rect 10508 2592 10560 2644
rect 18788 2592 18840 2644
rect 4804 2456 4856 2508
rect 7012 2456 7064 2508
rect 9220 2456 9272 2508
rect 10416 2456 10468 2508
rect 5080 2388 5132 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 7748 2431 7800 2440
rect 5448 2388 5500 2397
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 12624 2499 12676 2508
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 10324 2388 10376 2397
rect 13820 2524 13872 2576
rect 13912 2499 13964 2508
rect 13912 2465 13921 2499
rect 13921 2465 13955 2499
rect 13955 2465 13964 2499
rect 13912 2456 13964 2465
rect 17868 2524 17920 2576
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 19616 2456 19668 2508
rect 5724 2320 5776 2372
rect 7196 2320 7248 2372
rect 8116 2320 8168 2372
rect 9772 2320 9824 2372
rect 10140 2320 10192 2372
rect 10876 2320 10928 2372
rect 11796 2320 11848 2372
rect 20996 2320 21048 2372
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 17684 2252 17736 2304
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3056 2048 3108 2100
rect 13176 2048 13228 2100
rect 5080 1980 5132 2032
rect 17960 1980 18012 2032
rect 10784 1912 10836 1964
rect 15936 1912 15988 1964
rect 9404 1300 9456 1352
rect 18144 1300 18196 1352
rect 10416 1232 10468 1284
rect 18052 1232 18104 1284
rect 9680 1164 9732 1216
rect 10968 1164 11020 1216
rect 17960 1164 18012 1216
<< metal2 >>
rect 294 22520 350 23000
rect 846 22520 902 23000
rect 1398 22520 1454 23000
rect 1950 22520 2006 23000
rect 2502 22520 2558 23000
rect 3054 22520 3110 23000
rect 3606 22520 3662 23000
rect 4158 22520 4214 23000
rect 4710 22520 4766 23000
rect 5262 22520 5318 23000
rect 5814 22520 5870 23000
rect 6458 22520 6514 23000
rect 7010 22520 7066 23000
rect 7562 22520 7618 23000
rect 8114 22520 8170 23000
rect 8666 22520 8722 23000
rect 9218 22520 9274 23000
rect 9770 22520 9826 23000
rect 10322 22520 10378 23000
rect 10782 22536 10838 22545
rect 308 11014 336 22520
rect 860 19242 888 22520
rect 1412 19666 1440 22520
rect 1964 20890 1992 22520
rect 2516 21162 2544 22520
rect 2516 21134 2728 21162
rect 1964 20862 2084 20890
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1964 20602 1992 20742
rect 1952 20596 2004 20602
rect 1952 20538 2004 20544
rect 1412 19638 1532 19666
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 848 19236 900 19242
rect 848 19178 900 19184
rect 1412 18222 1440 19450
rect 1504 18630 1532 19638
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1766 17096 1822 17105
rect 1766 17031 1822 17040
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 15570 1624 16934
rect 1780 16794 1808 17031
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 15706 1808 16390
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1582 15056 1638 15065
rect 1582 14991 1638 15000
rect 1398 13560 1454 13569
rect 1398 13495 1400 13504
rect 1452 13495 1454 13504
rect 1400 13466 1452 13472
rect 1596 12986 1624 14991
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 11665 1440 12718
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 296 11008 348 11014
rect 296 10950 348 10956
rect 1688 10033 1716 13806
rect 1780 13394 1808 14418
rect 2056 14278 2084 20862
rect 2228 20868 2280 20874
rect 2228 20810 2280 20816
rect 2240 20058 2268 20810
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2228 20052 2280 20058
rect 2228 19994 2280 20000
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1860 14000 1912 14006
rect 1858 13968 1860 13977
rect 1912 13968 1914 13977
rect 1858 13903 1914 13912
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1674 10024 1730 10033
rect 1674 9959 1730 9968
rect 2424 8498 2452 19246
rect 2516 19174 2544 20198
rect 2596 19304 2648 19310
rect 2596 19246 2648 19252
rect 2504 19168 2556 19174
rect 2504 19110 2556 19116
rect 2608 18986 2636 19246
rect 2516 18958 2636 18986
rect 2516 18222 2544 18958
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 2608 18222 2636 18770
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2596 18216 2648 18222
rect 2596 18158 2648 18164
rect 2516 17066 2544 18158
rect 2700 18034 2728 21134
rect 2872 20936 2924 20942
rect 2872 20878 2924 20884
rect 2884 20262 2912 20878
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2700 18006 2820 18034
rect 2792 17882 2820 18006
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2884 17762 2912 19178
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2792 17734 2912 17762
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 17134 2636 17614
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 2516 13462 2544 16594
rect 2594 16008 2650 16017
rect 2594 15943 2596 15952
rect 2648 15943 2650 15952
rect 2596 15914 2648 15920
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2516 6730 2544 13398
rect 2700 12714 2728 13806
rect 2792 13326 2820 17734
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2884 14385 2912 17002
rect 2976 16114 3004 18566
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2870 14376 2926 14385
rect 2870 14311 2926 14320
rect 2884 13870 2912 14311
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2688 12708 2740 12714
rect 2688 12650 2740 12656
rect 2884 8838 2912 13466
rect 2976 11762 3004 15370
rect 3068 13530 3096 22520
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 3160 20602 3188 20946
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12782 3096 13262
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 3054 12200 3110 12209
rect 3054 12135 3056 12144
rect 3108 12135 3110 12144
rect 3056 12106 3108 12112
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 848 4004 900 4010
rect 848 3946 900 3952
rect 296 3528 348 3534
rect 296 3470 348 3476
rect 308 480 336 3470
rect 860 480 888 3946
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1412 480 1440 3402
rect 1964 480 1992 6666
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4758 2176 4966
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2700 3602 2728 6598
rect 2884 5794 2912 8774
rect 3160 7546 3188 20334
rect 3252 18970 3280 20538
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3344 17762 3372 19314
rect 3516 18148 3568 18154
rect 3516 18090 3568 18096
rect 3252 17734 3372 17762
rect 3252 12714 3280 17734
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 17270 3372 17614
rect 3528 17610 3556 18090
rect 3516 17604 3568 17610
rect 3516 17546 3568 17552
rect 3528 17338 3556 17546
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3332 17264 3384 17270
rect 3332 17206 3384 17212
rect 3514 17232 3570 17241
rect 3514 17167 3570 17176
rect 3332 15632 3384 15638
rect 3332 15574 3384 15580
rect 3344 15473 3372 15574
rect 3330 15464 3386 15473
rect 3330 15399 3386 15408
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3436 14521 3464 14894
rect 3422 14512 3478 14521
rect 3422 14447 3478 14456
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3528 9722 3556 17167
rect 3620 16046 3648 22520
rect 4172 19394 4200 22520
rect 4724 20890 4752 22520
rect 4724 20862 4844 20890
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4816 20466 4844 20862
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4264 19530 4292 19790
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4264 19502 4384 19530
rect 4172 19366 4292 19394
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3804 18086 3832 18566
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 4080 17921 4108 18770
rect 4172 18086 4200 19178
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4066 17912 4122 17921
rect 4066 17847 4122 17856
rect 3700 17536 3752 17542
rect 3700 17478 3752 17484
rect 3712 16658 3740 17478
rect 3792 17332 3844 17338
rect 3792 17274 3844 17280
rect 3804 16726 3832 17274
rect 4172 17202 4200 18022
rect 4264 17864 4292 19366
rect 4356 19174 4384 19502
rect 4816 19446 4844 19926
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4344 19168 4396 19174
rect 4344 19110 4396 19116
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4344 17876 4396 17882
rect 4264 17836 4344 17864
rect 4344 17818 4396 17824
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 3792 16720 3844 16726
rect 3792 16662 3844 16668
rect 3700 16652 3752 16658
rect 3700 16594 3752 16600
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3700 14952 3752 14958
rect 3700 14894 3752 14900
rect 3712 14385 3740 14894
rect 3698 14376 3754 14385
rect 3698 14311 3754 14320
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3712 14074 3740 14214
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 10674 3648 12650
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3606 9616 3662 9625
rect 3606 9551 3662 9560
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3056 7268 3108 7274
rect 3056 7210 3108 7216
rect 3332 7268 3384 7274
rect 3332 7210 3384 7216
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2976 5914 3004 6054
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 3068 5817 3096 7210
rect 3054 5808 3110 5817
rect 2884 5766 3004 5794
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2044 3120 2096 3126
rect 2042 3088 2044 3097
rect 2096 3088 2098 3097
rect 2042 3023 2098 3032
rect 2792 2802 2820 4626
rect 2870 3496 2926 3505
rect 2870 3431 2926 3440
rect 2884 3398 2912 3431
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2976 2990 3004 5766
rect 3054 5743 3110 5752
rect 3344 5574 3372 7210
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3160 5234 3188 5510
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3160 4282 3188 5170
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3054 3768 3110 3777
rect 3054 3703 3110 3712
rect 3068 3398 3096 3703
rect 3056 3392 3108 3398
rect 3056 3334 3108 3340
rect 3160 2990 3188 4218
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3252 3738 3280 3946
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2516 2774 2820 2802
rect 2516 480 2544 2774
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 2106 3096 2246
rect 3056 2100 3108 2106
rect 3056 2042 3108 2048
rect 3344 1986 3372 5306
rect 3068 1958 3372 1986
rect 3068 480 3096 1958
rect 3620 480 3648 9551
rect 3712 6662 3740 14010
rect 3884 13796 3936 13802
rect 3884 13738 3936 13744
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 11694 3832 13670
rect 3896 12918 3924 13738
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3896 10606 3924 12650
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3988 6905 4016 15982
rect 4172 15570 4200 16934
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 14006 4108 14826
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4080 11762 4108 13942
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4172 11694 4200 12582
rect 4264 11898 4292 13330
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 4172 5370 4200 11494
rect 4264 11354 4292 11630
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4356 7750 4384 17818
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4816 16590 4844 17546
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17134 4936 17478
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4908 16522 4936 16934
rect 4896 16516 4948 16522
rect 4896 16458 4948 16464
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 5000 16250 5028 17614
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5092 15688 5120 20198
rect 5184 19990 5212 20402
rect 5276 20262 5304 22520
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5172 19984 5224 19990
rect 5172 19926 5224 19932
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5184 18426 5212 18838
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 18465 5304 18634
rect 5262 18456 5318 18465
rect 5172 18420 5224 18426
rect 5262 18391 5318 18400
rect 5172 18362 5224 18368
rect 5368 18358 5396 18702
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5184 16726 5212 18022
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 5172 16720 5224 16726
rect 5172 16662 5224 16668
rect 5276 16114 5304 17546
rect 5368 17524 5396 18022
rect 5460 17678 5488 20470
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18834 5580 19110
rect 5644 18902 5672 19654
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5538 18320 5594 18329
rect 5538 18255 5594 18264
rect 5552 18222 5580 18255
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5538 18048 5594 18057
rect 5538 17983 5594 17992
rect 5552 17814 5580 17983
rect 5644 17814 5672 18838
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5632 17808 5684 17814
rect 5632 17750 5684 17756
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5368 17496 5580 17524
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5000 15660 5120 15688
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4908 14618 4936 14758
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4804 14408 4856 14414
rect 4802 14376 4804 14385
rect 4856 14376 4858 14385
rect 4802 14311 4858 14320
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4540 12170 4568 12718
rect 4816 12442 4844 13738
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4712 12368 4764 12374
rect 5000 12322 5028 15660
rect 5276 15502 5304 16050
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5276 15162 5304 15438
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5276 14618 5304 15098
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5184 12850 5212 13126
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4712 12310 4764 12316
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4724 12084 4752 12310
rect 4908 12294 5028 12322
rect 4724 12056 4844 12084
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4434 11792 4490 11801
rect 4434 11727 4490 11736
rect 4448 11354 4476 11727
rect 4816 11558 4844 12056
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4908 11370 4936 12294
rect 5092 11898 5120 12582
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4436 11348 4488 11354
rect 4908 11342 5028 11370
rect 4436 11290 4488 11296
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4802 10976 4858 10985
rect 4421 10908 4717 10928
rect 4802 10911 4858 10920
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4618 10568 4674 10577
rect 4618 10503 4620 10512
rect 4672 10503 4674 10512
rect 4620 10474 4672 10480
rect 4816 10266 4844 10911
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4802 9480 4858 9489
rect 4802 9415 4804 9424
rect 4856 9415 4858 9424
rect 4804 9386 4856 9392
rect 4908 9178 4936 11018
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4434 8392 4490 8401
rect 4434 8327 4490 8336
rect 4448 8090 4476 8327
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5778 4384 6258
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5370 4384 5714
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4172 4622 4200 5034
rect 4816 4826 4844 6054
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4172 4282 4200 4558
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4264 3466 4292 4626
rect 4908 4554 4936 5238
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 5000 4486 5028 11342
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4436 3528 4488 3534
rect 4356 3476 4436 3482
rect 4356 3470 4488 3476
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4356 3454 4476 3470
rect 4356 3210 4384 3454
rect 4802 3360 4858 3369
rect 4421 3292 4717 3312
rect 4802 3295 4858 3304
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4080 3182 4384 3210
rect 4080 2990 4108 3182
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4816 2666 4844 3295
rect 4172 2638 4844 2666
rect 4172 480 4200 2638
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1306 4844 2450
rect 5092 2446 5120 11494
rect 5184 11218 5212 12038
rect 5276 11234 5304 13262
rect 5368 11370 5396 15506
rect 5460 15434 5488 17002
rect 5552 15722 5580 17496
rect 5632 16584 5684 16590
rect 5632 16526 5684 16532
rect 5644 15892 5672 16526
rect 5736 16046 5764 20334
rect 5828 19394 5856 22520
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 5828 19366 6040 19394
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 18970 5856 19110
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5816 18284 5868 18290
rect 5816 18226 5868 18232
rect 5828 17202 5856 18226
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5828 16114 5856 17138
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5644 15864 5764 15892
rect 5552 15694 5672 15722
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5552 13734 5580 15574
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12764 5488 13126
rect 5552 12918 5580 13330
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5460 12736 5580 12764
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5460 12306 5488 12378
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5552 12170 5580 12736
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 5552 11762 5580 12106
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5644 11558 5672 15694
rect 5736 15162 5764 15864
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5736 14385 5764 15098
rect 5814 14920 5870 14929
rect 5814 14855 5870 14864
rect 5722 14376 5778 14385
rect 5722 14311 5778 14320
rect 5736 12918 5764 14311
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12306 5764 12854
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5368 11342 5488 11370
rect 5172 11212 5224 11218
rect 5276 11206 5396 11234
rect 5172 11154 5224 11160
rect 5264 11144 5316 11150
rect 5264 11086 5316 11092
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 6458 5212 7278
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5170 4040 5226 4049
rect 5170 3975 5226 3984
rect 5184 3942 5212 3975
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5092 2038 5120 2382
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 4724 1278 4844 1306
rect 4724 480 4752 1278
rect 5276 480 5304 11086
rect 5368 9994 5396 11206
rect 5460 11121 5488 11342
rect 5828 11150 5856 14855
rect 5816 11144 5868 11150
rect 5446 11112 5502 11121
rect 5816 11086 5868 11092
rect 5446 11047 5502 11056
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5460 9874 5488 11047
rect 5816 10736 5868 10742
rect 5814 10704 5816 10713
rect 5868 10704 5870 10713
rect 5814 10639 5870 10648
rect 5368 9846 5488 9874
rect 5368 5302 5396 9846
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5460 7342 5488 7482
rect 5644 7478 5672 8298
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5460 5642 5488 5782
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5356 5296 5408 5302
rect 5356 5238 5408 5244
rect 5460 4622 5488 5578
rect 5736 4826 5764 6734
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 2650 5396 3878
rect 5552 3738 5580 4626
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3194 5488 3538
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5460 2446 5488 3130
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5736 2378 5764 3946
rect 5828 3738 5856 4014
rect 5920 3942 5948 19246
rect 6012 18902 6040 19366
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 6000 18216 6052 18222
rect 6000 18158 6052 18164
rect 6012 18057 6040 18158
rect 5998 18048 6054 18057
rect 5998 17983 6054 17992
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6012 9586 6040 16186
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 6104 4049 6132 19246
rect 6196 17882 6224 20334
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6288 17338 6316 17818
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6276 16992 6328 16998
rect 6276 16934 6328 16940
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6196 15638 6224 16050
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6196 14278 6224 15574
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6196 13938 6224 14214
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 6182 12336 6238 12345
rect 6182 12271 6238 12280
rect 6196 11354 6224 12271
rect 6288 11354 6316 16934
rect 6380 16250 6408 20198
rect 6472 19174 6500 22520
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6644 19916 6696 19922
rect 6644 19858 6696 19864
rect 6656 19242 6684 19858
rect 6644 19236 6696 19242
rect 6644 19178 6696 19184
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6656 18766 6684 18838
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6748 18426 6776 20266
rect 6840 19922 6868 20402
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6840 18698 6868 19858
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6644 18420 6696 18426
rect 6644 18362 6696 18368
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6472 17338 6500 17682
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6368 16040 6420 16046
rect 6368 15982 6420 15988
rect 6380 15178 6408 15982
rect 6472 15910 6500 16186
rect 6460 15904 6512 15910
rect 6460 15846 6512 15852
rect 6380 15162 6500 15178
rect 6380 15156 6512 15162
rect 6380 15150 6460 15156
rect 6380 12889 6408 15150
rect 6460 15098 6512 15104
rect 6564 14822 6592 17682
rect 6656 17270 6684 18362
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6748 17814 6776 18226
rect 6826 18184 6882 18193
rect 6826 18119 6882 18128
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6840 16810 6868 18119
rect 6748 16782 6868 16810
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6552 14816 6604 14822
rect 6748 14770 6776 16782
rect 6828 16720 6880 16726
rect 6932 16708 6960 20470
rect 7024 18902 7052 22520
rect 7576 20534 7604 22520
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 8128 20346 8156 22520
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8128 20318 8248 20346
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19378 7512 19858
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 8036 19446 8064 19722
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 8024 19440 8076 19446
rect 8024 19382 8076 19388
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7012 18896 7064 18902
rect 7012 18838 7064 18844
rect 7012 18760 7064 18766
rect 7064 18708 7236 18714
rect 7012 18702 7236 18708
rect 7024 18698 7236 18702
rect 7024 18692 7248 18698
rect 7024 18686 7196 18692
rect 7196 18634 7248 18640
rect 7288 18216 7340 18222
rect 7024 18176 7288 18204
rect 7024 18086 7052 18176
rect 7288 18158 7340 18164
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7010 17912 7066 17921
rect 7010 17847 7066 17856
rect 7024 17814 7052 17847
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 7116 17134 7144 18022
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 7024 16726 7052 16934
rect 6880 16680 6960 16708
rect 7012 16720 7064 16726
rect 6828 16662 6880 16668
rect 7012 16662 7064 16668
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15706 6868 15846
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6552 14758 6604 14764
rect 6472 14550 6500 14758
rect 6656 14742 6776 14770
rect 6460 14544 6512 14550
rect 6460 14486 6512 14492
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6366 12880 6422 12889
rect 6366 12815 6422 12824
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6380 11082 6408 12718
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6288 5710 6316 6258
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6288 5574 6316 5646
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5234 6316 5510
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6368 4752 6420 4758
rect 6368 4694 6420 4700
rect 6380 4282 6408 4694
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5828 480 5856 3470
rect 5920 2990 5948 3674
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6472 480 6500 13398
rect 6564 4758 6592 13670
rect 6656 11626 6684 14742
rect 6840 13954 6868 15302
rect 6932 14958 6960 15982
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14056 6960 14894
rect 7024 14226 7052 16186
rect 7116 16153 7144 17070
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7102 16144 7158 16153
rect 7102 16079 7158 16088
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15700 7156 15706
rect 7104 15642 7156 15648
rect 7116 14618 7144 15642
rect 7208 15026 7236 15846
rect 7300 15706 7328 16594
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15162 7328 15302
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7024 14198 7144 14226
rect 6932 14028 7052 14056
rect 6840 13926 6960 13954
rect 6932 13870 6960 13926
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6840 12986 6868 13806
rect 7024 13258 7052 14028
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7116 12986 7144 14198
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 7102 12880 7158 12889
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6748 10606 6776 12854
rect 7102 12815 7158 12824
rect 7116 12646 7144 12815
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6840 11762 6868 12242
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 7208 11286 7236 14826
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 14006 7328 14418
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7300 12646 7328 12922
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7392 12458 7420 17614
rect 7484 13569 7512 17682
rect 7576 15881 7604 19382
rect 8128 19310 8156 19654
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 8220 18426 8248 20318
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19310 8432 19654
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 7562 15872 7618 15881
rect 7562 15807 7618 15816
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7576 14362 7604 15642
rect 7668 14550 7696 17478
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7760 16454 7788 17138
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8220 16658 8248 17478
rect 8312 17202 8340 19178
rect 8496 18154 8524 20402
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7852 15960 7880 16594
rect 7760 15932 7880 15960
rect 7760 14890 7788 15932
rect 8312 15910 8340 17138
rect 8484 17128 8536 17134
rect 8484 17070 8536 17076
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8208 15564 8260 15570
rect 8312 15552 8340 15846
rect 8260 15524 8340 15552
rect 8208 15506 8260 15512
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7656 14544 7708 14550
rect 7840 14544 7892 14550
rect 7656 14486 7708 14492
rect 7746 14512 7802 14521
rect 7840 14486 7892 14492
rect 7746 14447 7802 14456
rect 7760 14414 7788 14447
rect 7656 14408 7708 14414
rect 7576 14356 7656 14362
rect 7576 14350 7708 14356
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7576 14334 7696 14350
rect 7852 13802 7880 14486
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7470 13560 7526 13569
rect 7886 13552 8182 13572
rect 7470 13495 7526 13504
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12850 7512 13262
rect 7562 13016 7618 13025
rect 7562 12951 7618 12960
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7300 12430 7420 12458
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 11014 6960 11086
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6840 10169 6868 10202
rect 7116 10198 7144 10474
rect 7208 10470 7236 10746
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7104 10192 7156 10198
rect 6826 10160 6882 10169
rect 7104 10134 7156 10140
rect 6826 10095 6882 10104
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9761 7144 9862
rect 7102 9752 7158 9761
rect 7102 9687 7158 9696
rect 7208 9602 7236 10406
rect 7300 9625 7328 12430
rect 7199 9574 7236 9602
rect 7286 9616 7342 9625
rect 6644 9512 6696 9518
rect 7199 9500 7227 9574
rect 7286 9551 7342 9560
rect 7199 9472 7236 9500
rect 6644 9454 6696 9460
rect 6656 9042 6684 9454
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6656 8022 6684 8978
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 8090 6960 8230
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6656 7546 6684 7958
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6656 6322 6684 7482
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6840 7002 6868 7278
rect 6932 7206 6960 7890
rect 7024 7410 7052 8434
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6866 6960 7142
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6642 4040 6698 4049
rect 6642 3975 6698 3984
rect 6656 3942 6684 3975
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6748 3602 6776 5170
rect 6918 5128 6974 5137
rect 6918 5063 6974 5072
rect 6932 4554 6960 5063
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6826 4176 6882 4185
rect 6826 4111 6882 4120
rect 6840 3602 6868 4111
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6748 3058 6776 3538
rect 6918 3224 6974 3233
rect 6918 3159 6974 3168
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6932 2922 6960 3159
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7024 480 7052 2450
rect 7208 2378 7236 9472
rect 7484 7426 7512 12582
rect 7576 10130 7604 12951
rect 7760 12850 7788 13330
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 7748 12844 7800 12850
rect 8220 12832 8248 13942
rect 8298 13696 8354 13705
rect 8298 13631 8354 13640
rect 8312 13530 8340 13631
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 7748 12786 7800 12792
rect 8128 12804 8248 12832
rect 7760 12442 7788 12786
rect 8128 12714 8156 12804
rect 8116 12708 8168 12714
rect 8116 12650 8168 12656
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7748 12436 7800 12442
rect 7748 12378 7800 12384
rect 7668 12152 7696 12378
rect 8220 12306 8248 12650
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7748 12164 7800 12170
rect 7668 12124 7748 12152
rect 7748 12106 7800 12112
rect 8220 11898 8248 12242
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8404 11830 8432 16594
rect 8496 14618 8524 17070
rect 8588 15638 8616 20334
rect 8680 19394 8708 22520
rect 8680 19366 8984 19394
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8680 18834 8708 19246
rect 8956 18834 8984 19366
rect 9232 19310 9260 22520
rect 9784 20482 9812 22520
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 9784 20454 10088 20482
rect 9864 20324 9916 20330
rect 9864 20266 9916 20272
rect 9876 20233 9904 20266
rect 9862 20224 9918 20233
rect 9862 20159 9918 20168
rect 9678 20088 9734 20097
rect 9678 20023 9680 20032
rect 9732 20023 9734 20032
rect 9680 19994 9732 20000
rect 9772 19984 9824 19990
rect 9770 19952 9772 19961
rect 9956 19984 10008 19990
rect 9824 19952 9826 19961
rect 9956 19926 10008 19932
rect 9770 19887 9826 19896
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9692 19378 9720 19790
rect 9770 19680 9826 19689
rect 9770 19615 9826 19624
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9312 19168 9364 19174
rect 9310 19136 9312 19145
rect 9496 19168 9548 19174
rect 9364 19136 9366 19145
rect 9496 19110 9548 19116
rect 9310 19071 9366 19080
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8760 18692 8812 18698
rect 8760 18634 8812 18640
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8680 16114 8708 18022
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8576 15632 8628 15638
rect 8576 15574 8628 15580
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8680 15473 8708 15574
rect 8666 15464 8722 15473
rect 8666 15399 8722 15408
rect 8772 15314 8800 18634
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9140 18290 9168 18566
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8864 17066 8892 18158
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9140 17105 9168 18022
rect 9126 17096 9182 17105
rect 8852 17060 8904 17066
rect 9126 17031 9182 17040
rect 8852 17002 8904 17008
rect 8864 16590 8892 17002
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8850 16144 8906 16153
rect 8850 16079 8906 16088
rect 8588 15286 8800 15314
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8482 14376 8538 14385
rect 8482 14311 8538 14320
rect 8496 13530 8524 14311
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8482 12064 8538 12073
rect 8482 11999 8538 12008
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8220 11558 8248 11698
rect 8496 11626 8524 11999
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8390 11520 8446 11529
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 7930 11248 7986 11257
rect 7930 11183 7986 11192
rect 7944 11082 7972 11183
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 8220 11014 8248 11086
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 8220 10266 8248 10542
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7392 7398 7512 7426
rect 7392 5137 7420 7398
rect 7576 6934 7604 10066
rect 8206 9616 8262 9625
rect 8206 9551 8262 9560
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7760 9178 7788 9386
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8220 9178 8248 9551
rect 8312 9518 8340 11494
rect 8390 11455 8446 11464
rect 8404 11354 8432 11455
rect 8496 11354 8524 11562
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8588 11286 8616 15286
rect 8864 14929 8892 16079
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9232 14958 9260 15846
rect 9324 15065 9352 18566
rect 9508 18290 9536 19110
rect 9692 18766 9720 19314
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9586 18456 9642 18465
rect 9586 18391 9642 18400
rect 9600 18290 9628 18391
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9692 16046 9720 16390
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9310 15056 9366 15065
rect 9310 14991 9366 15000
rect 9220 14952 9272 14958
rect 8850 14920 8906 14929
rect 9220 14894 9272 14900
rect 9312 14952 9364 14958
rect 9364 14912 9536 14940
rect 9312 14894 9364 14900
rect 9508 14906 9536 14912
rect 8850 14855 8906 14864
rect 8852 14816 8904 14822
rect 8758 14784 8814 14793
rect 8852 14758 8904 14764
rect 8758 14719 8814 14728
rect 8772 13977 8800 14719
rect 8758 13968 8814 13977
rect 8758 13903 8814 13912
rect 8864 13802 8892 14758
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8942 13832 8998 13841
rect 8852 13796 8904 13802
rect 8942 13767 8998 13776
rect 8852 13738 8904 13744
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12617 8708 13262
rect 8772 13161 8800 13670
rect 8758 13152 8814 13161
rect 8758 13087 8814 13096
rect 8760 12640 8812 12646
rect 8666 12608 8722 12617
rect 8760 12582 8812 12588
rect 8666 12543 8722 12552
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8680 12102 8708 12242
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8772 11898 8800 12582
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8772 11558 8800 11630
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 8758 11248 8814 11257
rect 8392 11212 8444 11218
rect 8758 11183 8814 11192
rect 8392 11154 8444 11160
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8300 9376 8352 9382
rect 8298 9344 8300 9353
rect 8352 9344 8354 9353
rect 8298 9279 8354 9288
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7668 8430 7696 8978
rect 7760 8498 7788 9114
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 7954 7696 8366
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8220 8022 8248 8298
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 7656 7948 7708 7954
rect 7656 7890 7708 7896
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7002 7788 7822
rect 8312 7818 8340 8230
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 5692 7604 6870
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6186 7696 6734
rect 7656 6180 7708 6186
rect 7656 6122 7708 6128
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7668 5914 7696 6122
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7576 5664 7696 5692
rect 7472 5160 7524 5166
rect 7378 5128 7434 5137
rect 7472 5102 7524 5108
rect 7378 5063 7434 5072
rect 7484 4622 7512 5102
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7378 2952 7434 2961
rect 7378 2887 7380 2896
rect 7432 2887 7434 2896
rect 7380 2858 7432 2864
rect 7484 2650 7512 4014
rect 7576 3233 7604 4082
rect 7562 3224 7618 3233
rect 7562 3159 7618 3168
rect 7668 3108 7696 5664
rect 7760 4758 7788 6054
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8220 5166 8248 6054
rect 8312 5778 8340 6122
rect 8404 6118 8432 11154
rect 8576 11144 8628 11150
rect 8628 11104 8708 11132
rect 8576 11086 8628 11092
rect 8482 10840 8538 10849
rect 8482 10775 8538 10784
rect 8496 10266 8524 10775
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8484 10056 8536 10062
rect 8588 10044 8616 10202
rect 8536 10016 8616 10044
rect 8484 9998 8536 10004
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8496 8090 8524 9590
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8588 7954 8616 8774
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8496 7342 8524 7822
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8588 7274 8616 7890
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8680 7206 8708 11104
rect 8772 9654 8800 11183
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8864 9382 8892 13738
rect 8956 12306 8984 13767
rect 9048 13569 9076 13874
rect 9034 13560 9090 13569
rect 9034 13495 9090 13504
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9048 12102 9076 13330
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12481 9168 13194
rect 9126 12472 9182 12481
rect 9126 12407 9182 12416
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 7268 8812 7274
rect 8760 7210 8812 7216
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8482 6896 8538 6905
rect 8482 6831 8538 6840
rect 8496 6798 8524 6831
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8496 5778 8524 6734
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8772 5370 8800 7210
rect 8956 6458 8984 11222
rect 9048 9042 9076 12038
rect 9140 11393 9168 12242
rect 9126 11384 9182 11393
rect 9126 11319 9182 11328
rect 9232 10674 9260 14894
rect 9508 14890 9628 14906
rect 9508 14884 9640 14890
rect 9508 14878 9588 14884
rect 9588 14826 9640 14832
rect 9680 14272 9732 14278
rect 9678 14240 9680 14249
rect 9732 14240 9734 14249
rect 9678 14175 9734 14184
rect 9588 13796 9640 13802
rect 9416 13756 9588 13784
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9324 12850 9352 13670
rect 9416 13569 9444 13756
rect 9588 13738 9640 13744
rect 9784 13569 9812 19615
rect 9968 19514 9996 19926
rect 9956 19508 10008 19514
rect 9956 19450 10008 19456
rect 10060 18873 10088 20454
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10152 20097 10180 20266
rect 10138 20088 10194 20097
rect 10138 20023 10194 20032
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10046 18864 10102 18873
rect 10046 18799 10102 18808
rect 10152 17864 10180 19450
rect 10060 17836 10180 17864
rect 10060 17338 10088 17836
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9876 14414 9904 16390
rect 10060 16130 10088 17274
rect 9968 16114 10088 16130
rect 9956 16108 10088 16114
rect 10008 16102 10088 16108
rect 9956 16050 10008 16056
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 14550 9996 15846
rect 10046 14648 10102 14657
rect 10046 14583 10102 14592
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9864 14408 9916 14414
rect 9916 14368 9996 14396
rect 9864 14350 9916 14356
rect 9968 14113 9996 14368
rect 9954 14104 10010 14113
rect 9864 14068 9916 14074
rect 9954 14039 10010 14048
rect 9864 14010 9916 14016
rect 9402 13560 9458 13569
rect 9402 13495 9458 13504
rect 9770 13560 9826 13569
rect 9770 13495 9826 13504
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9416 12050 9444 13398
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9324 12022 9444 12050
rect 9324 11694 9352 12022
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9416 11529 9444 11834
rect 9508 11762 9536 12650
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9402 11520 9458 11529
rect 9402 11455 9458 11464
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9416 10810 9444 11290
rect 9600 11218 9628 13330
rect 9876 13326 9904 14010
rect 9954 13696 10010 13705
rect 9954 13631 10010 13640
rect 9968 13530 9996 13631
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9954 13288 10010 13297
rect 9692 12073 9720 13262
rect 9954 13223 10010 13232
rect 9862 13016 9918 13025
rect 9862 12951 9918 12960
rect 9770 12880 9826 12889
rect 9770 12815 9826 12824
rect 9678 12064 9734 12073
rect 9678 11999 9734 12008
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9692 10588 9720 11154
rect 9324 10560 9720 10588
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10062 9168 10406
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9518 9168 9998
rect 9128 9512 9180 9518
rect 9220 9512 9272 9518
rect 9128 9454 9180 9460
rect 9218 9480 9220 9489
rect 9272 9480 9274 9489
rect 9140 9042 9168 9454
rect 9218 9415 9274 9424
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9140 8090 9168 8978
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7760 3777 7788 3878
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7746 3768 7802 3777
rect 7886 3760 8182 3780
rect 7746 3703 7802 3712
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7576 3080 7696 3108
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7576 480 7604 3080
rect 7760 2961 7788 3334
rect 8114 3224 8170 3233
rect 8114 3159 8116 3168
rect 8168 3159 8170 3168
rect 8116 3130 8168 3136
rect 8220 2990 8248 4966
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 4146 8524 4422
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 3369 8340 3470
rect 8298 3360 8354 3369
rect 8298 3295 8354 3304
rect 8300 3120 8352 3126
rect 8298 3088 8300 3097
rect 8352 3088 8354 3097
rect 8298 3023 8354 3032
rect 8208 2984 8260 2990
rect 7746 2952 7802 2961
rect 8208 2926 8260 2932
rect 7746 2887 7802 2896
rect 7760 2446 7788 2887
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8128 480 8156 2314
rect 8680 480 8708 5170
rect 8772 4622 8800 5306
rect 9048 5234 9076 8026
rect 9140 7886 9168 8026
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 6322 9168 7822
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5778 9168 6258
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 5914 9260 6190
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4826 9076 5034
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 9324 3534 9352 10560
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9692 9994 9720 10406
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9496 9376 9548 9382
rect 9600 9353 9628 9386
rect 9496 9318 9548 9324
rect 9586 9344 9642 9353
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 5166 9444 7686
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9508 5012 9536 9318
rect 9586 9279 9642 9288
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9416 4984 9536 5012
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9232 480 9260 2450
rect 9416 1358 9444 4984
rect 9692 4622 9720 5714
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4298 9720 4558
rect 9784 4554 9812 12815
rect 9876 12306 9904 12951
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 10282 9904 12106
rect 9968 10470 9996 13223
rect 10060 12170 10088 14583
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 10060 11694 10088 11766
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10046 11520 10102 11529
rect 10046 11455 10102 11464
rect 10060 11354 10088 11455
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 10046 10296 10102 10305
rect 9876 10254 9996 10282
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9876 8430 9904 8774
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9772 4548 9824 4554
rect 9772 4490 9824 4496
rect 9876 4486 9904 8026
rect 9864 4480 9916 4486
rect 9864 4422 9916 4428
rect 9968 4298 9996 10254
rect 10046 10231 10048 10240
rect 10100 10231 10102 10240
rect 10048 10202 10100 10208
rect 10152 9058 10180 17682
rect 10244 14521 10272 21082
rect 10336 20505 10364 22520
rect 10874 22522 10930 23000
rect 10838 22520 10930 22522
rect 11426 22520 11482 23000
rect 12070 22520 12126 23000
rect 12622 22520 12678 23000
rect 13174 22520 13230 23000
rect 13726 22520 13782 23000
rect 14278 22520 14334 23000
rect 14830 22520 14886 23000
rect 15382 22520 15438 23000
rect 15934 22520 15990 23000
rect 16486 22520 16542 23000
rect 17038 22520 17094 23000
rect 17682 22520 17738 23000
rect 18234 22520 18290 23000
rect 18326 22672 18382 22681
rect 18326 22607 18382 22616
rect 10838 22494 10916 22520
rect 10782 22471 10838 22480
rect 11440 20890 11468 22520
rect 11440 20862 11744 20890
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11060 20528 11112 20534
rect 10322 20496 10378 20505
rect 11060 20470 11112 20476
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 10322 20431 10378 20440
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10336 19689 10364 20334
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10322 19680 10378 19689
rect 10322 19615 10378 19624
rect 10612 19514 10640 20198
rect 11072 19854 11100 20470
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10980 19378 11008 19654
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10336 18737 10364 19110
rect 10428 18902 10456 19314
rect 10506 19272 10562 19281
rect 10506 19207 10562 19216
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10322 18728 10378 18737
rect 10322 18663 10378 18672
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10230 14512 10286 14521
rect 10230 14447 10286 14456
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 14278 10272 14350
rect 10336 14278 10364 14418
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10060 9030 10180 9058
rect 10060 8090 10088 9030
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 10060 7478 10088 7890
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 10152 4808 10180 8910
rect 9508 4270 9720 4298
rect 9876 4270 9996 4298
rect 10060 4780 10180 4808
rect 9508 4010 9536 4270
rect 9600 4134 9812 4162
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9508 3534 9536 3946
rect 9600 3738 9628 4134
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9692 3194 9720 4014
rect 9784 3913 9812 4134
rect 9770 3904 9826 3913
rect 9770 3839 9826 3848
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9784 3602 9812 3674
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9784 3058 9812 3538
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9692 1222 9720 2586
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 9784 480 9812 2314
rect 9876 2258 9904 4270
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3602 9996 3878
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10060 2854 10088 4780
rect 10244 3942 10272 14214
rect 10428 13870 10456 16934
rect 10520 15910 10548 19207
rect 10876 19168 10928 19174
rect 10874 19136 10876 19145
rect 10928 19136 10930 19145
rect 10874 19071 10930 19080
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 10704 17338 10732 18362
rect 10888 18154 10916 19071
rect 10980 18902 11008 19314
rect 10968 18896 11020 18902
rect 10968 18838 11020 18844
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11072 18290 11100 18838
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11164 18222 11192 20470
rect 11716 20058 11744 20862
rect 11796 20324 11848 20330
rect 11796 20266 11848 20272
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11702 18728 11758 18737
rect 11256 18698 11376 18714
rect 11256 18692 11388 18698
rect 11256 18686 11336 18692
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10782 18048 10838 18057
rect 10782 17983 10838 17992
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10612 15706 10640 15846
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10520 14618 10548 15506
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 15094 10640 15438
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10506 14512 10562 14521
rect 10506 14447 10562 14456
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10520 13734 10548 14447
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10322 13560 10378 13569
rect 10322 13495 10324 13504
rect 10376 13495 10378 13504
rect 10324 13466 10376 13472
rect 10336 13161 10364 13466
rect 10322 13152 10378 13161
rect 10322 13087 10378 13096
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10336 11898 10364 12582
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10414 12064 10470 12073
rect 10414 11999 10470 12008
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10428 11778 10456 11999
rect 10336 11762 10456 11778
rect 10324 11756 10456 11762
rect 10376 11750 10456 11756
rect 10324 11698 10376 11704
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10849 10364 10950
rect 10322 10840 10378 10849
rect 10322 10775 10378 10784
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10266 10364 10406
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10336 4185 10364 8366
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10244 2394 10272 3130
rect 10336 2446 10364 3538
rect 10428 2514 10456 11630
rect 10520 11218 10548 12378
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10520 6322 10548 6666
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10612 4214 10640 15030
rect 10796 14958 10824 17983
rect 11058 17776 11114 17785
rect 11256 17746 11284 18686
rect 11702 18663 11758 18672
rect 11336 18634 11388 18640
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11058 17711 11114 17720
rect 11244 17740 11296 17746
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10980 16697 11008 17614
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 11072 16232 11100 17711
rect 11244 17682 11296 17688
rect 11256 17270 11284 17682
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 16794 11284 16934
rect 11716 16794 11744 18663
rect 11808 18222 11836 20266
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 18408 11928 19790
rect 12084 18986 12112 22520
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 11992 18958 12112 18986
rect 11992 18902 12020 18958
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 11900 18380 12020 18408
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11702 16688 11758 16697
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11244 16652 11296 16658
rect 11702 16623 11704 16632
rect 11244 16594 11296 16600
rect 11756 16623 11758 16632
rect 11704 16594 11756 16600
rect 10980 16204 11100 16232
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10704 13394 10732 13874
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10704 11898 10732 12174
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10704 11121 10732 11562
rect 10690 11112 10746 11121
rect 10690 11047 10746 11056
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10704 10441 10732 10678
rect 10690 10432 10746 10441
rect 10690 10367 10746 10376
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 8906 10732 9386
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10796 8294 10824 14894
rect 10888 14822 10916 16050
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 14482 10916 14758
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10980 14346 11008 16204
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11060 14340 11112 14346
rect 11060 14282 11112 14288
rect 10966 14104 11022 14113
rect 10966 14039 11022 14048
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 11286 10916 13670
rect 10980 11676 11008 14039
rect 11072 12764 11100 14282
rect 11164 12918 11192 16594
rect 11256 16454 11284 16594
rect 11244 16448 11296 16454
rect 11716 16436 11744 16594
rect 11808 16590 11836 17206
rect 11900 16794 11928 18226
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11716 16408 11836 16436
rect 11244 16390 11296 16396
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11440 15910 11468 16050
rect 11704 15972 11756 15978
rect 11704 15914 11756 15920
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 11256 15162 11284 15846
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11716 15065 11744 15914
rect 11808 15502 11836 16408
rect 11900 15570 11928 16730
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11702 15056 11758 15065
rect 11702 14991 11758 15000
rect 11808 14822 11836 15438
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11702 14376 11758 14385
rect 11702 14311 11758 14320
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11716 13870 11744 14311
rect 11244 13864 11296 13870
rect 11704 13864 11756 13870
rect 11244 13806 11296 13812
rect 11334 13832 11390 13841
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11072 12736 11192 12764
rect 11060 11688 11112 11694
rect 10980 11648 11060 11676
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10980 11132 11008 11648
rect 11060 11630 11112 11636
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10888 11104 11008 11132
rect 10888 9602 10916 11104
rect 11072 10538 11100 11154
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9722 11008 9998
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10888 9574 11008 9602
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10704 7546 10732 8230
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10888 6254 10916 6802
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10704 4128 10732 4966
rect 10796 4729 10824 5102
rect 10782 4720 10838 4729
rect 10782 4655 10838 4664
rect 10704 4100 10824 4128
rect 10690 4040 10746 4049
rect 10600 4004 10652 4010
rect 10690 3975 10692 3984
rect 10600 3946 10652 3952
rect 10744 3975 10746 3984
rect 10692 3946 10744 3952
rect 10612 2854 10640 3946
rect 10508 2848 10560 2854
rect 10508 2790 10560 2796
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10520 2650 10548 2790
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10152 2378 10272 2394
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10140 2372 10272 2378
rect 10192 2366 10272 2372
rect 10140 2314 10192 2320
rect 9876 2230 10364 2258
rect 10336 480 10364 2230
rect 10428 1290 10456 2450
rect 10796 1970 10824 4100
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3194 10916 4014
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10888 480 10916 2314
rect 10980 1222 11008 9574
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 7410 11100 7754
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 6934 11100 7346
rect 11164 6934 11192 12736
rect 11256 11354 11284 13806
rect 11704 13806 11756 13812
rect 11334 13767 11390 13776
rect 11348 13734 11376 13767
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11704 12912 11756 12918
rect 11702 12880 11704 12889
rect 11756 12880 11758 12889
rect 11702 12815 11758 12824
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11716 11880 11744 12815
rect 11808 12646 11836 13330
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11794 12064 11850 12073
rect 11794 11999 11850 12008
rect 11624 11852 11744 11880
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11624 11286 11652 11852
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11336 10532 11388 10538
rect 11336 10474 11388 10480
rect 11348 9994 11376 10474
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11256 7750 11284 8978
rect 11716 8974 11744 11698
rect 11808 10305 11836 11999
rect 11900 11558 11928 14418
rect 11992 14346 12020 18380
rect 12084 14550 12112 18838
rect 12164 18080 12216 18086
rect 12162 18048 12164 18057
rect 12216 18048 12218 18057
rect 12162 17983 12218 17992
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11980 14340 12032 14346
rect 11980 14282 12032 14288
rect 12084 14074 12112 14350
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12070 13832 12126 13841
rect 12070 13767 12126 13776
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12617 12020 13330
rect 11978 12608 12034 12617
rect 11978 12543 12034 12552
rect 11992 12170 12020 12543
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 11888 11552 11940 11558
rect 11992 11529 12020 11863
rect 11888 11494 11940 11500
rect 11978 11520 12034 11529
rect 11978 11455 12034 11464
rect 11978 11384 12034 11393
rect 11978 11319 11980 11328
rect 12032 11319 12034 11328
rect 11980 11290 12032 11296
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11794 10296 11850 10305
rect 11794 10231 11850 10240
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 7410 11744 7686
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 7002 11284 7142
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 11164 6662 11192 6734
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11072 5234 11100 5510
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11072 4758 11100 5170
rect 11164 5166 11192 5510
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 3670 11192 4422
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11256 1986 11284 3878
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11808 2378 11836 10231
rect 11900 8430 11928 11222
rect 11978 9616 12034 9625
rect 11978 9551 11980 9560
rect 12032 9551 12034 9560
rect 11980 9522 12032 9528
rect 12084 9466 12112 13767
rect 12176 13433 12204 14282
rect 12162 13424 12218 13433
rect 12162 13359 12218 13368
rect 12162 13288 12218 13297
rect 12162 13223 12218 13232
rect 12176 13190 12204 13223
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12176 12374 12204 12854
rect 12164 12368 12216 12374
rect 12164 12310 12216 12316
rect 12268 12322 12296 20198
rect 12636 19310 12664 22520
rect 13188 20074 13216 22520
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 12728 20046 13216 20074
rect 13280 20058 13308 20198
rect 13268 20052 13320 20058
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12348 18828 12400 18834
rect 12348 18770 12400 18776
rect 12624 18828 12676 18834
rect 12624 18770 12676 18776
rect 12360 16153 12388 18770
rect 12532 18760 12584 18766
rect 12530 18728 12532 18737
rect 12584 18728 12586 18737
rect 12530 18663 12586 18672
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12346 16144 12402 16153
rect 12346 16079 12402 16088
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12360 14822 12388 14894
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12360 13326 12388 14758
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12918 12388 13262
rect 12452 12986 12480 18158
rect 12532 18080 12584 18086
rect 12530 18048 12532 18057
rect 12584 18048 12586 18057
rect 12530 17983 12586 17992
rect 12636 17882 12664 18770
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12636 17202 12664 17818
rect 12624 17196 12676 17202
rect 12624 17138 12676 17144
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 15162 12664 15846
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 13530 12664 14758
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12624 13184 12676 13190
rect 12624 13126 12676 13132
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12912 12400 12918
rect 12636 12866 12664 13126
rect 12348 12854 12400 12860
rect 12544 12838 12664 12866
rect 12438 12744 12494 12753
rect 12438 12679 12494 12688
rect 12268 12294 12388 12322
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 10742 12204 12174
rect 12164 10736 12216 10742
rect 12164 10678 12216 10684
rect 12164 9920 12216 9926
rect 12162 9888 12164 9897
rect 12216 9888 12218 9897
rect 12162 9823 12218 9832
rect 11992 9438 12112 9466
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 3602 11928 7686
rect 11992 4078 12020 9438
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 8362 12112 8774
rect 12360 8566 12388 12294
rect 12452 10441 12480 12679
rect 12544 12646 12572 12838
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12530 12472 12586 12481
rect 12530 12407 12586 12416
rect 12544 12170 12572 12407
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12544 11257 12572 11494
rect 12636 11354 12664 12174
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12530 11248 12586 11257
rect 12530 11183 12586 11192
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12452 10062 12480 10367
rect 12728 10266 12756 20046
rect 13268 19994 13320 20000
rect 13372 19922 13584 19938
rect 13360 19916 13584 19922
rect 13412 19910 13584 19916
rect 13360 19858 13412 19864
rect 13452 19848 13504 19854
rect 13556 19836 13584 19910
rect 13636 19848 13688 19854
rect 13556 19808 13636 19836
rect 13452 19790 13504 19796
rect 13636 19790 13688 19796
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12912 18737 12940 19246
rect 13096 18834 13124 19450
rect 13268 19304 13320 19310
rect 13268 19246 13320 19252
rect 13280 18970 13308 19246
rect 13464 19242 13492 19790
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18970 13492 19178
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12898 18728 12954 18737
rect 13634 18728 13690 18737
rect 12898 18663 12954 18672
rect 13188 18698 13584 18714
rect 13188 18692 13596 18698
rect 13188 18686 13544 18692
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12820 17134 12848 17478
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12912 16658 12940 18663
rect 13188 18630 13216 18686
rect 13634 18663 13690 18672
rect 13544 18634 13596 18640
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12912 16182 12940 16594
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 12990 16144 13046 16153
rect 12990 16079 13046 16088
rect 13004 14550 13032 16079
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12820 11898 12848 14418
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12912 14006 12940 14350
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12912 12850 12940 13670
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12544 9625 12572 10066
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12440 9512 12492 9518
rect 12820 9500 12848 11834
rect 12912 9654 12940 12650
rect 13004 11898 13032 13806
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 9654 13032 11494
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12492 9472 12848 9500
rect 12440 9454 12492 9460
rect 13004 9178 13032 9590
rect 12992 9172 13044 9178
rect 12992 9114 13044 9120
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12072 8356 12124 8362
rect 13096 8344 13124 18158
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 14890 13216 15302
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13176 14544 13228 14550
rect 13176 14486 13228 14492
rect 12072 8298 12124 8304
rect 13004 8316 13124 8344
rect 12084 7886 12112 8298
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12360 7546 12388 7890
rect 13004 7546 13032 8316
rect 13188 8242 13216 14486
rect 13280 12714 13308 18566
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13372 13297 13400 16934
rect 13452 14952 13504 14958
rect 13450 14920 13452 14929
rect 13504 14920 13506 14929
rect 13450 14855 13506 14864
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13358 13288 13414 13297
rect 13464 13258 13492 14350
rect 13358 13223 13414 13232
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 13268 11280 13320 11286
rect 13268 11222 13320 11228
rect 13280 9586 13308 11222
rect 13372 10130 13400 12786
rect 13464 12594 13492 13194
rect 13556 12850 13584 18090
rect 13648 14793 13676 18663
rect 13740 18086 13768 22520
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14200 20346 14228 20402
rect 14016 20330 14228 20346
rect 14004 20324 14228 20330
rect 14056 20318 14228 20324
rect 14004 20266 14056 20272
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13634 14784 13690 14793
rect 13634 14719 13690 14728
rect 13740 14634 13768 16050
rect 13832 15473 13860 20198
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 13910 19544 13966 19553
rect 13910 19479 13966 19488
rect 13924 16946 13952 19479
rect 14200 18290 14228 19654
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14016 17134 14044 18226
rect 14094 18184 14150 18193
rect 14094 18119 14096 18128
rect 14148 18119 14150 18128
rect 14096 18090 14148 18096
rect 14188 17740 14240 17746
rect 14188 17682 14240 17688
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17338 14136 17614
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13924 16918 14044 16946
rect 13910 16824 13966 16833
rect 13910 16759 13966 16768
rect 13818 15464 13874 15473
rect 13818 15399 13874 15408
rect 13832 14657 13860 15399
rect 13648 14606 13768 14634
rect 13818 14648 13874 14657
rect 13648 13462 13676 14606
rect 13818 14583 13874 14592
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13636 13456 13688 13462
rect 13636 13398 13688 13404
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13648 12714 13676 13398
rect 13636 12708 13688 12714
rect 13636 12650 13688 12656
rect 13464 12566 13676 12594
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13464 11354 13492 12242
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13648 9602 13676 12566
rect 13740 12374 13768 13874
rect 13832 12374 13860 14418
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11150 13768 11698
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13740 10810 13768 11086
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13464 9574 13676 9602
rect 13464 9382 13492 9574
rect 13542 9480 13598 9489
rect 13542 9415 13598 9424
rect 13556 9382 13584 9415
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13832 8906 13860 11766
rect 13924 8906 13952 16759
rect 14016 15994 14044 16918
rect 14016 15966 14136 15994
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 14016 9042 14044 15846
rect 14108 13190 14136 15966
rect 14200 14618 14228 17682
rect 14292 17241 14320 22520
rect 14844 20618 14872 22520
rect 14660 20590 14872 20618
rect 14372 20324 14424 20330
rect 14372 20266 14424 20272
rect 14384 20233 14412 20266
rect 14370 20224 14426 20233
rect 14370 20159 14426 20168
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18290 14412 19110
rect 14660 18630 14688 20590
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14278 17232 14334 17241
rect 14278 17167 14334 17176
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16250 14412 16934
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14476 16096 14504 17070
rect 14384 16068 14504 16096
rect 14278 15600 14334 15609
rect 14278 15535 14280 15544
rect 14332 15535 14334 15544
rect 14280 15506 14332 15512
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14384 13002 14412 16068
rect 14464 15972 14516 15978
rect 14464 15914 14516 15920
rect 14476 15570 14504 15914
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14476 14482 14504 14826
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14568 13938 14596 17138
rect 14752 16590 14780 20402
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15106 19408 15162 19417
rect 15106 19343 15162 19352
rect 15120 19310 15148 19343
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15304 18222 15332 19654
rect 15292 18216 15344 18222
rect 15292 18158 15344 18164
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15212 16658 15240 17750
rect 15396 17490 15424 22520
rect 15566 20496 15622 20505
rect 15566 20431 15622 20440
rect 15580 20330 15608 20431
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15488 18154 15516 18906
rect 15566 18864 15622 18873
rect 15566 18799 15622 18808
rect 15580 18154 15608 18799
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15568 18148 15620 18154
rect 15568 18090 15620 18096
rect 15396 17462 15516 17490
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 16266 14780 16526
rect 14752 16250 14872 16266
rect 14752 16244 14884 16250
rect 14752 16238 14832 16244
rect 14832 16186 14884 16192
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15212 15162 15240 15642
rect 15304 15570 15332 16118
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 14648 14884 14700 14890
rect 14648 14826 14700 14832
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14108 12974 14412 13002
rect 14108 9382 14136 12974
rect 14476 12832 14504 13806
rect 14660 13025 14688 14826
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15304 14618 15332 14962
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14752 13530 14780 14418
rect 15304 14346 15332 14418
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14646 13016 14702 13025
rect 14646 12951 14702 12960
rect 14292 12804 14504 12832
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14200 11014 14228 12378
rect 14292 12102 14320 12804
rect 14660 12730 14688 12951
rect 14476 12702 14688 12730
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 13820 8900 13872 8906
rect 13820 8842 13872 8848
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 14016 8838 14044 8978
rect 14200 8974 14228 9522
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 14200 8566 14228 8910
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 13096 8214 13216 8242
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12084 5166 12112 6054
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 12070 3496 12126 3505
rect 12070 3431 12126 3440
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11256 1958 11468 1986
rect 10968 1216 11020 1222
rect 10968 1158 11020 1164
rect 11440 480 11468 1958
rect 12084 480 12112 3431
rect 12360 2990 12388 6870
rect 12636 6798 12664 7414
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12820 6934 12848 7142
rect 12808 6928 12860 6934
rect 12808 6870 12860 6876
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12452 5710 12480 6326
rect 12728 5914 12756 6666
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5914 12848 6054
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 13004 5166 13032 7482
rect 13096 6934 13124 8214
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13188 7002 13216 7822
rect 14108 7410 14136 7822
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 14016 6934 14044 7278
rect 14292 7002 14320 11154
rect 14384 11150 14412 12310
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 13740 5166 13768 6870
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13924 5710 13952 6122
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5370 13952 5646
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 14016 5030 14044 6870
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14200 6458 14228 6598
rect 14292 6458 14320 6734
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 5234 14228 6190
rect 14292 5710 14320 6394
rect 14384 6254 14412 11086
rect 14476 7410 14504 12702
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 9518 14596 11290
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14188 5228 14240 5234
rect 14188 5170 14240 5176
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14292 5114 14320 5170
rect 14200 5086 14320 5114
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12544 4554 12572 4762
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12544 4078 12572 4490
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12544 1034 12572 3062
rect 12636 2514 12664 4966
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 13176 2100 13228 2106
rect 13176 2042 13228 2048
rect 12544 1006 12664 1034
rect 12636 480 12664 1006
rect 13188 480 13216 2042
rect 13740 480 13768 2790
rect 13832 2582 13860 4694
rect 13924 4146 13952 4966
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 4026 14044 4966
rect 14200 4554 14228 5086
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14292 4758 14320 4966
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13924 3998 14044 4026
rect 13924 3602 13952 3998
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 3738 14044 3878
rect 14108 3738 14136 4422
rect 14292 4214 14320 4558
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 14292 3618 14320 4014
rect 14384 3738 14412 5782
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 14004 3596 14056 3602
rect 14292 3590 14412 3618
rect 14004 3538 14056 3544
rect 14016 3398 14044 3538
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 13924 2514 13952 3334
rect 14384 3097 14412 3590
rect 14476 3534 14504 6258
rect 14568 5778 14596 9318
rect 14660 7818 14688 12310
rect 14752 12102 14780 13330
rect 15212 13274 15240 13874
rect 15304 13870 15332 14282
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15120 13246 15240 13274
rect 15120 12986 15148 13246
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12442 15240 13126
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14752 10130 14780 12038
rect 15304 11914 15332 12582
rect 15396 12442 15424 15506
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15120 11898 15332 11914
rect 15108 11892 15332 11898
rect 15160 11886 15332 11892
rect 15108 11834 15160 11840
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15304 11257 15332 11698
rect 15382 11384 15438 11393
rect 15382 11319 15438 11328
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 15396 11150 15424 11319
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 15304 10062 15332 10542
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15488 9654 15516 17462
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15580 16726 15608 16934
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 12714 15608 15846
rect 15672 15366 15700 20198
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15856 19242 15884 19722
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15844 18216 15896 18222
rect 15844 18158 15896 18164
rect 15856 16017 15884 18158
rect 15842 16008 15898 16017
rect 15842 15943 15898 15952
rect 15842 15736 15898 15745
rect 15842 15671 15898 15680
rect 15856 15638 15884 15671
rect 15844 15632 15896 15638
rect 15844 15574 15896 15580
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 13734 15700 15302
rect 15948 14770 15976 22520
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16040 18426 16068 19858
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16132 19553 16160 19790
rect 16118 19544 16174 19553
rect 16118 19479 16174 19488
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 16132 18766 16160 19246
rect 16120 18760 16172 18766
rect 16120 18702 16172 18708
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 16132 17678 16160 18702
rect 16028 17672 16080 17678
rect 16028 17614 16080 17620
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 15764 14742 15976 14770
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15672 11642 15700 13330
rect 15764 11937 15792 14742
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15856 13920 15884 14554
rect 16040 14550 16068 17614
rect 16132 16590 16160 17614
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15856 13892 15976 13920
rect 15844 13456 15896 13462
rect 15844 13398 15896 13404
rect 15750 11928 15806 11937
rect 15750 11863 15806 11872
rect 15580 11614 15700 11642
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 8537 14780 9454
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14738 8528 14794 8537
rect 14738 8463 14794 8472
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14752 5914 14780 8463
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15304 7410 15332 9318
rect 15396 9178 15424 9318
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15580 8276 15608 11614
rect 15658 11520 15714 11529
rect 15658 11455 15714 11464
rect 15672 11218 15700 11455
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15658 9480 15714 9489
rect 15658 9415 15660 9424
rect 15712 9415 15714 9424
rect 15660 9386 15712 9392
rect 15764 8634 15792 9522
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15672 8430 15700 8570
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15580 8248 15700 8276
rect 15672 7818 15700 8248
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15212 6322 15240 6802
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14370 3088 14426 3097
rect 14280 3052 14332 3058
rect 14370 3023 14372 3032
rect 14280 2994 14332 3000
rect 14424 3023 14426 3032
rect 14372 2994 14424 3000
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14292 480 14320 2994
rect 14568 2854 14596 5238
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14752 3942 14780 4150
rect 14740 3936 14792 3942
rect 14646 3904 14702 3913
rect 14740 3878 14792 3884
rect 14646 3839 14702 3848
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14660 2258 14688 3839
rect 14752 2922 14780 3878
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3097 14872 3402
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 14660 2230 14872 2258
rect 14844 480 14872 2230
rect 15396 480 15424 3674
rect 15488 3534 15516 3674
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15580 2990 15608 7142
rect 15672 5166 15700 7754
rect 15856 7426 15884 13398
rect 15948 11150 15976 13892
rect 16026 13832 16082 13841
rect 16026 13767 16082 13776
rect 16040 13462 16068 13767
rect 16028 13456 16080 13462
rect 16028 13398 16080 13404
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 11626 16068 13194
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 16132 11506 16160 12650
rect 16040 11478 16160 11506
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 15948 10198 15976 11086
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 16040 8022 16068 11478
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 16132 7886 16160 8570
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15764 7398 15884 7426
rect 15660 5160 15712 5166
rect 15660 5102 15712 5108
rect 15764 5030 15792 7398
rect 15948 7342 15976 7686
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16132 6934 16160 7822
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16224 5098 16252 20198
rect 16500 19281 16528 22520
rect 17052 19394 17080 22520
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17144 19514 17172 19790
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 16868 19366 17080 19394
rect 16486 19272 16542 19281
rect 16486 19207 16542 19216
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16776 18902 16804 19110
rect 16764 18896 16816 18902
rect 16764 18838 16816 18844
rect 16776 18290 16804 18838
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17134 16528 17478
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16500 16250 16528 16526
rect 16868 16454 16896 19366
rect 16948 19304 17000 19310
rect 16948 19246 17000 19252
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16500 15502 16528 16050
rect 16764 16040 16816 16046
rect 16764 15982 16816 15988
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16396 15496 16448 15502
rect 16394 15464 16396 15473
rect 16488 15496 16540 15502
rect 16448 15464 16450 15473
rect 16488 15438 16540 15444
rect 16394 15399 16450 15408
rect 16302 15056 16358 15065
rect 16302 14991 16358 15000
rect 16316 13870 16344 14991
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16408 14006 16436 14486
rect 16396 14000 16448 14006
rect 16396 13942 16448 13948
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 9058 16344 13670
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12986 16436 13262
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16500 10606 16528 15438
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 14958 16620 15302
rect 16684 15026 16712 15846
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16776 14226 16804 15982
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16868 15706 16896 15846
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16960 15162 16988 19246
rect 17132 19236 17184 19242
rect 17132 19178 17184 19184
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16684 14198 16804 14226
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 13297 16620 13330
rect 16578 13288 16634 13297
rect 16578 13223 16634 13232
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16396 10192 16448 10198
rect 16396 10134 16448 10140
rect 16408 9178 16436 10134
rect 16500 9994 16528 10542
rect 16592 10266 16620 12174
rect 16684 11354 16712 14198
rect 16762 12880 16818 12889
rect 16762 12815 16818 12824
rect 16776 12782 16804 12815
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16776 11121 16804 11494
rect 16868 11286 16896 14962
rect 16856 11280 16908 11286
rect 16856 11222 16908 11228
rect 16762 11112 16818 11121
rect 16762 11047 16818 11056
rect 16868 10810 16896 11222
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16960 10810 16988 11086
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16960 10538 16988 10746
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 17052 9110 17080 17002
rect 17144 14278 17172 19178
rect 17236 18970 17264 20334
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17132 14272 17184 14278
rect 17132 14214 17184 14220
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17144 11762 17172 12242
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17144 9897 17172 10474
rect 17130 9888 17186 9897
rect 17130 9823 17186 9832
rect 17040 9104 17092 9110
rect 16316 9030 16436 9058
rect 17040 9046 17092 9052
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16316 7478 16344 8434
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16212 5092 16264 5098
rect 16212 5034 16264 5040
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 16224 4826 16252 5034
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 15764 4729 15792 4762
rect 15750 4720 15806 4729
rect 15750 4655 15806 4664
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15672 3194 15700 3538
rect 15764 3534 15792 4014
rect 16408 3602 16436 9030
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16776 8362 16804 8502
rect 17236 8430 17264 17478
rect 17328 12782 17356 19722
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 17512 16250 17540 18158
rect 17604 17354 17632 18566
rect 17696 17542 17724 22520
rect 18142 22264 18198 22273
rect 18142 22199 18198 22208
rect 18050 21720 18106 21729
rect 18050 21655 18106 21664
rect 17958 21312 18014 21321
rect 17958 21247 18014 21256
rect 17972 20942 18000 21247
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 18064 20874 18092 21655
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 18156 20806 18184 22199
rect 18248 20890 18276 22520
rect 18340 21146 18368 22607
rect 18786 22520 18842 23000
rect 19338 22520 19394 23000
rect 19890 22520 19946 23000
rect 20442 22520 20498 23000
rect 20994 22520 21050 23000
rect 21546 22520 21602 23000
rect 22098 22520 22154 23000
rect 22650 22520 22706 23000
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18696 21004 18748 21010
rect 18696 20946 18748 20952
rect 18248 20862 18644 20890
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17684 17536 17736 17542
rect 17684 17478 17736 17484
rect 17604 17326 17724 17354
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17406 16144 17462 16153
rect 17406 16079 17462 16088
rect 17420 16046 17448 16079
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17406 15736 17462 15745
rect 17406 15671 17462 15680
rect 17420 15638 17448 15671
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17512 15502 17540 16186
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17512 14958 17540 15438
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17604 13258 17632 17002
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 10742 17448 12582
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17512 10130 17540 13126
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17420 8430 17448 9862
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 6662 16528 7346
rect 16776 6866 16804 8298
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16500 6254 16528 6598
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 15948 480 15976 1906
rect 16500 480 16528 6054
rect 16776 5710 16804 6802
rect 17132 6724 17184 6730
rect 17132 6666 17184 6672
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 16776 4078 16804 5646
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16592 2990 16620 3878
rect 16776 3738 16804 3878
rect 16764 3732 16816 3738
rect 16764 3674 16816 3680
rect 16868 3058 16896 6122
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 17052 480 17080 3334
rect 17144 2514 17172 6666
rect 17512 6254 17540 8230
rect 17604 7954 17632 11494
rect 17696 10985 17724 17326
rect 17788 16697 17816 20198
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17880 17649 17908 19994
rect 18052 19916 18104 19922
rect 18052 19858 18104 19864
rect 17958 18864 18014 18873
rect 17958 18799 17960 18808
rect 18012 18799 18014 18808
rect 17960 18770 18012 18776
rect 17866 17640 17922 17649
rect 17866 17575 17922 17584
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17774 16688 17830 16697
rect 17774 16623 17830 16632
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 15570 17816 16390
rect 17880 16153 17908 17206
rect 18064 17082 18092 19858
rect 18156 19825 18184 20538
rect 18142 19816 18198 19825
rect 18142 19751 18198 19760
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18156 18630 18184 18770
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 17972 17054 18092 17082
rect 17866 16144 17922 16153
rect 17866 16079 17922 16088
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17880 15609 17908 15642
rect 17866 15600 17922 15609
rect 17776 15564 17828 15570
rect 17866 15535 17922 15544
rect 17776 15506 17828 15512
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14482 17908 14894
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17880 12782 17908 14418
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17880 12306 17908 12718
rect 17972 12646 18000 17054
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16794 18092 16934
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18052 16652 18104 16658
rect 18052 16594 18104 16600
rect 18064 15065 18092 16594
rect 18156 15609 18184 18022
rect 18616 17785 18644 20862
rect 18708 20777 18736 20946
rect 18694 20768 18750 20777
rect 18694 20703 18750 20712
rect 18800 18737 18828 22520
rect 18972 18760 19024 18766
rect 18786 18728 18842 18737
rect 18972 18702 19024 18708
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 18786 18663 18842 18672
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18694 18456 18750 18465
rect 18694 18391 18750 18400
rect 18602 17776 18658 17785
rect 18602 17711 18658 17720
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18616 17202 18644 17546
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18616 16726 18644 17138
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18616 16114 18644 16662
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18142 15600 18198 15609
rect 18142 15535 18198 15544
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18050 15056 18106 15065
rect 18050 14991 18106 15000
rect 18708 14822 18736 18391
rect 18800 17882 18828 18566
rect 18788 17876 18840 17882
rect 18788 17818 18840 17824
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18892 17338 18920 17614
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 18786 17096 18842 17105
rect 18786 17031 18842 17040
rect 18800 15366 18828 17031
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18786 14240 18842 14249
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17972 11830 18000 12242
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17682 10976 17738 10985
rect 17682 10911 17738 10920
rect 17684 10056 17736 10062
rect 17682 10024 17684 10033
rect 17736 10024 17738 10033
rect 17682 9959 17738 9968
rect 17788 9897 17816 11562
rect 17972 11354 18000 11766
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17958 11248 18014 11257
rect 17958 11183 18014 11192
rect 17868 10600 17920 10606
rect 17868 10542 17920 10548
rect 17880 9926 17908 10542
rect 17972 10146 18000 11183
rect 18064 11150 18092 12378
rect 18156 11694 18184 14214
rect 18282 14172 18578 14192
rect 18786 14175 18842 14184
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18800 14074 18828 14175
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18788 13932 18840 13938
rect 18788 13874 18840 13880
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13530 18276 13670
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18602 13288 18658 13297
rect 18602 13223 18658 13232
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18144 11688 18196 11694
rect 18340 11665 18368 11698
rect 18144 11630 18196 11636
rect 18326 11656 18382 11665
rect 18326 11591 18382 11600
rect 18144 11212 18196 11218
rect 18144 11154 18196 11160
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17972 10118 18092 10146
rect 17960 9988 18012 9994
rect 17960 9930 18012 9936
rect 17868 9920 17920 9926
rect 17774 9888 17830 9897
rect 17868 9862 17920 9868
rect 17774 9823 17830 9832
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 8974 17724 9522
rect 17788 9178 17816 9823
rect 17972 9518 18000 9930
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17958 9072 18014 9081
rect 17788 9030 17958 9058
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 7993 17724 8910
rect 17788 8838 17816 9030
rect 17958 9007 18014 9016
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17682 7984 17738 7993
rect 17592 7948 17644 7954
rect 17682 7919 17738 7928
rect 17592 7890 17644 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17696 7274 17724 7822
rect 17684 7268 17736 7274
rect 17684 7210 17736 7216
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6322 17632 6666
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17512 4078 17540 6190
rect 17696 4593 17724 7210
rect 17788 5846 17816 7822
rect 17776 5840 17828 5846
rect 17880 5817 17908 8842
rect 18064 8378 18092 10118
rect 18156 9489 18184 11154
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18616 9654 18644 13223
rect 18800 12850 18828 13874
rect 18878 13832 18934 13841
rect 18878 13767 18934 13776
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18708 12073 18736 12650
rect 18694 12064 18750 12073
rect 18694 11999 18750 12008
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18142 9480 18198 9489
rect 18142 9415 18198 9424
rect 18156 8430 18184 9415
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17972 8350 18092 8378
rect 18144 8424 18196 8430
rect 18144 8366 18196 8372
rect 17972 8022 18000 8350
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 18064 8090 18092 8230
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 18050 7984 18106 7993
rect 18050 7919 18106 7928
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17776 5782 17828 5788
rect 17866 5808 17922 5817
rect 17788 4622 17816 5782
rect 17866 5743 17922 5752
rect 17776 4616 17828 4622
rect 17682 4584 17738 4593
rect 17776 4558 17828 4564
rect 17682 4519 17738 4528
rect 17500 4072 17552 4078
rect 17500 4014 17552 4020
rect 17788 3534 17816 4558
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 2582 17908 3402
rect 17972 2922 18000 7686
rect 18064 7410 18092 7919
rect 18248 7732 18276 8502
rect 18604 8356 18656 8362
rect 18708 8344 18736 11018
rect 18800 10010 18828 11086
rect 18892 10810 18920 13767
rect 18984 12753 19012 18702
rect 19168 18222 19196 18702
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19168 17202 19196 18158
rect 19246 18048 19302 18057
rect 19246 17983 19302 17992
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 16250 19196 16526
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19260 16130 19288 17983
rect 19352 17270 19380 22520
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19536 19514 19564 19858
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17746 19472 18022
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19340 17264 19392 17270
rect 19340 17206 19392 17212
rect 19168 16102 19288 16130
rect 19168 12986 19196 16102
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19260 15366 19288 15982
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19260 14958 19288 15302
rect 19248 14952 19300 14958
rect 19248 14894 19300 14900
rect 19260 13938 19288 14894
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 13433 19288 13670
rect 19352 13462 19380 15914
rect 19536 13870 19564 18090
rect 19628 15706 19656 20402
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19720 17814 19748 20334
rect 19708 17808 19760 17814
rect 19708 17750 19760 17756
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19340 13456 19392 13462
rect 19246 13424 19302 13433
rect 19340 13398 19392 13404
rect 19246 13359 19302 13368
rect 19524 13388 19576 13394
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19260 12866 19288 13359
rect 19524 13330 19576 13336
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19352 12986 19380 13262
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19260 12838 19380 12866
rect 19248 12776 19300 12782
rect 18970 12744 19026 12753
rect 19248 12718 19300 12724
rect 18970 12679 19026 12688
rect 19260 12442 19288 12718
rect 19248 12436 19300 12442
rect 19248 12378 19300 12384
rect 19352 12322 19380 12838
rect 19444 12374 19472 13262
rect 19076 12294 19380 12322
rect 19432 12368 19484 12374
rect 19432 12310 19484 12316
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18984 11626 19012 12106
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18800 9982 18920 10010
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18656 8316 18736 8344
rect 18604 8298 18656 8304
rect 18326 8120 18382 8129
rect 18326 8055 18382 8064
rect 18340 7818 18368 8055
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18156 7704 18276 7732
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18064 6934 18092 7346
rect 18052 6928 18104 6934
rect 18052 6870 18104 6876
rect 18156 5710 18184 7704
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18616 6225 18644 8298
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7721 18736 7890
rect 18694 7712 18750 7721
rect 18694 7647 18750 7656
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18602 6216 18658 6225
rect 18602 6151 18658 6160
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18064 5273 18092 5306
rect 18050 5264 18106 5273
rect 18050 5199 18106 5208
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4865 18092 4966
rect 18050 4856 18106 4865
rect 18050 4791 18106 4800
rect 18156 4758 18184 5510
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18708 5234 18736 6870
rect 18696 5228 18748 5234
rect 18524 5188 18696 5216
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18524 4622 18552 5188
rect 18696 5170 18748 5176
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3194 18092 3878
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18156 2990 18184 4422
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18616 3534 18644 4694
rect 18800 3602 18828 9862
rect 18892 7177 18920 9982
rect 18878 7168 18934 7177
rect 18878 7103 18934 7112
rect 18892 5846 18920 7103
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18878 5128 18934 5137
rect 18878 5063 18934 5072
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18788 3596 18840 3602
rect 18788 3538 18840 3544
rect 18604 3528 18656 3534
rect 18708 3505 18736 3538
rect 18604 3470 18656 3476
rect 18694 3496 18750 3505
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18616 3058 18644 3470
rect 18694 3431 18750 3440
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 17868 2576 17920 2582
rect 17868 2518 17920 2524
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 480 17724 2246
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 17972 1601 18000 1974
rect 17958 1592 18014 1601
rect 17958 1527 18014 1536
rect 18156 1442 18184 2790
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1414 18276 1442
rect 18144 1352 18196 1358
rect 18144 1294 18196 1300
rect 18052 1284 18104 1290
rect 18052 1226 18104 1232
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 17972 1057 18000 1158
rect 17958 1048 18014 1057
rect 17958 983 18014 992
rect 18064 649 18092 1226
rect 18050 640 18106 649
rect 18050 575 18106 584
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6458 0 6514 480
rect 7010 0 7066 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 12070 0 12126 480
rect 12622 0 12678 480
rect 13174 0 13230 480
rect 13726 0 13782 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17682 0 17738 480
rect 18156 241 18184 1294
rect 18248 480 18276 1414
rect 18800 480 18828 2586
rect 18892 2553 18920 5063
rect 18984 2938 19012 11562
rect 19076 7426 19104 12294
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19260 11098 19288 11630
rect 19536 11354 19564 13330
rect 19524 11348 19576 11354
rect 19524 11290 19576 11296
rect 19260 11070 19380 11098
rect 19628 11082 19656 14418
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 13530 19748 14350
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19720 11694 19748 12922
rect 19812 12345 19840 17478
rect 19904 15450 19932 22520
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19996 16250 20024 19178
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19904 15422 20024 15450
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 14657 19932 15302
rect 19890 14648 19946 14657
rect 19890 14583 19946 14592
rect 19996 13954 20024 15422
rect 20088 14074 20116 19110
rect 20180 16182 20208 19314
rect 20364 18290 20392 20470
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 20272 16658 20300 18158
rect 20456 17542 20484 22520
rect 21008 18902 21036 22520
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20812 17536 20864 17542
rect 21560 17490 21588 22520
rect 22112 17542 22140 22520
rect 20812 17478 20864 17484
rect 20444 17264 20496 17270
rect 20444 17206 20496 17212
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20180 15162 20208 16118
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 19996 13926 20116 13954
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19798 12336 19854 12345
rect 19798 12271 19854 12280
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19246 10976 19302 10985
rect 19246 10911 19302 10920
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19168 9586 19196 10610
rect 19260 10146 19288 10911
rect 19352 10810 19380 11070
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19260 10118 19472 10146
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19248 9988 19300 9994
rect 19248 9930 19300 9936
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19156 9036 19208 9042
rect 19156 8978 19208 8984
rect 19168 7818 19196 8978
rect 19260 8090 19288 9930
rect 19352 9722 19380 9998
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19352 9178 19380 9658
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19248 7880 19300 7886
rect 19300 7840 19380 7868
rect 19248 7822 19300 7828
rect 19156 7812 19208 7818
rect 19156 7754 19208 7760
rect 19168 7546 19196 7754
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19076 7398 19196 7426
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 19076 6662 19104 7210
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 3058 19104 6598
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19168 2961 19196 7398
rect 19260 6769 19288 7686
rect 19352 7478 19380 7840
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19246 6760 19302 6769
rect 19246 6695 19302 6704
rect 19444 6610 19472 10118
rect 19536 8566 19564 10202
rect 19812 9450 19840 12038
rect 19904 11150 19932 13262
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10538 19932 11086
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19890 8392 19946 8401
rect 19890 8327 19892 8336
rect 19944 8327 19946 8336
rect 19892 8298 19944 8304
rect 19996 7342 20024 13806
rect 20088 10577 20116 13926
rect 20074 10568 20130 10577
rect 20074 10503 20130 10512
rect 20180 10470 20208 14350
rect 20168 10464 20220 10470
rect 20272 10441 20300 15846
rect 20364 12170 20392 17002
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20456 10690 20484 17206
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20364 10662 20484 10690
rect 20168 10406 20220 10412
rect 20258 10432 20314 10441
rect 20258 10367 20314 10376
rect 20364 9761 20392 10662
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20350 9752 20406 9761
rect 20350 9687 20406 9696
rect 20456 9654 20484 10474
rect 20548 10441 20576 13330
rect 20824 12209 20852 17478
rect 20916 17462 21588 17490
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 20810 12200 20866 12209
rect 20810 12135 20866 12144
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11898 20668 12038
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20916 11801 20944 17462
rect 22664 17338 22692 22520
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 22652 17332 22704 17338
rect 22652 17274 22704 17280
rect 20902 11792 20958 11801
rect 20902 11727 20958 11736
rect 20534 10432 20590 10441
rect 20534 10367 20590 10376
rect 20444 9648 20496 9654
rect 20444 9590 20496 9596
rect 20548 8498 20576 10367
rect 21008 10169 21036 17274
rect 20994 10160 21050 10169
rect 20994 10095 21050 10104
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20628 8492 20680 8498
rect 20628 8434 20680 8440
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19260 6582 19472 6610
rect 19260 3738 19288 6582
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19708 6112 19760 6118
rect 19708 6054 19760 6060
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19628 3924 19656 5578
rect 19720 4570 19748 6054
rect 19812 5914 19840 6054
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 19904 5710 19932 6258
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19904 5098 19932 5646
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19720 4542 19840 4570
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19720 4078 19748 4422
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19628 3896 19748 3924
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19340 3120 19392 3126
rect 19340 3062 19392 3068
rect 19154 2952 19210 2961
rect 18984 2910 19104 2938
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 19076 2009 19104 2910
rect 19154 2887 19210 2896
rect 19062 2000 19118 2009
rect 19062 1935 19118 1944
rect 19352 480 19380 3062
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19628 2514 19656 2790
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19720 762 19748 3896
rect 19812 2854 19840 4542
rect 19904 3942 19932 5034
rect 19892 3936 19944 3942
rect 19996 3913 20024 5578
rect 19892 3878 19944 3884
rect 19982 3904 20038 3913
rect 19982 3839 20038 3848
rect 20088 2990 20116 8230
rect 20536 7336 20588 7342
rect 20536 7278 20588 7284
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 3602 20300 4966
rect 20260 3596 20312 3602
rect 20260 3538 20312 3544
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19720 734 19932 762
rect 19904 480 19932 734
rect 20456 480 20484 5306
rect 20548 4690 20576 7278
rect 20640 6866 20668 8434
rect 21548 7200 21600 7206
rect 21548 7142 21600 7148
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 6322 20668 6802
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5370 20668 6258
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20996 2372 21048 2378
rect 20996 2314 21048 2320
rect 21008 480 21036 2314
rect 21560 480 21588 7142
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22100 3596 22152 3602
rect 22100 3538 22152 3544
rect 22112 480 22140 3538
rect 22664 480 22692 3946
rect 18142 232 18198 241
rect 18142 167 18198 176
rect 18234 0 18290 480
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19890 0 19946 480
rect 20442 0 20498 480
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
<< via2 >>
rect 1766 17040 1822 17096
rect 1582 15000 1638 15056
rect 1398 13524 1454 13560
rect 1398 13504 1400 13524
rect 1400 13504 1452 13524
rect 1452 13504 1454 13524
rect 1398 11600 1454 11656
rect 1858 13948 1860 13968
rect 1860 13948 1912 13968
rect 1912 13948 1914 13968
rect 1858 13912 1914 13948
rect 1674 9968 1730 10024
rect 2594 15972 2650 16008
rect 2594 15952 2596 15972
rect 2596 15952 2648 15972
rect 2648 15952 2650 15972
rect 2870 14320 2926 14376
rect 3054 12164 3110 12200
rect 3054 12144 3056 12164
rect 3056 12144 3108 12164
rect 3108 12144 3110 12164
rect 3514 17176 3570 17232
rect 3330 15408 3386 15464
rect 3422 14456 3478 14512
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4066 17856 4122 17912
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 3698 14320 3754 14376
rect 3606 9560 3662 9616
rect 2042 3068 2044 3088
rect 2044 3068 2096 3088
rect 2096 3068 2098 3088
rect 2042 3032 2098 3068
rect 2870 3440 2926 3496
rect 3054 5752 3110 5808
rect 3054 3712 3110 3768
rect 3974 6840 4030 6896
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 5262 18400 5318 18456
rect 5538 18264 5594 18320
rect 5538 17992 5594 18048
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4802 14356 4804 14376
rect 4804 14356 4856 14376
rect 4856 14356 4858 14376
rect 4802 14320 4858 14356
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4434 11736 4490 11792
rect 4802 10920 4858 10976
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4618 10532 4674 10568
rect 4618 10512 4620 10532
rect 4620 10512 4672 10532
rect 4672 10512 4674 10532
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4802 9444 4858 9480
rect 4802 9424 4804 9444
rect 4804 9424 4856 9444
rect 4856 9424 4858 9444
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4434 8336 4490 8392
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4802 3304 4858 3360
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 5814 14864 5870 14920
rect 5722 14320 5778 14376
rect 5170 3984 5226 4040
rect 5446 11056 5502 11112
rect 5814 10684 5816 10704
rect 5816 10684 5868 10704
rect 5868 10684 5870 10704
rect 5814 10648 5870 10684
rect 5998 17992 6054 18048
rect 6182 12280 6238 12336
rect 6826 18128 6882 18184
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7010 17856 7066 17912
rect 6366 12824 6422 12880
rect 6090 3984 6146 4040
rect 7102 16088 7158 16144
rect 7102 12824 7158 12880
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 7562 15816 7618 15872
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7746 14456 7802 14512
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7470 13504 7526 13560
rect 7562 12960 7618 13016
rect 6826 10104 6882 10160
rect 7102 9696 7158 9752
rect 7286 9560 7342 9616
rect 6642 3984 6698 4040
rect 6918 5072 6974 5128
rect 6826 4120 6882 4176
rect 6918 3168 6974 3224
rect 8298 13640 8354 13696
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 9862 20168 9918 20224
rect 9678 20052 9734 20088
rect 9678 20032 9680 20052
rect 9680 20032 9732 20052
rect 9732 20032 9734 20052
rect 9770 19932 9772 19952
rect 9772 19932 9824 19952
rect 9824 19932 9826 19952
rect 9770 19896 9826 19932
rect 9770 19624 9826 19680
rect 9310 19116 9312 19136
rect 9312 19116 9364 19136
rect 9364 19116 9366 19136
rect 9310 19080 9366 19116
rect 8666 15408 8722 15464
rect 9126 17040 9182 17096
rect 8850 16088 8906 16144
rect 8482 14320 8538 14376
rect 8482 12008 8538 12064
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7930 11192 7986 11248
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8206 9560 8262 9616
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 8390 11464 8446 11520
rect 9586 18400 9642 18456
rect 9310 15000 9366 15056
rect 8850 14864 8906 14920
rect 8758 14728 8814 14784
rect 8758 13912 8814 13968
rect 8942 13776 8998 13832
rect 8758 13096 8814 13152
rect 8666 12552 8722 12608
rect 8758 11192 8814 11248
rect 8298 9324 8300 9344
rect 8300 9324 8352 9344
rect 8352 9324 8354 9344
rect 8298 9288 8354 9324
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7378 5072 7434 5128
rect 7378 2916 7434 2952
rect 7378 2896 7380 2916
rect 7380 2896 7432 2916
rect 7432 2896 7434 2916
rect 7562 3168 7618 3224
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 8482 10784 8538 10840
rect 9034 13504 9090 13560
rect 9126 12416 9182 12472
rect 8482 6840 8538 6896
rect 9126 11328 9182 11384
rect 9678 14220 9680 14240
rect 9680 14220 9732 14240
rect 9732 14220 9734 14240
rect 9678 14184 9734 14220
rect 10138 20032 10194 20088
rect 10046 18808 10102 18864
rect 10046 14592 10102 14648
rect 9954 14048 10010 14104
rect 9402 13504 9458 13560
rect 9770 13504 9826 13560
rect 9402 11464 9458 11520
rect 9954 13640 10010 13696
rect 9954 13232 10010 13288
rect 9862 12960 9918 13016
rect 9770 12824 9826 12880
rect 9678 12008 9734 12064
rect 9218 9460 9220 9480
rect 9220 9460 9272 9480
rect 9272 9460 9274 9480
rect 9218 9424 9274 9460
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7746 3712 7802 3768
rect 8114 3188 8170 3224
rect 8114 3168 8116 3188
rect 8116 3168 8168 3188
rect 8168 3168 8170 3188
rect 8298 3304 8354 3360
rect 8298 3068 8300 3088
rect 8300 3068 8352 3088
rect 8352 3068 8354 3088
rect 8298 3032 8354 3068
rect 7746 2896 7802 2952
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 9586 9288 9642 9344
rect 10046 11464 10102 11520
rect 10046 10260 10102 10296
rect 10046 10240 10048 10260
rect 10048 10240 10100 10260
rect 10100 10240 10102 10260
rect 10782 22480 10838 22536
rect 18326 22616 18382 22672
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10322 20440 10378 20496
rect 10322 19624 10378 19680
rect 10506 19216 10562 19272
rect 10322 18672 10378 18728
rect 10230 14456 10286 14512
rect 9770 3848 9826 3904
rect 10874 19116 10876 19136
rect 10876 19116 10928 19136
rect 10928 19116 10930 19136
rect 10874 19080 10930 19116
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10782 17992 10838 18048
rect 10506 14456 10562 14512
rect 10322 13524 10378 13560
rect 10322 13504 10324 13524
rect 10324 13504 10376 13524
rect 10376 13504 10378 13524
rect 10322 13096 10378 13152
rect 10414 12008 10470 12064
rect 10322 10784 10378 10840
rect 10322 4120 10378 4176
rect 11058 17720 11114 17776
rect 11702 18672 11758 18728
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10966 16632 11022 16688
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11702 16652 11758 16688
rect 11702 16632 11704 16652
rect 11704 16632 11756 16652
rect 11756 16632 11758 16652
rect 10690 11056 10746 11112
rect 10690 10376 10746 10432
rect 10966 14048 11022 14104
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11702 15000 11758 15056
rect 11702 14320 11758 14376
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 10782 4664 10838 4720
rect 10690 4004 10746 4040
rect 10690 3984 10692 4004
rect 10692 3984 10744 4004
rect 10744 3984 10746 4004
rect 11334 13776 11390 13832
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11702 12860 11704 12880
rect 11704 12860 11756 12880
rect 11756 12860 11758 12880
rect 11702 12824 11758 12860
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11794 12008 11850 12064
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 12162 18028 12164 18048
rect 12164 18028 12216 18048
rect 12216 18028 12218 18048
rect 12162 17992 12218 18028
rect 12070 13776 12126 13832
rect 11978 12552 12034 12608
rect 11978 11872 12034 11928
rect 11978 11464 12034 11520
rect 11978 11348 12034 11384
rect 11978 11328 11980 11348
rect 11980 11328 12032 11348
rect 12032 11328 12034 11348
rect 11794 10240 11850 10296
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11978 9580 12034 9616
rect 11978 9560 11980 9580
rect 11980 9560 12032 9580
rect 12032 9560 12034 9580
rect 12162 13368 12218 13424
rect 12162 13232 12218 13288
rect 12530 18708 12532 18728
rect 12532 18708 12584 18728
rect 12584 18708 12586 18728
rect 12530 18672 12586 18708
rect 12346 16088 12402 16144
rect 12530 18028 12532 18048
rect 12532 18028 12584 18048
rect 12584 18028 12586 18048
rect 12530 17992 12586 18028
rect 12438 12688 12494 12744
rect 12162 9868 12164 9888
rect 12164 9868 12216 9888
rect 12216 9868 12218 9888
rect 12162 9832 12218 9868
rect 12530 12416 12586 12472
rect 12530 11192 12586 11248
rect 12438 10376 12494 10432
rect 12898 18672 12954 18728
rect 13634 18672 13690 18728
rect 12990 16088 13046 16144
rect 12530 9560 12586 9616
rect 13450 14900 13452 14920
rect 13452 14900 13504 14920
rect 13504 14900 13506 14920
rect 13450 14864 13506 14900
rect 13358 13232 13414 13288
rect 13634 14728 13690 14784
rect 13910 19488 13966 19544
rect 14094 18148 14150 18184
rect 14094 18128 14096 18148
rect 14096 18128 14148 18148
rect 14148 18128 14150 18148
rect 13910 16768 13966 16824
rect 13818 15408 13874 15464
rect 13818 14592 13874 14648
rect 13542 9424 13598 9480
rect 14370 20168 14426 20224
rect 14278 17176 14334 17232
rect 14278 15564 14334 15600
rect 14278 15544 14280 15564
rect 14280 15544 14332 15564
rect 14332 15544 14334 15564
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 15106 19352 15162 19408
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 15566 20440 15622 20496
rect 15566 18808 15622 18864
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14646 12960 14702 13016
rect 12070 3440 12126 3496
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15382 11328 15438 11384
rect 15290 11192 15346 11248
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 15842 15952 15898 16008
rect 15842 15680 15898 15736
rect 16118 19488 16174 19544
rect 15750 11872 15806 11928
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14738 8472 14794 8528
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15658 11464 15714 11520
rect 15658 9444 15714 9480
rect 15658 9424 15660 9444
rect 15660 9424 15712 9444
rect 15712 9424 15714 9444
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 14370 3052 14426 3088
rect 14370 3032 14372 3052
rect 14372 3032 14424 3052
rect 14424 3032 14426 3052
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14646 3848 14702 3904
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14830 3032 14886 3088
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 16026 13776 16082 13832
rect 16486 19216 16542 19272
rect 16394 15444 16396 15464
rect 16396 15444 16448 15464
rect 16448 15444 16450 15464
rect 16394 15408 16450 15444
rect 16302 15000 16358 15056
rect 16578 13232 16634 13288
rect 16762 12824 16818 12880
rect 16762 11056 16818 11112
rect 17130 9832 17186 9888
rect 15750 4664 15806 4720
rect 18142 22208 18198 22264
rect 18050 21664 18106 21720
rect 17958 21256 18014 21312
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 17406 16088 17462 16144
rect 17406 15680 17462 15736
rect 17958 18828 18014 18864
rect 17958 18808 17960 18828
rect 17960 18808 18012 18828
rect 18012 18808 18014 18828
rect 17866 17584 17922 17640
rect 17774 16632 17830 16688
rect 18142 19760 18198 19816
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 17866 16088 17922 16144
rect 17866 15544 17922 15600
rect 18694 20712 18750 20768
rect 18786 18672 18842 18728
rect 18694 18400 18750 18456
rect 18602 17720 18658 17776
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18142 15544 18198 15600
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18050 15000 18106 15056
rect 18786 17040 18842 17096
rect 17682 10920 17738 10976
rect 17682 10004 17684 10024
rect 17684 10004 17736 10024
rect 17736 10004 17738 10024
rect 17682 9968 17738 10004
rect 17958 11192 18014 11248
rect 18786 14184 18842 14240
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18602 13232 18658 13288
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18326 11600 18382 11656
rect 17774 9832 17830 9888
rect 17958 9016 18014 9072
rect 17682 7928 17738 7984
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18878 13776 18934 13832
rect 18694 12008 18750 12064
rect 18142 9424 18198 9480
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18050 7928 18106 7984
rect 17866 5752 17922 5808
rect 17682 4528 17738 4584
rect 19246 17992 19302 18048
rect 19246 13368 19302 13424
rect 18970 12688 19026 12744
rect 18326 8064 18382 8120
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18694 7656 18750 7712
rect 18602 6160 18658 6216
rect 18050 5208 18106 5264
rect 18050 4800 18106 4856
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18878 7112 18934 7168
rect 18878 5072 18934 5128
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18694 3440 18750 3496
rect 17958 1536 18014 1592
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 17958 992 18014 1048
rect 18050 584 18106 640
rect 19890 14592 19946 14648
rect 19798 12280 19854 12336
rect 19246 10920 19302 10976
rect 19246 6704 19302 6760
rect 19890 8356 19946 8392
rect 19890 8336 19892 8356
rect 19892 8336 19944 8356
rect 19944 8336 19946 8356
rect 20074 10512 20130 10568
rect 20258 10376 20314 10432
rect 20350 9696 20406 9752
rect 20810 12144 20866 12200
rect 20902 11736 20958 11792
rect 20534 10376 20590 10432
rect 20994 10104 21050 10160
rect 18878 2488 18934 2544
rect 19154 2896 19210 2952
rect 19062 1944 19118 2000
rect 19982 3848 20038 3904
rect 18142 176 18198 232
<< metal3 >>
rect 18321 22674 18387 22677
rect 22520 22674 23000 22704
rect 18321 22672 23000 22674
rect 18321 22616 18326 22672
rect 18382 22616 23000 22672
rect 18321 22614 23000 22616
rect 18321 22611 18387 22614
rect 22520 22584 23000 22614
rect 10777 22540 10843 22541
rect 10726 22538 10732 22540
rect 10686 22478 10732 22538
rect 10796 22536 10843 22540
rect 10838 22480 10843 22536
rect 10726 22476 10732 22478
rect 10796 22476 10843 22480
rect 10777 22475 10843 22476
rect 18137 22266 18203 22269
rect 22520 22266 23000 22296
rect 18137 22264 23000 22266
rect 18137 22208 18142 22264
rect 18198 22208 23000 22264
rect 18137 22206 23000 22208
rect 18137 22203 18203 22206
rect 22520 22176 23000 22206
rect 18045 21722 18111 21725
rect 22520 21722 23000 21752
rect 18045 21720 23000 21722
rect 18045 21664 18050 21720
rect 18106 21664 23000 21720
rect 18045 21662 23000 21664
rect 18045 21659 18111 21662
rect 22520 21632 23000 21662
rect 17953 21314 18019 21317
rect 22520 21314 23000 21344
rect 17953 21312 23000 21314
rect 17953 21256 17958 21312
rect 18014 21256 23000 21312
rect 17953 21254 23000 21256
rect 17953 21251 18019 21254
rect 22520 21224 23000 21254
rect 18689 20770 18755 20773
rect 22520 20770 23000 20800
rect 18689 20768 23000 20770
rect 18689 20712 18694 20768
rect 18750 20712 23000 20768
rect 18689 20710 23000 20712
rect 18689 20707 18755 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22520 20680 23000 20710
rect 18270 20639 18590 20640
rect 10317 20498 10383 20501
rect 15561 20498 15627 20501
rect 10317 20496 15627 20498
rect 10317 20440 10322 20496
rect 10378 20440 15566 20496
rect 15622 20440 15627 20496
rect 10317 20438 15627 20440
rect 10317 20435 10383 20438
rect 15561 20435 15627 20438
rect 22520 20362 23000 20392
rect 14598 20302 23000 20362
rect 9857 20226 9923 20229
rect 14365 20226 14431 20229
rect 9857 20224 14431 20226
rect 9857 20168 9862 20224
rect 9918 20168 14370 20224
rect 14426 20168 14431 20224
rect 9857 20166 14431 20168
rect 9857 20163 9923 20166
rect 14365 20163 14431 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 9673 20090 9739 20093
rect 10133 20090 10199 20093
rect 9673 20088 10199 20090
rect 9673 20032 9678 20088
rect 9734 20032 10138 20088
rect 10194 20032 10199 20088
rect 9673 20030 10199 20032
rect 9673 20027 9739 20030
rect 10133 20027 10199 20030
rect 9765 19954 9831 19957
rect 14598 19954 14658 20302
rect 22520 20272 23000 20302
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 9765 19952 14658 19954
rect 9765 19896 9770 19952
rect 9826 19896 14658 19952
rect 9765 19894 14658 19896
rect 9765 19891 9831 19894
rect 18137 19818 18203 19821
rect 22520 19818 23000 19848
rect 18137 19816 23000 19818
rect 18137 19760 18142 19816
rect 18198 19760 23000 19816
rect 18137 19758 23000 19760
rect 18137 19755 18203 19758
rect 22520 19728 23000 19758
rect 9765 19682 9831 19685
rect 10317 19682 10383 19685
rect 9765 19680 10383 19682
rect 9765 19624 9770 19680
rect 9826 19624 10322 19680
rect 10378 19624 10383 19680
rect 9765 19622 10383 19624
rect 9765 19619 9831 19622
rect 10317 19619 10383 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 13905 19546 13971 19549
rect 16113 19546 16179 19549
rect 13905 19544 16179 19546
rect 13905 19488 13910 19544
rect 13966 19488 16118 19544
rect 16174 19488 16179 19544
rect 13905 19486 16179 19488
rect 13905 19483 13971 19486
rect 16113 19483 16179 19486
rect 15101 19410 15167 19413
rect 22520 19410 23000 19440
rect 15101 19408 23000 19410
rect 15101 19352 15106 19408
rect 15162 19352 23000 19408
rect 15101 19350 23000 19352
rect 15101 19347 15167 19350
rect 22520 19320 23000 19350
rect 10501 19274 10567 19277
rect 16481 19274 16547 19277
rect 10501 19272 16547 19274
rect 10501 19216 10506 19272
rect 10562 19216 16486 19272
rect 16542 19216 16547 19272
rect 10501 19214 16547 19216
rect 10501 19211 10567 19214
rect 16481 19211 16547 19214
rect 9305 19138 9371 19141
rect 10869 19138 10935 19141
rect 9305 19136 10935 19138
rect 9305 19080 9310 19136
rect 9366 19080 10874 19136
rect 10930 19080 10935 19136
rect 9305 19078 10935 19080
rect 9305 19075 9371 19078
rect 10869 19075 10935 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 10041 18866 10107 18869
rect 15561 18866 15627 18869
rect 10041 18864 15627 18866
rect 10041 18808 10046 18864
rect 10102 18808 15566 18864
rect 15622 18808 15627 18864
rect 10041 18806 15627 18808
rect 10041 18803 10107 18806
rect 15561 18803 15627 18806
rect 17953 18866 18019 18869
rect 22520 18866 23000 18896
rect 17953 18864 23000 18866
rect 17953 18808 17958 18864
rect 18014 18808 23000 18864
rect 17953 18806 23000 18808
rect 17953 18803 18019 18806
rect 22520 18776 23000 18806
rect 10317 18730 10383 18733
rect 11697 18730 11763 18733
rect 10317 18728 11763 18730
rect 10317 18672 10322 18728
rect 10378 18672 11702 18728
rect 11758 18672 11763 18728
rect 10317 18670 11763 18672
rect 10317 18667 10383 18670
rect 11697 18667 11763 18670
rect 12525 18730 12591 18733
rect 12893 18730 12959 18733
rect 12525 18728 12959 18730
rect 12525 18672 12530 18728
rect 12586 18672 12898 18728
rect 12954 18672 12959 18728
rect 12525 18670 12959 18672
rect 12525 18667 12591 18670
rect 12893 18667 12959 18670
rect 13629 18730 13695 18733
rect 18781 18730 18847 18733
rect 13629 18728 18847 18730
rect 13629 18672 13634 18728
rect 13690 18672 18786 18728
rect 18842 18672 18847 18728
rect 13629 18670 18847 18672
rect 13629 18667 13695 18670
rect 18781 18667 18847 18670
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 5257 18458 5323 18461
rect 9581 18458 9647 18461
rect 5257 18456 9647 18458
rect 5257 18400 5262 18456
rect 5318 18400 9586 18456
rect 9642 18400 9647 18456
rect 5257 18398 9647 18400
rect 5257 18395 5323 18398
rect 9581 18395 9647 18398
rect 18689 18458 18755 18461
rect 22520 18458 23000 18488
rect 18689 18456 23000 18458
rect 18689 18400 18694 18456
rect 18750 18400 23000 18456
rect 18689 18398 23000 18400
rect 18689 18395 18755 18398
rect 22520 18368 23000 18398
rect 5533 18320 5599 18325
rect 5533 18264 5538 18320
rect 5594 18264 5599 18320
rect 5533 18259 5599 18264
rect 5536 18186 5596 18259
rect 6821 18186 6887 18189
rect 14089 18186 14155 18189
rect 5536 18184 14155 18186
rect 5536 18128 6826 18184
rect 6882 18128 14094 18184
rect 14150 18128 14155 18184
rect 5536 18126 14155 18128
rect 6821 18123 6887 18126
rect 14089 18123 14155 18126
rect 5533 18050 5599 18053
rect 5993 18050 6059 18053
rect 10777 18052 10843 18053
rect 5533 18048 6059 18050
rect 5533 17992 5538 18048
rect 5594 17992 5998 18048
rect 6054 17992 6059 18048
rect 5533 17990 6059 17992
rect 5533 17987 5599 17990
rect 5993 17987 6059 17990
rect 10726 17988 10732 18052
rect 10796 18050 10843 18052
rect 12157 18050 12223 18053
rect 12525 18050 12591 18053
rect 10796 18048 10888 18050
rect 10838 17992 10888 18048
rect 10796 17990 10888 17992
rect 12157 18048 12591 18050
rect 12157 17992 12162 18048
rect 12218 17992 12530 18048
rect 12586 17992 12591 18048
rect 12157 17990 12591 17992
rect 10796 17988 10843 17990
rect 10777 17987 10843 17988
rect 12157 17987 12223 17990
rect 12525 17987 12591 17990
rect 19241 18050 19307 18053
rect 22520 18050 23000 18080
rect 19241 18048 23000 18050
rect 19241 17992 19246 18048
rect 19302 17992 23000 18048
rect 19241 17990 23000 17992
rect 19241 17987 19307 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22520 17960 23000 17990
rect 14805 17919 15125 17920
rect 4061 17914 4127 17917
rect 7005 17914 7071 17917
rect 4061 17912 7071 17914
rect 4061 17856 4066 17912
rect 4122 17856 7010 17912
rect 7066 17856 7071 17912
rect 4061 17854 7071 17856
rect 4061 17851 4127 17854
rect 7005 17851 7071 17854
rect 11053 17778 11119 17781
rect 18597 17778 18663 17781
rect 11053 17776 18663 17778
rect 11053 17720 11058 17776
rect 11114 17720 18602 17776
rect 18658 17720 18663 17776
rect 11053 17718 18663 17720
rect 11053 17715 11119 17718
rect 18597 17715 18663 17718
rect 17861 17642 17927 17645
rect 17861 17640 18890 17642
rect 17861 17584 17866 17640
rect 17922 17584 18890 17640
rect 17861 17582 18890 17584
rect 17861 17579 17927 17582
rect 18830 17506 18890 17582
rect 22520 17506 23000 17536
rect 18830 17446 23000 17506
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22520 17416 23000 17446
rect 18270 17375 18590 17376
rect 0 17234 480 17264
rect 3509 17234 3575 17237
rect 14273 17234 14339 17237
rect 0 17232 3575 17234
rect 0 17176 3514 17232
rect 3570 17176 3575 17232
rect 0 17174 3575 17176
rect 0 17144 480 17174
rect 3509 17171 3575 17174
rect 14046 17232 14339 17234
rect 14046 17176 14278 17232
rect 14334 17176 14339 17232
rect 14046 17174 14339 17176
rect 1761 17098 1827 17101
rect 9121 17098 9187 17101
rect 1761 17096 9187 17098
rect 1761 17040 1766 17096
rect 1822 17040 9126 17096
rect 9182 17040 9187 17096
rect 1761 17038 9187 17040
rect 1761 17035 1827 17038
rect 9121 17035 9187 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 13905 16826 13971 16829
rect 14046 16826 14106 17174
rect 14273 17171 14339 17174
rect 18781 17098 18847 17101
rect 22520 17098 23000 17128
rect 18781 17096 23000 17098
rect 18781 17040 18786 17096
rect 18842 17040 23000 17096
rect 18781 17038 23000 17040
rect 18781 17035 18847 17038
rect 22520 17008 23000 17038
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 13905 16824 14106 16826
rect 13905 16768 13910 16824
rect 13966 16768 14106 16824
rect 13905 16766 14106 16768
rect 13905 16763 13971 16766
rect 10961 16690 11027 16693
rect 11697 16690 11763 16693
rect 10961 16688 11763 16690
rect 10961 16632 10966 16688
rect 11022 16632 11702 16688
rect 11758 16632 11763 16688
rect 10961 16630 11763 16632
rect 10961 16627 11027 16630
rect 11697 16627 11763 16630
rect 17769 16690 17835 16693
rect 17769 16688 17970 16690
rect 17769 16632 17774 16688
rect 17830 16632 17970 16688
rect 17769 16630 17970 16632
rect 17769 16627 17835 16630
rect 17910 16554 17970 16630
rect 22520 16554 23000 16584
rect 17910 16494 23000 16554
rect 22520 16464 23000 16494
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 7097 16146 7163 16149
rect 8845 16146 8911 16149
rect 7097 16144 8911 16146
rect 7097 16088 7102 16144
rect 7158 16088 8850 16144
rect 8906 16088 8911 16144
rect 7097 16086 8911 16088
rect 7097 16083 7163 16086
rect 8845 16083 8911 16086
rect 12341 16146 12407 16149
rect 12985 16146 13051 16149
rect 17401 16146 17467 16149
rect 12341 16144 17467 16146
rect 12341 16088 12346 16144
rect 12402 16088 12990 16144
rect 13046 16088 17406 16144
rect 17462 16088 17467 16144
rect 12341 16086 17467 16088
rect 12341 16083 12407 16086
rect 12985 16083 13051 16086
rect 17401 16083 17467 16086
rect 17861 16146 17927 16149
rect 22520 16146 23000 16176
rect 17861 16144 23000 16146
rect 17861 16088 17866 16144
rect 17922 16088 23000 16144
rect 17861 16086 23000 16088
rect 17861 16083 17927 16086
rect 22520 16056 23000 16086
rect 2589 16010 2655 16013
rect 15837 16010 15903 16013
rect 2589 16008 15903 16010
rect 2589 15952 2594 16008
rect 2650 15952 15842 16008
rect 15898 15952 15903 16008
rect 2589 15950 15903 15952
rect 2589 15947 2655 15950
rect 15837 15947 15903 15950
rect 7557 15876 7623 15877
rect 7557 15872 7604 15876
rect 7668 15874 7674 15876
rect 7557 15816 7562 15872
rect 7557 15812 7604 15816
rect 7668 15814 7714 15874
rect 7668 15812 7674 15814
rect 7557 15811 7623 15812
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 15837 15738 15903 15741
rect 17401 15738 17467 15741
rect 15837 15736 17467 15738
rect 15837 15680 15842 15736
rect 15898 15680 17406 15736
rect 17462 15680 17467 15736
rect 15837 15678 17467 15680
rect 15837 15675 15903 15678
rect 17401 15675 17467 15678
rect 14273 15602 14339 15605
rect 17861 15602 17927 15605
rect 14273 15600 17927 15602
rect 14273 15544 14278 15600
rect 14334 15544 17866 15600
rect 17922 15544 17927 15600
rect 14273 15542 17927 15544
rect 14273 15539 14339 15542
rect 17861 15539 17927 15542
rect 18137 15602 18203 15605
rect 22520 15602 23000 15632
rect 18137 15600 23000 15602
rect 18137 15544 18142 15600
rect 18198 15544 23000 15600
rect 18137 15542 23000 15544
rect 18137 15539 18203 15542
rect 22520 15512 23000 15542
rect 3325 15466 3391 15469
rect 8661 15466 8727 15469
rect 3325 15464 8727 15466
rect 3325 15408 3330 15464
rect 3386 15408 8666 15464
rect 8722 15408 8727 15464
rect 3325 15406 8727 15408
rect 3325 15403 3391 15406
rect 8661 15403 8727 15406
rect 13813 15466 13879 15469
rect 16389 15466 16455 15469
rect 13813 15464 16455 15466
rect 13813 15408 13818 15464
rect 13874 15408 16394 15464
rect 16450 15408 16455 15464
rect 13813 15406 16455 15408
rect 13813 15403 13879 15406
rect 16389 15403 16455 15406
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 22520 15194 23000 15224
rect 18830 15134 23000 15194
rect 1577 15058 1643 15061
rect 9305 15058 9371 15061
rect 1577 15056 9371 15058
rect 1577 15000 1582 15056
rect 1638 15000 9310 15056
rect 9366 15000 9371 15056
rect 1577 14998 9371 15000
rect 1577 14995 1643 14998
rect 9305 14995 9371 14998
rect 11697 15058 11763 15061
rect 11830 15058 11836 15060
rect 11697 15056 11836 15058
rect 11697 15000 11702 15056
rect 11758 15000 11836 15056
rect 11697 14998 11836 15000
rect 11697 14995 11763 14998
rect 11830 14996 11836 14998
rect 11900 15058 11906 15060
rect 16297 15058 16363 15061
rect 11900 15056 16363 15058
rect 11900 15000 16302 15056
rect 16358 15000 16363 15056
rect 11900 14998 16363 15000
rect 11900 14996 11906 14998
rect 16297 14995 16363 14998
rect 18045 15058 18111 15061
rect 18830 15058 18890 15134
rect 22520 15104 23000 15134
rect 18045 15056 18890 15058
rect 18045 15000 18050 15056
rect 18106 15000 18890 15056
rect 18045 14998 18890 15000
rect 18045 14995 18111 14998
rect 5809 14922 5875 14925
rect 8845 14922 8911 14925
rect 13445 14922 13511 14925
rect 5809 14920 13511 14922
rect 5809 14864 5814 14920
rect 5870 14864 8850 14920
rect 8906 14864 13450 14920
rect 13506 14864 13511 14920
rect 5809 14862 13511 14864
rect 5809 14859 5875 14862
rect 8845 14859 8911 14862
rect 13445 14859 13511 14862
rect 8753 14786 8819 14789
rect 13629 14786 13695 14789
rect 8753 14784 13695 14786
rect 8753 14728 8758 14784
rect 8814 14728 13634 14784
rect 13690 14728 13695 14784
rect 8753 14726 13695 14728
rect 8753 14723 8819 14726
rect 13629 14723 13695 14726
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 10041 14650 10107 14653
rect 13813 14650 13879 14653
rect 10041 14648 13879 14650
rect 10041 14592 10046 14648
rect 10102 14592 13818 14648
rect 13874 14592 13879 14648
rect 10041 14590 13879 14592
rect 10041 14587 10107 14590
rect 13813 14587 13879 14590
rect 19885 14650 19951 14653
rect 22520 14650 23000 14680
rect 19885 14648 23000 14650
rect 19885 14592 19890 14648
rect 19946 14592 23000 14648
rect 19885 14590 23000 14592
rect 19885 14587 19951 14590
rect 22520 14560 23000 14590
rect 3417 14514 3483 14517
rect 7741 14514 7807 14517
rect 3417 14512 7807 14514
rect 3417 14456 3422 14512
rect 3478 14456 7746 14512
rect 7802 14456 7807 14512
rect 3417 14454 7807 14456
rect 3417 14451 3483 14454
rect 7741 14451 7807 14454
rect 10225 14514 10291 14517
rect 10501 14514 10567 14517
rect 10225 14512 10567 14514
rect 10225 14456 10230 14512
rect 10286 14456 10506 14512
rect 10562 14456 10567 14512
rect 10225 14454 10567 14456
rect 10225 14451 10291 14454
rect 10501 14451 10567 14454
rect 2865 14378 2931 14381
rect 3693 14378 3759 14381
rect 4797 14378 4863 14381
rect 5717 14378 5783 14381
rect 2865 14376 5783 14378
rect 2865 14320 2870 14376
rect 2926 14320 3698 14376
rect 3754 14320 4802 14376
rect 4858 14320 5722 14376
rect 5778 14320 5783 14376
rect 2865 14318 5783 14320
rect 2865 14315 2931 14318
rect 3693 14315 3759 14318
rect 4797 14315 4863 14318
rect 5717 14315 5783 14318
rect 8477 14378 8543 14381
rect 11697 14378 11763 14381
rect 8477 14376 11763 14378
rect 8477 14320 8482 14376
rect 8538 14320 11702 14376
rect 11758 14320 11763 14376
rect 8477 14318 11763 14320
rect 8477 14315 8543 14318
rect 11697 14315 11763 14318
rect 9673 14242 9739 14245
rect 9990 14242 9996 14244
rect 9673 14240 9996 14242
rect 9673 14184 9678 14240
rect 9734 14184 9996 14240
rect 9673 14182 9996 14184
rect 9673 14179 9739 14182
rect 9990 14180 9996 14182
rect 10060 14180 10066 14244
rect 18781 14242 18847 14245
rect 22520 14242 23000 14272
rect 18781 14240 23000 14242
rect 18781 14184 18786 14240
rect 18842 14184 23000 14240
rect 18781 14182 23000 14184
rect 18781 14179 18847 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22520 14152 23000 14182
rect 18270 14111 18590 14112
rect 9949 14106 10015 14109
rect 10961 14106 11027 14109
rect 9949 14104 11027 14106
rect 9949 14048 9954 14104
rect 10010 14048 10966 14104
rect 11022 14048 11027 14104
rect 9949 14046 11027 14048
rect 9949 14043 10015 14046
rect 10961 14043 11027 14046
rect 1853 13970 1919 13973
rect 8753 13970 8819 13973
rect 1853 13968 8819 13970
rect 1853 13912 1858 13968
rect 1914 13912 8758 13968
rect 8814 13912 8819 13968
rect 1853 13910 8819 13912
rect 1853 13907 1919 13910
rect 8753 13907 8819 13910
rect 8937 13834 9003 13837
rect 11329 13834 11395 13837
rect 12065 13834 12131 13837
rect 16021 13834 16087 13837
rect 8937 13832 16087 13834
rect 8937 13776 8942 13832
rect 8998 13776 11334 13832
rect 11390 13776 12070 13832
rect 12126 13776 16026 13832
rect 16082 13776 16087 13832
rect 8937 13774 16087 13776
rect 8937 13771 9003 13774
rect 11329 13771 11395 13774
rect 12065 13771 12131 13774
rect 16021 13771 16087 13774
rect 18873 13834 18939 13837
rect 22520 13834 23000 13864
rect 18873 13832 23000 13834
rect 18873 13776 18878 13832
rect 18934 13776 23000 13832
rect 18873 13774 23000 13776
rect 18873 13771 18939 13774
rect 22520 13744 23000 13774
rect 8293 13698 8359 13701
rect 9949 13698 10015 13701
rect 8293 13696 10015 13698
rect 8293 13640 8298 13696
rect 8354 13640 9954 13696
rect 10010 13640 10015 13696
rect 8293 13638 10015 13640
rect 8293 13635 8359 13638
rect 9949 13635 10015 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 1393 13562 1459 13565
rect 7465 13562 7531 13565
rect 1393 13560 7531 13562
rect 1393 13504 1398 13560
rect 1454 13504 7470 13560
rect 7526 13504 7531 13560
rect 1393 13502 7531 13504
rect 1393 13499 1459 13502
rect 7465 13499 7531 13502
rect 9029 13562 9095 13565
rect 9397 13562 9463 13565
rect 9029 13560 9463 13562
rect 9029 13504 9034 13560
rect 9090 13504 9402 13560
rect 9458 13504 9463 13560
rect 9029 13502 9463 13504
rect 9029 13499 9095 13502
rect 9397 13499 9463 13502
rect 9622 13500 9628 13564
rect 9692 13562 9698 13564
rect 9765 13562 9831 13565
rect 9692 13560 9831 13562
rect 9692 13504 9770 13560
rect 9826 13504 9831 13560
rect 9692 13502 9831 13504
rect 9692 13500 9698 13502
rect 9765 13499 9831 13502
rect 10317 13562 10383 13565
rect 10317 13560 12404 13562
rect 10317 13504 10322 13560
rect 10378 13504 12404 13560
rect 10317 13502 12404 13504
rect 10317 13499 10383 13502
rect 12157 13426 12223 13429
rect 9998 13424 12223 13426
rect 9998 13368 12162 13424
rect 12218 13368 12223 13424
rect 9998 13366 12223 13368
rect 12344 13426 12404 13502
rect 19241 13426 19307 13429
rect 12344 13424 19307 13426
rect 12344 13368 19246 13424
rect 19302 13368 19307 13424
rect 12344 13366 19307 13368
rect 9998 13293 10058 13366
rect 12157 13363 12223 13366
rect 19241 13363 19307 13366
rect 9949 13288 10058 13293
rect 9949 13232 9954 13288
rect 10010 13232 10058 13288
rect 9949 13230 10058 13232
rect 12157 13290 12223 13293
rect 13353 13290 13419 13293
rect 16573 13290 16639 13293
rect 12157 13288 16639 13290
rect 12157 13232 12162 13288
rect 12218 13232 13358 13288
rect 13414 13232 16578 13288
rect 16634 13232 16639 13288
rect 12157 13230 16639 13232
rect 9949 13227 10015 13230
rect 12157 13227 12223 13230
rect 13353 13227 13419 13230
rect 16573 13227 16639 13230
rect 18597 13290 18663 13293
rect 22520 13290 23000 13320
rect 18597 13288 23000 13290
rect 18597 13232 18602 13288
rect 18658 13232 23000 13288
rect 18597 13230 23000 13232
rect 18597 13227 18663 13230
rect 22520 13200 23000 13230
rect 8753 13154 8819 13157
rect 10317 13154 10383 13157
rect 8753 13152 10383 13154
rect 8753 13096 8758 13152
rect 8814 13096 10322 13152
rect 10378 13096 10383 13152
rect 8753 13094 10383 13096
rect 8753 13091 8819 13094
rect 10317 13091 10383 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 7557 13020 7623 13021
rect 7557 13018 7604 13020
rect 7512 13016 7604 13018
rect 7512 12960 7562 13016
rect 7512 12958 7604 12960
rect 7557 12956 7604 12958
rect 7668 12956 7674 13020
rect 9857 13018 9923 13021
rect 9990 13018 9996 13020
rect 9857 13016 9996 13018
rect 9857 12960 9862 13016
rect 9918 12960 9996 13016
rect 9857 12958 9996 12960
rect 7557 12955 7623 12956
rect 9857 12955 9923 12958
rect 9990 12956 9996 12958
rect 10060 12956 10066 13020
rect 14641 13018 14707 13021
rect 14641 13016 17050 13018
rect 14641 12960 14646 13016
rect 14702 12960 17050 13016
rect 14641 12958 17050 12960
rect 14641 12955 14707 12958
rect 6361 12882 6427 12885
rect 7097 12882 7163 12885
rect 6361 12880 7163 12882
rect 6361 12824 6366 12880
rect 6422 12824 7102 12880
rect 7158 12824 7163 12880
rect 6361 12822 7163 12824
rect 6361 12819 6427 12822
rect 7097 12819 7163 12822
rect 9622 12820 9628 12884
rect 9692 12882 9698 12884
rect 9765 12882 9831 12885
rect 9692 12880 9831 12882
rect 9692 12824 9770 12880
rect 9826 12824 9831 12880
rect 9692 12822 9831 12824
rect 9692 12820 9698 12822
rect 9765 12819 9831 12822
rect 11697 12882 11763 12885
rect 16757 12882 16823 12885
rect 11697 12880 16823 12882
rect 11697 12824 11702 12880
rect 11758 12824 16762 12880
rect 16818 12824 16823 12880
rect 11697 12822 16823 12824
rect 16990 12882 17050 12958
rect 22520 12882 23000 12912
rect 16990 12822 23000 12882
rect 11697 12819 11763 12822
rect 16757 12819 16823 12822
rect 22520 12792 23000 12822
rect 12433 12746 12499 12749
rect 18965 12746 19031 12749
rect 12433 12744 19031 12746
rect 12433 12688 12438 12744
rect 12494 12688 18970 12744
rect 19026 12688 19031 12744
rect 12433 12686 19031 12688
rect 12433 12683 12499 12686
rect 18965 12683 19031 12686
rect 8661 12610 8727 12613
rect 11973 12610 12039 12613
rect 8661 12608 12039 12610
rect 8661 12552 8666 12608
rect 8722 12552 11978 12608
rect 12034 12552 12039 12608
rect 8661 12550 12039 12552
rect 8661 12547 8727 12550
rect 11973 12547 12039 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 9121 12474 9187 12477
rect 12525 12474 12591 12477
rect 9121 12472 12591 12474
rect 9121 12416 9126 12472
rect 9182 12416 12530 12472
rect 12586 12416 12591 12472
rect 9121 12414 12591 12416
rect 9121 12411 9187 12414
rect 12525 12411 12591 12414
rect 6177 12338 6243 12341
rect 19793 12338 19859 12341
rect 22520 12338 23000 12368
rect 6177 12336 19859 12338
rect 6177 12280 6182 12336
rect 6238 12280 19798 12336
rect 19854 12280 19859 12336
rect 6177 12278 19859 12280
rect 6177 12275 6243 12278
rect 19793 12275 19859 12278
rect 21038 12278 23000 12338
rect 3049 12202 3115 12205
rect 20805 12202 20871 12205
rect 3049 12200 20871 12202
rect 3049 12144 3054 12200
rect 3110 12144 20810 12200
rect 20866 12144 20871 12200
rect 3049 12142 20871 12144
rect 3049 12139 3115 12142
rect 20805 12139 20871 12142
rect 8477 12066 8543 12069
rect 9673 12066 9739 12069
rect 10409 12066 10475 12069
rect 11789 12068 11855 12069
rect 11789 12066 11836 12068
rect 8477 12064 10475 12066
rect 8477 12008 8482 12064
rect 8538 12008 9678 12064
rect 9734 12008 10414 12064
rect 10470 12008 10475 12064
rect 8477 12006 10475 12008
rect 11744 12064 11836 12066
rect 11744 12008 11794 12064
rect 11744 12006 11836 12008
rect 8477 12003 8543 12006
rect 9673 12003 9739 12006
rect 10409 12003 10475 12006
rect 11789 12004 11836 12006
rect 11900 12004 11906 12068
rect 18689 12066 18755 12069
rect 21038 12066 21098 12278
rect 22520 12248 23000 12278
rect 18689 12064 21098 12066
rect 18689 12008 18694 12064
rect 18750 12008 21098 12064
rect 18689 12006 21098 12008
rect 11789 12003 11855 12004
rect 18689 12003 18755 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 11973 11930 12039 11933
rect 15745 11930 15811 11933
rect 22520 11930 23000 11960
rect 11973 11928 15811 11930
rect 11973 11872 11978 11928
rect 12034 11872 15750 11928
rect 15806 11872 15811 11928
rect 11973 11870 15811 11872
rect 11973 11867 12039 11870
rect 15745 11867 15811 11870
rect 21038 11870 23000 11930
rect 4429 11794 4495 11797
rect 20897 11794 20963 11797
rect 4429 11792 20963 11794
rect 4429 11736 4434 11792
rect 4490 11736 20902 11792
rect 20958 11736 20963 11792
rect 4429 11734 20963 11736
rect 4429 11731 4495 11734
rect 20897 11731 20963 11734
rect 1393 11658 1459 11661
rect 18321 11658 18387 11661
rect 1393 11656 18387 11658
rect 1393 11600 1398 11656
rect 1454 11600 18326 11656
rect 18382 11600 18387 11656
rect 1393 11598 18387 11600
rect 1393 11595 1459 11598
rect 18321 11595 18387 11598
rect 8385 11522 8451 11525
rect 9397 11522 9463 11525
rect 8385 11520 9463 11522
rect 8385 11464 8390 11520
rect 8446 11464 9402 11520
rect 9458 11464 9463 11520
rect 8385 11462 9463 11464
rect 8385 11459 8451 11462
rect 9397 11459 9463 11462
rect 10041 11522 10107 11525
rect 11973 11522 12039 11525
rect 10041 11520 12039 11522
rect 10041 11464 10046 11520
rect 10102 11464 11978 11520
rect 12034 11464 12039 11520
rect 10041 11462 12039 11464
rect 10041 11459 10107 11462
rect 11973 11459 12039 11462
rect 15653 11522 15719 11525
rect 21038 11522 21098 11870
rect 22520 11840 23000 11870
rect 15653 11520 21098 11522
rect 15653 11464 15658 11520
rect 15714 11464 21098 11520
rect 15653 11462 21098 11464
rect 15653 11459 15719 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9121 11386 9187 11389
rect 11973 11386 12039 11389
rect 9121 11384 12039 11386
rect 9121 11328 9126 11384
rect 9182 11328 11978 11384
rect 12034 11328 12039 11384
rect 9121 11326 12039 11328
rect 9121 11323 9187 11326
rect 11973 11323 12039 11326
rect 15377 11386 15443 11389
rect 22520 11386 23000 11416
rect 15377 11384 23000 11386
rect 15377 11328 15382 11384
rect 15438 11328 23000 11384
rect 15377 11326 23000 11328
rect 15377 11323 15443 11326
rect 22520 11296 23000 11326
rect 7925 11250 7991 11253
rect 8753 11250 8819 11253
rect 12525 11250 12591 11253
rect 7925 11248 12591 11250
rect 7925 11192 7930 11248
rect 7986 11192 8758 11248
rect 8814 11192 12530 11248
rect 12586 11192 12591 11248
rect 7925 11190 12591 11192
rect 7925 11187 7991 11190
rect 8753 11187 8819 11190
rect 12525 11187 12591 11190
rect 15285 11250 15351 11253
rect 17953 11250 18019 11253
rect 15285 11248 18019 11250
rect 15285 11192 15290 11248
rect 15346 11192 17958 11248
rect 18014 11192 18019 11248
rect 15285 11190 18019 11192
rect 15285 11187 15351 11190
rect 17953 11187 18019 11190
rect 5441 11114 5507 11117
rect 10685 11114 10751 11117
rect 16757 11114 16823 11117
rect 5441 11112 10751 11114
rect 5441 11056 5446 11112
rect 5502 11056 10690 11112
rect 10746 11056 10751 11112
rect 5441 11054 10751 11056
rect 5441 11051 5507 11054
rect 10685 11051 10751 11054
rect 11148 11054 16682 11114
rect 4797 10978 4863 10981
rect 11148 10978 11208 11054
rect 4797 10976 11208 10978
rect 4797 10920 4802 10976
rect 4858 10920 11208 10976
rect 4797 10918 11208 10920
rect 16622 10978 16682 11054
rect 16757 11112 18890 11114
rect 16757 11056 16762 11112
rect 16818 11056 18890 11112
rect 16757 11054 18890 11056
rect 16757 11051 16823 11054
rect 17677 10978 17743 10981
rect 16622 10976 17743 10978
rect 16622 10920 17682 10976
rect 17738 10920 17743 10976
rect 16622 10918 17743 10920
rect 18830 10978 18890 11054
rect 19241 10978 19307 10981
rect 22520 10978 23000 11008
rect 18830 10976 23000 10978
rect 18830 10920 19246 10976
rect 19302 10920 23000 10976
rect 18830 10918 23000 10920
rect 4797 10915 4863 10918
rect 17677 10915 17743 10918
rect 19241 10915 19307 10918
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 22520 10888 23000 10918
rect 18270 10847 18590 10848
rect 8477 10842 8543 10845
rect 10317 10842 10383 10845
rect 8477 10840 10383 10842
rect 8477 10784 8482 10840
rect 8538 10784 10322 10840
rect 10378 10784 10383 10840
rect 8477 10782 10383 10784
rect 8477 10779 8543 10782
rect 10317 10779 10383 10782
rect 5809 10706 5875 10709
rect 5809 10704 15578 10706
rect 5809 10648 5814 10704
rect 5870 10648 15578 10704
rect 5809 10646 15578 10648
rect 5809 10643 5875 10646
rect 4613 10570 4679 10573
rect 15518 10570 15578 10646
rect 20069 10570 20135 10573
rect 4613 10568 15394 10570
rect 4613 10512 4618 10568
rect 4674 10512 15394 10568
rect 4613 10510 15394 10512
rect 15518 10568 20135 10570
rect 15518 10512 20074 10568
rect 20130 10512 20135 10568
rect 15518 10510 20135 10512
rect 4613 10507 4679 10510
rect 10685 10434 10751 10437
rect 12433 10434 12499 10437
rect 10685 10432 12499 10434
rect 10685 10376 10690 10432
rect 10746 10376 12438 10432
rect 12494 10376 12499 10432
rect 10685 10374 12499 10376
rect 15334 10434 15394 10510
rect 20069 10507 20135 10510
rect 20253 10434 20319 10437
rect 15334 10432 20319 10434
rect 15334 10376 20258 10432
rect 20314 10376 20319 10432
rect 15334 10374 20319 10376
rect 10685 10371 10751 10374
rect 12433 10371 12499 10374
rect 20253 10371 20319 10374
rect 20529 10434 20595 10437
rect 22520 10434 23000 10464
rect 20529 10432 23000 10434
rect 20529 10376 20534 10432
rect 20590 10376 23000 10432
rect 20529 10374 23000 10376
rect 20529 10371 20595 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22520 10344 23000 10374
rect 14805 10303 15125 10304
rect 10041 10298 10107 10301
rect 11789 10298 11855 10301
rect 10041 10296 11855 10298
rect 10041 10240 10046 10296
rect 10102 10240 11794 10296
rect 11850 10240 11855 10296
rect 10041 10238 11855 10240
rect 10041 10235 10107 10238
rect 11789 10235 11855 10238
rect 6821 10162 6887 10165
rect 20989 10162 21055 10165
rect 6821 10160 21055 10162
rect 6821 10104 6826 10160
rect 6882 10104 20994 10160
rect 21050 10104 21055 10160
rect 6821 10102 21055 10104
rect 6821 10099 6887 10102
rect 20989 10099 21055 10102
rect 1669 10026 1735 10029
rect 17677 10026 17743 10029
rect 22520 10026 23000 10056
rect 1669 10024 17743 10026
rect 1669 9968 1674 10024
rect 1730 9968 17682 10024
rect 17738 9968 17743 10024
rect 1669 9966 17743 9968
rect 1669 9963 1735 9966
rect 17677 9963 17743 9966
rect 18094 9966 23000 10026
rect 12157 9890 12223 9893
rect 17125 9890 17191 9893
rect 12157 9888 17191 9890
rect 12157 9832 12162 9888
rect 12218 9832 17130 9888
rect 17186 9832 17191 9888
rect 12157 9830 17191 9832
rect 12157 9827 12223 9830
rect 17125 9827 17191 9830
rect 17769 9890 17835 9893
rect 18094 9890 18154 9966
rect 22520 9936 23000 9966
rect 17769 9888 18154 9890
rect 17769 9832 17774 9888
rect 17830 9832 18154 9888
rect 17769 9830 18154 9832
rect 17769 9827 17835 9830
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 7097 9754 7163 9757
rect 20345 9754 20411 9757
rect 7097 9752 11208 9754
rect 7097 9696 7102 9752
rect 7158 9696 11208 9752
rect 7097 9694 11208 9696
rect 7097 9691 7163 9694
rect 3601 9618 3667 9621
rect 7281 9618 7347 9621
rect 8201 9618 8267 9621
rect 3601 9616 8267 9618
rect 3601 9560 3606 9616
rect 3662 9560 7286 9616
rect 7342 9560 8206 9616
rect 8262 9560 8267 9616
rect 3601 9558 8267 9560
rect 11148 9618 11208 9694
rect 11792 9694 18154 9754
rect 11792 9618 11852 9694
rect 11148 9558 11852 9618
rect 11973 9618 12039 9621
rect 12525 9618 12591 9621
rect 11973 9616 12591 9618
rect 11973 9560 11978 9616
rect 12034 9560 12530 9616
rect 12586 9560 12591 9616
rect 11973 9558 12591 9560
rect 18094 9618 18154 9694
rect 18830 9752 20411 9754
rect 18830 9696 20350 9752
rect 20406 9696 20411 9752
rect 18830 9694 20411 9696
rect 18830 9618 18890 9694
rect 20345 9691 20411 9694
rect 18094 9558 18890 9618
rect 3601 9555 3667 9558
rect 7281 9555 7347 9558
rect 8201 9555 8267 9558
rect 11973 9555 12039 9558
rect 12525 9555 12591 9558
rect 4797 9482 4863 9485
rect 9213 9482 9279 9485
rect 4797 9480 9279 9482
rect 4797 9424 4802 9480
rect 4858 9424 9218 9480
rect 9274 9424 9279 9480
rect 4797 9422 9279 9424
rect 4797 9419 4863 9422
rect 9213 9419 9279 9422
rect 13537 9482 13603 9485
rect 15653 9482 15719 9485
rect 13537 9480 15719 9482
rect 13537 9424 13542 9480
rect 13598 9424 15658 9480
rect 15714 9424 15719 9480
rect 13537 9422 15719 9424
rect 13537 9419 13603 9422
rect 15653 9419 15719 9422
rect 18137 9482 18203 9485
rect 22520 9482 23000 9512
rect 18137 9480 23000 9482
rect 18137 9424 18142 9480
rect 18198 9424 23000 9480
rect 18137 9422 23000 9424
rect 18137 9419 18203 9422
rect 22520 9392 23000 9422
rect 8293 9346 8359 9349
rect 9581 9346 9647 9349
rect 8293 9344 9647 9346
rect 8293 9288 8298 9344
rect 8354 9288 9586 9344
rect 9642 9288 9647 9344
rect 8293 9286 9647 9288
rect 8293 9283 8359 9286
rect 9581 9283 9647 9286
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 17953 9074 18019 9077
rect 22520 9074 23000 9104
rect 17953 9072 23000 9074
rect 17953 9016 17958 9072
rect 18014 9016 23000 9072
rect 17953 9014 23000 9016
rect 17953 9011 18019 9014
rect 22520 8984 23000 9014
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 22520 8666 23000 8696
rect 18692 8606 23000 8666
rect 14733 8530 14799 8533
rect 18692 8530 18752 8606
rect 22520 8576 23000 8606
rect 14733 8528 18752 8530
rect 14733 8472 14738 8528
rect 14794 8472 18752 8528
rect 14733 8470 18752 8472
rect 14733 8467 14799 8470
rect 4429 8394 4495 8397
rect 19885 8394 19951 8397
rect 4429 8392 19951 8394
rect 4429 8336 4434 8392
rect 4490 8336 19890 8392
rect 19946 8336 19951 8392
rect 4429 8334 19951 8336
rect 4429 8331 4495 8334
rect 19885 8331 19951 8334
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 18321 8122 18387 8125
rect 22520 8122 23000 8152
rect 18321 8120 23000 8122
rect 18321 8064 18326 8120
rect 18382 8064 23000 8120
rect 18321 8062 23000 8064
rect 18321 8059 18387 8062
rect 22520 8032 23000 8062
rect 17677 7986 17743 7989
rect 18045 7986 18111 7989
rect 17677 7984 18111 7986
rect 17677 7928 17682 7984
rect 17738 7928 18050 7984
rect 18106 7928 18111 7984
rect 17677 7926 18111 7928
rect 17677 7923 17743 7926
rect 18045 7923 18111 7926
rect 18689 7714 18755 7717
rect 22520 7714 23000 7744
rect 18689 7712 23000 7714
rect 18689 7656 18694 7712
rect 18750 7656 23000 7712
rect 18689 7654 23000 7656
rect 18689 7651 18755 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22520 7624 23000 7654
rect 18270 7583 18590 7584
rect 18873 7170 18939 7173
rect 22520 7170 23000 7200
rect 18873 7168 23000 7170
rect 18873 7112 18878 7168
rect 18934 7112 23000 7168
rect 18873 7110 23000 7112
rect 18873 7107 18939 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22520 7080 23000 7110
rect 14805 7039 15125 7040
rect 3969 6898 4035 6901
rect 8477 6898 8543 6901
rect 3969 6896 8543 6898
rect 3969 6840 3974 6896
rect 4030 6840 8482 6896
rect 8538 6840 8543 6896
rect 3969 6838 8543 6840
rect 3969 6835 4035 6838
rect 8477 6835 8543 6838
rect 19241 6762 19307 6765
rect 22520 6762 23000 6792
rect 19241 6760 23000 6762
rect 19241 6704 19246 6760
rect 19302 6704 23000 6760
rect 19241 6702 23000 6704
rect 19241 6699 19307 6702
rect 22520 6672 23000 6702
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 18597 6218 18663 6221
rect 22520 6218 23000 6248
rect 18597 6216 23000 6218
rect 18597 6160 18602 6216
rect 18658 6160 23000 6216
rect 18597 6158 23000 6160
rect 18597 6155 18663 6158
rect 22520 6128 23000 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5810 480 5840
rect 3049 5810 3115 5813
rect 0 5808 3115 5810
rect 0 5752 3054 5808
rect 3110 5752 3115 5808
rect 0 5750 3115 5752
rect 0 5720 480 5750
rect 3049 5747 3115 5750
rect 17861 5810 17927 5813
rect 22520 5810 23000 5840
rect 17861 5808 23000 5810
rect 17861 5752 17866 5808
rect 17922 5752 23000 5808
rect 17861 5750 23000 5752
rect 17861 5747 17927 5750
rect 22520 5720 23000 5750
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 18045 5266 18111 5269
rect 22520 5266 23000 5296
rect 18045 5264 23000 5266
rect 18045 5208 18050 5264
rect 18106 5208 23000 5264
rect 18045 5206 23000 5208
rect 18045 5203 18111 5206
rect 22520 5176 23000 5206
rect 6913 5130 6979 5133
rect 7373 5130 7439 5133
rect 18873 5130 18939 5133
rect 6913 5128 18939 5130
rect 6913 5072 6918 5128
rect 6974 5072 7378 5128
rect 7434 5072 18878 5128
rect 18934 5072 18939 5128
rect 6913 5070 18939 5072
rect 6913 5067 6979 5070
rect 7373 5067 7439 5070
rect 18873 5067 18939 5070
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 18045 4858 18111 4861
rect 22520 4858 23000 4888
rect 18045 4856 23000 4858
rect 18045 4800 18050 4856
rect 18106 4800 23000 4856
rect 18045 4798 23000 4800
rect 18045 4795 18111 4798
rect 22520 4768 23000 4798
rect 10777 4722 10843 4725
rect 15745 4722 15811 4725
rect 10777 4720 15811 4722
rect 10777 4664 10782 4720
rect 10838 4664 15750 4720
rect 15806 4664 15811 4720
rect 10777 4662 15811 4664
rect 10777 4659 10843 4662
rect 15745 4659 15811 4662
rect 17677 4586 17743 4589
rect 17677 4584 18890 4586
rect 17677 4528 17682 4584
rect 17738 4528 18890 4584
rect 17677 4526 18890 4528
rect 17677 4523 17743 4526
rect 18830 4450 18890 4526
rect 22520 4450 23000 4480
rect 18830 4390 23000 4450
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22520 4360 23000 4390
rect 18270 4319 18590 4320
rect 6821 4178 6887 4181
rect 10317 4178 10383 4181
rect 6821 4176 10383 4178
rect 6821 4120 6826 4176
rect 6882 4120 10322 4176
rect 10378 4120 10383 4176
rect 6821 4118 10383 4120
rect 6821 4115 6887 4118
rect 10317 4115 10383 4118
rect 5165 4042 5231 4045
rect 6085 4042 6151 4045
rect 5165 4040 6151 4042
rect 5165 3984 5170 4040
rect 5226 3984 6090 4040
rect 6146 3984 6151 4040
rect 5165 3982 6151 3984
rect 5165 3979 5231 3982
rect 6085 3979 6151 3982
rect 6637 4042 6703 4045
rect 10685 4042 10751 4045
rect 6637 4040 10751 4042
rect 6637 3984 6642 4040
rect 6698 3984 10690 4040
rect 10746 3984 10751 4040
rect 6637 3982 10751 3984
rect 6637 3979 6703 3982
rect 10685 3979 10751 3982
rect 9765 3906 9831 3909
rect 14641 3906 14707 3909
rect 9765 3904 14707 3906
rect 9765 3848 9770 3904
rect 9826 3848 14646 3904
rect 14702 3848 14707 3904
rect 9765 3846 14707 3848
rect 9765 3843 9831 3846
rect 14641 3843 14707 3846
rect 19977 3906 20043 3909
rect 22520 3906 23000 3936
rect 19977 3904 23000 3906
rect 19977 3848 19982 3904
rect 20038 3848 23000 3904
rect 19977 3846 23000 3848
rect 19977 3843 20043 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22520 3816 23000 3846
rect 14805 3775 15125 3776
rect 3049 3770 3115 3773
rect 7741 3770 7807 3773
rect 3049 3768 7807 3770
rect 3049 3712 3054 3768
rect 3110 3712 7746 3768
rect 7802 3712 7807 3768
rect 3049 3710 7807 3712
rect 3049 3707 3115 3710
rect 7741 3707 7807 3710
rect 2865 3498 2931 3501
rect 12065 3498 12131 3501
rect 2865 3496 12131 3498
rect 2865 3440 2870 3496
rect 2926 3440 12070 3496
rect 12126 3440 12131 3496
rect 2865 3438 12131 3440
rect 2865 3435 2931 3438
rect 12065 3435 12131 3438
rect 18689 3498 18755 3501
rect 22520 3498 23000 3528
rect 18689 3496 23000 3498
rect 18689 3440 18694 3496
rect 18750 3440 23000 3496
rect 18689 3438 23000 3440
rect 18689 3435 18755 3438
rect 22520 3408 23000 3438
rect 4797 3362 4863 3365
rect 8293 3362 8359 3365
rect 4797 3360 8359 3362
rect 4797 3304 4802 3360
rect 4858 3304 8298 3360
rect 8354 3304 8359 3360
rect 4797 3302 8359 3304
rect 4797 3299 4863 3302
rect 8293 3299 8359 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 6913 3226 6979 3229
rect 7557 3226 7623 3229
rect 8109 3226 8175 3229
rect 6913 3224 8175 3226
rect 6913 3168 6918 3224
rect 6974 3168 7562 3224
rect 7618 3168 8114 3224
rect 8170 3168 8175 3224
rect 6913 3166 8175 3168
rect 6913 3163 6979 3166
rect 7557 3163 7623 3166
rect 8109 3163 8175 3166
rect 2037 3090 2103 3093
rect 8293 3090 8359 3093
rect 2037 3088 8359 3090
rect 2037 3032 2042 3088
rect 2098 3032 8298 3088
rect 8354 3032 8359 3088
rect 2037 3030 8359 3032
rect 2037 3027 2103 3030
rect 8293 3027 8359 3030
rect 14365 3090 14431 3093
rect 14825 3090 14891 3093
rect 14365 3088 14891 3090
rect 14365 3032 14370 3088
rect 14426 3032 14830 3088
rect 14886 3032 14891 3088
rect 14365 3030 14891 3032
rect 14365 3027 14431 3030
rect 14825 3027 14891 3030
rect 7373 2954 7439 2957
rect 7741 2954 7807 2957
rect 7373 2952 7807 2954
rect 7373 2896 7378 2952
rect 7434 2896 7746 2952
rect 7802 2896 7807 2952
rect 7373 2894 7807 2896
rect 7373 2891 7439 2894
rect 7741 2891 7807 2894
rect 19149 2954 19215 2957
rect 22520 2954 23000 2984
rect 19149 2952 23000 2954
rect 19149 2896 19154 2952
rect 19210 2896 23000 2952
rect 19149 2894 23000 2896
rect 19149 2891 19215 2894
rect 22520 2864 23000 2894
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 18873 2546 18939 2549
rect 22520 2546 23000 2576
rect 18873 2544 23000 2546
rect 18873 2488 18878 2544
rect 18934 2488 23000 2544
rect 18873 2486 23000 2488
rect 18873 2483 18939 2486
rect 22520 2456 23000 2486
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 19057 2002 19123 2005
rect 22520 2002 23000 2032
rect 19057 2000 23000 2002
rect 19057 1944 19062 2000
rect 19118 1944 23000 2000
rect 19057 1942 23000 1944
rect 19057 1939 19123 1942
rect 22520 1912 23000 1942
rect 17953 1594 18019 1597
rect 22520 1594 23000 1624
rect 17953 1592 23000 1594
rect 17953 1536 17958 1592
rect 18014 1536 23000 1592
rect 17953 1534 23000 1536
rect 17953 1531 18019 1534
rect 22520 1504 23000 1534
rect 17953 1050 18019 1053
rect 22520 1050 23000 1080
rect 17953 1048 23000 1050
rect 17953 992 17958 1048
rect 18014 992 23000 1048
rect 17953 990 23000 992
rect 17953 987 18019 990
rect 22520 960 23000 990
rect 18045 642 18111 645
rect 22520 642 23000 672
rect 18045 640 23000 642
rect 18045 584 18050 640
rect 18106 584 23000 640
rect 18045 582 23000 584
rect 18045 579 18111 582
rect 22520 552 23000 582
rect 18137 234 18203 237
rect 22520 234 23000 264
rect 18137 232 23000 234
rect 18137 176 18142 232
rect 18198 176 23000 232
rect 18137 174 23000 176
rect 18137 171 18203 174
rect 22520 144 23000 174
<< via3 >>
rect 10732 22536 10796 22540
rect 10732 22480 10782 22536
rect 10782 22480 10796 22536
rect 10732 22476 10796 22480
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 10732 18048 10796 18052
rect 10732 17992 10782 18048
rect 10782 17992 10796 18048
rect 10732 17988 10796 17992
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7604 15872 7668 15876
rect 7604 15816 7618 15872
rect 7618 15816 7668 15872
rect 7604 15812 7668 15816
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 11836 14996 11900 15060
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 9996 14180 10060 14244
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 9628 13500 9692 13564
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7604 13016 7668 13020
rect 7604 12960 7618 13016
rect 7618 12960 7668 13016
rect 7604 12956 7668 12960
rect 9996 12956 10060 13020
rect 9628 12820 9692 12884
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 11836 12064 11900 12068
rect 11836 12008 11850 12064
rect 11850 12008 11900 12064
rect 11836 12004 11900 12008
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 10731 22540 10797 22541
rect 10731 22476 10732 22540
rect 10796 22476 10797 22540
rect 10731 22475 10797 22476
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 10734 18053 10794 22475
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 10731 18052 10797 18053
rect 10731 17988 10732 18052
rect 10796 17988 10797 18052
rect 10731 17987 10797 17988
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7603 15876 7669 15877
rect 7603 15812 7604 15876
rect 7668 15812 7669 15876
rect 7603 15811 7669 15812
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 7606 13021 7666 15811
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 9995 14244 10061 14245
rect 9995 14180 9996 14244
rect 10060 14180 10061 14244
rect 9995 14179 10061 14180
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7603 13020 7669 13021
rect 7603 12956 7604 13020
rect 7668 12956 7669 13020
rect 7603 12955 7669 12956
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 12544 8195 13568
rect 9627 13564 9693 13565
rect 9627 13500 9628 13564
rect 9692 13500 9693 13564
rect 9627 13499 9693 13500
rect 9630 12885 9690 13499
rect 9998 13021 10058 14179
rect 11340 14176 11660 15200
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 11835 15060 11901 15061
rect 11835 14996 11836 15060
rect 11900 14996 11901 15060
rect 11835 14995 11901 14996
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 9995 13020 10061 13021
rect 9995 12956 9996 13020
rect 10060 12956 10061 13020
rect 9995 12955 10061 12956
rect 9627 12884 9693 12885
rect 9627 12820 9628 12884
rect 9692 12820 9693 12884
rect 9627 12819 9693 12820
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 12000 11660 13024
rect 11838 12069 11898 14995
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 11835 12068 11901 12069
rect 11835 12004 11836 12068
rect 11900 12004 11901 12068
rect 11835 12003 11901 12004
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _038_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_12 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 2944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4048 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_24
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_50 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_48
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 1604681595
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_78
timestamp 1604681595
transform 1 0 8280 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1604681595
transform 1 0 10580 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1604681595
transform 1 0 11316 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12696 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_131
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_132
timestamp 1604681595
transform 1 0 13248 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_166
timestamp 1604681595
transform 1 0 16376 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1604681595
transform 1 0 15824 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_168
timestamp 1604681595
transform 1 0 16560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_175
timestamp 1604681595
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18952 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_193
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_200
timestamp 1604681595
transform 1 0 19504 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_193
timestamp 1604681595
transform 1 0 18860 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1604681595
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1604681595
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_210
timestamp 1604681595
transform 1 0 20424 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1604681595
transform 1 0 21528 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_2_52
timestamp 1604681595
transform 1 0 5888 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_60
timestamp 1604681595
transform 1 0 6624 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_109
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1604681595
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1604681595
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_158
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17940 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 17756 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_175
timestamp 1604681595
transform 1 0 17204 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_192
timestamp 1604681595
transform 1 0 18768 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_10
timestamp 1604681595
transform 1 0 2024 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_42
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_53
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8556 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_73
timestamp 1604681595
transform 1 0 7820 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_97
timestamp 1604681595
transform 1 0 10028 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 10764 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_139
timestamp 1604681595
transform 1 0 13892 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_156
timestamp 1604681595
transform 1 0 15456 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_164
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_3_191
timestamp 1604681595
transform 1 0 18676 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_50
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_67
timestamp 1604681595
transform 1 0 7268 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 9752 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_84
timestamp 1604681595
transform 1 0 8832 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_98
timestamp 1604681595
transform 1 0 10120 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_4_122
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1604681595
transform 1 0 13432 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_163
timestamp 1604681595
transform 1 0 16100 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_171
timestamp 1604681595
transform 1 0 16836 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_181
timestamp 1604681595
transform 1 0 17756 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18492 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_205
timestamp 1604681595
transform 1 0 19964 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_14
timestamp 1604681595
transform 1 0 2392 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3128 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_38
timestamp 1604681595
transform 1 0 4600 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_46
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1604681595
transform 1 0 5980 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7360 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 9660 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_84
timestamp 1604681595
transform 1 0 8832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_92
timestamp 1604681595
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_97
timestamp 1604681595
transform 1 0 10028 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13708 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_129
timestamp 1604681595
transform 1 0 12972 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_146
timestamp 1604681595
transform 1 0 14536 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1604681595
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 18308 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_191
timestamp 1604681595
transform 1 0 18676 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_12
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1604681595
transform 1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3772 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_21
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 1604681595
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_72
timestamp 1604681595
transform 1 0 7728 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_84
timestamp 1604681595
transform 1 0 8832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 1604681595
transform 1 0 11132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1604681595
transform 1 0 10764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604681595
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_6_126
timestamp 1604681595
transform 1 0 12696 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_143
timestamp 1604681595
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_132
timestamp 1604681595
transform 1 0 13248 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_145
timestamp 1604681595
transform 1 0 14444 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 15640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15180 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_162
timestamp 1604681595
transform 1 0 16008 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16744 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1604681595
transform 1 0 18216 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1604681595
transform 1 0 16652 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19688 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_194
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_194
timestamp 1604681595
transform 1 0 18952 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_211
timestamp 1604681595
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_40
timestamp 1604681595
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 4968 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5980 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_45
timestamp 1604681595
transform 1 0 5244 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1604681595
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12052 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_111
timestamp 1604681595
transform 1 0 11316 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_128
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 17664 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_170
timestamp 1604681595
transform 1 0 16744 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1604681595
transform 1 0 19136 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_208
timestamp 1604681595
transform 1 0 20240 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_19
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1604681595
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_96
timestamp 1604681595
transform 1 0 9936 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_113
timestamp 1604681595
transform 1 0 11500 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604681595
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1604681595
transform 1 0 14812 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_166
timestamp 1604681595
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604681595
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_200
timestamp 1604681595
transform 1 0 19504 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1604681595
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_39
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7636 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_63
timestamp 1604681595
transform 1 0 6900 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9752 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 11960 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_110
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13524 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_10_127
timestamp 1604681595
transform 1 0 12788 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1604681595
transform 1 0 14352 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17204 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_174
timestamp 1604681595
transform 1 0 17112 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_184
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1604681595
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_42
timestamp 1604681595
transform 1 0 4968 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_53
timestamp 1604681595
transform 1 0 5980 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_83
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9476 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_100
timestamp 1604681595
transform 1 0 10304 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1604681595
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14996 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_167
timestamp 1604681595
transform 1 0 16468 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_178
timestamp 1604681595
transform 1 0 17480 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1604681595
transform 1 0 17848 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1604681595
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_193
timestamp 1604681595
transform 1 0 18860 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_201
timestamp 1604681595
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1604681595
transform 1 0 5612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6624 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_52
timestamp 1604681595
transform 1 0 5888 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10672 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1604681595
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_96
timestamp 1604681595
transform 1 0 9936 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_120
timestamp 1604681595
transform 1 0 12144 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_132
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_158
timestamp 1604681595
transform 1 0 15640 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_175
timestamp 1604681595
transform 1 0 17204 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_199
timestamp 1604681595
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_23
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_31
timestamp 1604681595
transform 1 0 3956 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_42
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_53
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_43
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_55
timestamp 1604681595
transform 1 0 6164 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 6900 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_67
timestamp 1604681595
transform 1 0 7268 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9108 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9936 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12144 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_112
timestamp 1604681595
transform 1 0 11408 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604681595
transform 1 0 13708 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_127
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_144
timestamp 1604681595
transform 1 0 14352 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15088 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_161
timestamp 1604681595
transform 1 0 15916 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 18308 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604681595
transform 1 0 16652 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_173
timestamp 1604681595
transform 1 0 17020 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_184
timestamp 1604681595
transform 1 0 18032 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18768 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_191
timestamp 1604681595
transform 1 0 18676 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_19
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 4600 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1604681595
transform 1 0 3588 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_30
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_41
timestamp 1604681595
transform 1 0 4876 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8096 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_68
timestamp 1604681595
transform 1 0 7360 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1604681595
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15456 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_15_151
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1604681595
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_188
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_212
timestamp 1604681595
transform 1 0 20608 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_12
timestamp 1604681595
transform 1 0 2208 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 4232 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_38
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_50
timestamp 1604681595
transform 1 0 5704 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_67
timestamp 1604681595
transform 1 0 7268 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_126
timestamp 1604681595
transform 1 0 12696 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15364 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_164
timestamp 1604681595
transform 1 0 16192 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16928 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1604681595
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_188
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_194
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1604681595
transform 1 0 1472 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_18
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_35
timestamp 1604681595
transform 1 0 4324 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_52
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1604681595
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_78
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_95
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_112
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_148
timestamp 1604681595
transform 1 0 14720 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1604681595
transform 1 0 15640 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18124 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_175
timestamp 1604681595
transform 1 0 17204 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1604681595
transform 1 0 18676 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 1840 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_11
timestamp 1604681595
transform 1 0 2116 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6716 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_18_43
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_55
timestamp 1604681595
transform 1 0 6164 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_99
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_123
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_140
timestamp 1604681595
transform 1 0 13984 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_157
timestamp 1604681595
transform 1 0 15548 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17848 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_174
timestamp 1604681595
transform 1 0 17112 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_198
timestamp 1604681595
transform 1 0 19320 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1604681595
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4140 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_39
timestamp 1604681595
transform 1 0 4692 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5428 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_48
timestamp 1604681595
transform 1 0 5520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604681595
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_63
timestamp 1604681595
transform 1 0 6900 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_88
timestamp 1604681595
transform 1 0 9200 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 11316 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_115
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1604681595
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 12512 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_105
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13616 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_128
timestamp 1604681595
transform 1 0 12880 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_139
timestamp 1604681595
transform 1 0 13892 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 14628 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_152
timestamp 1604681595
transform 1 0 15088 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_164
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1604681595
transform 1 0 17572 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_189
timestamp 1604681595
transform 1 0 18492 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_210
timestamp 1604681595
transform 1 0 20424 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1604681595
transform 1 0 21528 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_10
timestamp 1604681595
transform 1 0 2024 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7268 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1604681595
transform 1 0 7176 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_76
timestamp 1604681595
transform 1 0 8096 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_84
timestamp 1604681595
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_133
timestamp 1604681595
transform 1 0 13340 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_141
timestamp 1604681595
transform 1 0 14076 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_170
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19780 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_195
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_212
timestamp 1604681595
transform 1 0 20608 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 2852 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_11
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10028 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1604681595
transform 1 0 9844 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11592 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1604681595
transform 1 0 10856 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_123
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_140
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16192 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 14904 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_148
timestamp 1604681595
transform 1 0 14720 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_162
timestamp 1604681595
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_180
timestamp 1604681595
transform 1 0 17664 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_20
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3680 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_44
timestamp 1604681595
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_56
timestamp 1604681595
transform 1 0 6256 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1604681595
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1604681595
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_80
timestamp 1604681595
transform 1 0 8464 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9200 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1604681595
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_116
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_139
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_156
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1604681595
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18584 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_23_206
timestamp 1604681595
transform 1 0 20056 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1604681595
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_9
timestamp 1604681595
transform 1 0 1932 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4324 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5888 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_76
timestamp 1604681595
transform 1 0 8096 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1604681595
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11776 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_107
timestamp 1604681595
transform 1 0 10948 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_115
timestamp 1604681595
transform 1 0 11684 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1604681595
transform 1 0 13248 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_140
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15916 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_170
timestamp 1604681595
transform 1 0 16744 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_194
timestamp 1604681595
transform 1 0 18952 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_19
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_82
timestamp 1604681595
transform 1 0 8648 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_95
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604681595
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_134
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1604681595
transform 1 0 15640 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 19688 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_201
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_9
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6624 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_54
timestamp 1604681595
transform 1 0 6072 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_46
timestamp 1604681595
transform 1 0 5336 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_26_76
timestamp 1604681595
transform 1 0 8096 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_71
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_79
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_97
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 13984 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_144
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 15364 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15088 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_159
timestamp 1604681595
transform 1 0 15732 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_161
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16468 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_183
timestamp 1604681595
transform 1 0 17940 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18676 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_200
timestamp 1604681595
transform 1 0 19504 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_195
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1604681595
transform 1 0 21528 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4508 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_46
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_54
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_64
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_72
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_82
timestamp 1604681595
transform 1 0 8648 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_99
timestamp 1604681595
transform 1 0 10212 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_135
timestamp 1604681595
transform 1 0 13524 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_162
timestamp 1604681595
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_179
timestamp 1604681595
transform 1 0 17572 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_187
timestamp 1604681595
transform 1 0 18308 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1604681595
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1604681595
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_7
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_43
timestamp 1604681595
transform 1 0 5060 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_79
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_91
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13708 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_129
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_146
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1604681595
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 16836 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_200
timestamp 1604681595
transform 1 0 19504 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_222
timestamp 1604681595
transform 1 0 21528 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4140 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_39
timestamp 1604681595
transform 1 0 4692 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5428 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_63
timestamp 1604681595
transform 1 0 6900 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10304 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_99
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_30_116
timestamp 1604681595
transform 1 0 11776 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_140
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_157
timestamp 1604681595
transform 1 0 15548 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1604681595
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_181
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18492 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1604681595
transform 1 0 19320 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_17
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3404 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8096 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_68
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_92
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_109
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1604681595
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_190
timestamp 1604681595
transform 1 0 18584 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_198
timestamp 1604681595
transform 1 0 19320 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1604681595
transform 1 0 21528 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_11
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_50
timestamp 1604681595
transform 1 0 5704 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_62
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_32_79
timestamp 1604681595
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1604681595
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_136
timestamp 1604681595
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1604681595
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1604681595
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_163
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16836 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18124 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_191
timestamp 1604681595
transform 1 0 18676 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_199
timestamp 1604681595
transform 1 0 19412 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_206
timestamp 1604681595
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 2852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_32
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_47
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_33_72
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_80
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_100
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 12696 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_33_130
timestamp 1604681595
transform 1 0 13064 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_147
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_165
timestamp 1604681595
transform 1 0 16284 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 17112 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1604681595
transform 1 0 17020 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_178
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1604681595
transform 1 0 18860 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_201
timestamp 1604681595
transform 1 0 19596 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_216
timestamp 1604681595
transform 1 0 20976 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_1_
port 0 nsew default input
rlabel metal3 s 0 5720 480 5840 6 ccff_head
port 1 nsew default input
rlabel metal3 s 0 17144 480 17264 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 22520 3816 23000 3936 6 chanx_right_in[0]
port 3 nsew default input
rlabel metal3 s 22520 8576 23000 8696 6 chanx_right_in[10]
port 4 nsew default input
rlabel metal3 s 22520 8984 23000 9104 6 chanx_right_in[11]
port 5 nsew default input
rlabel metal3 s 22520 9392 23000 9512 6 chanx_right_in[12]
port 6 nsew default input
rlabel metal3 s 22520 9936 23000 10056 6 chanx_right_in[13]
port 7 nsew default input
rlabel metal3 s 22520 10344 23000 10464 6 chanx_right_in[14]
port 8 nsew default input
rlabel metal3 s 22520 10888 23000 11008 6 chanx_right_in[15]
port 9 nsew default input
rlabel metal3 s 22520 11296 23000 11416 6 chanx_right_in[16]
port 10 nsew default input
rlabel metal3 s 22520 11840 23000 11960 6 chanx_right_in[17]
port 11 nsew default input
rlabel metal3 s 22520 12248 23000 12368 6 chanx_right_in[18]
port 12 nsew default input
rlabel metal3 s 22520 12792 23000 12912 6 chanx_right_in[19]
port 13 nsew default input
rlabel metal3 s 22520 4360 23000 4480 6 chanx_right_in[1]
port 14 nsew default input
rlabel metal3 s 22520 4768 23000 4888 6 chanx_right_in[2]
port 15 nsew default input
rlabel metal3 s 22520 5176 23000 5296 6 chanx_right_in[3]
port 16 nsew default input
rlabel metal3 s 22520 5720 23000 5840 6 chanx_right_in[4]
port 17 nsew default input
rlabel metal3 s 22520 6128 23000 6248 6 chanx_right_in[5]
port 18 nsew default input
rlabel metal3 s 22520 6672 23000 6792 6 chanx_right_in[6]
port 19 nsew default input
rlabel metal3 s 22520 7080 23000 7200 6 chanx_right_in[7]
port 20 nsew default input
rlabel metal3 s 22520 7624 23000 7744 6 chanx_right_in[8]
port 21 nsew default input
rlabel metal3 s 22520 8032 23000 8152 6 chanx_right_in[9]
port 22 nsew default input
rlabel metal3 s 22520 13200 23000 13320 6 chanx_right_out[0]
port 23 nsew default tristate
rlabel metal3 s 22520 17960 23000 18080 6 chanx_right_out[10]
port 24 nsew default tristate
rlabel metal3 s 22520 18368 23000 18488 6 chanx_right_out[11]
port 25 nsew default tristate
rlabel metal3 s 22520 18776 23000 18896 6 chanx_right_out[12]
port 26 nsew default tristate
rlabel metal3 s 22520 19320 23000 19440 6 chanx_right_out[13]
port 27 nsew default tristate
rlabel metal3 s 22520 19728 23000 19848 6 chanx_right_out[14]
port 28 nsew default tristate
rlabel metal3 s 22520 20272 23000 20392 6 chanx_right_out[15]
port 29 nsew default tristate
rlabel metal3 s 22520 20680 23000 20800 6 chanx_right_out[16]
port 30 nsew default tristate
rlabel metal3 s 22520 21224 23000 21344 6 chanx_right_out[17]
port 31 nsew default tristate
rlabel metal3 s 22520 21632 23000 21752 6 chanx_right_out[18]
port 32 nsew default tristate
rlabel metal3 s 22520 22176 23000 22296 6 chanx_right_out[19]
port 33 nsew default tristate
rlabel metal3 s 22520 13744 23000 13864 6 chanx_right_out[1]
port 34 nsew default tristate
rlabel metal3 s 22520 14152 23000 14272 6 chanx_right_out[2]
port 35 nsew default tristate
rlabel metal3 s 22520 14560 23000 14680 6 chanx_right_out[3]
port 36 nsew default tristate
rlabel metal3 s 22520 15104 23000 15224 6 chanx_right_out[4]
port 37 nsew default tristate
rlabel metal3 s 22520 15512 23000 15632 6 chanx_right_out[5]
port 38 nsew default tristate
rlabel metal3 s 22520 16056 23000 16176 6 chanx_right_out[6]
port 39 nsew default tristate
rlabel metal3 s 22520 16464 23000 16584 6 chanx_right_out[7]
port 40 nsew default tristate
rlabel metal3 s 22520 17008 23000 17128 6 chanx_right_out[8]
port 41 nsew default tristate
rlabel metal3 s 22520 17416 23000 17536 6 chanx_right_out[9]
port 42 nsew default tristate
rlabel metal2 s 846 0 902 480 6 chany_bottom_in[0]
port 43 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[10]
port 44 nsew default input
rlabel metal2 s 7010 0 7066 480 6 chany_bottom_in[11]
port 45 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[12]
port 46 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[13]
port 47 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[14]
port 48 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[15]
port 49 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[16]
port 50 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[17]
port 51 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[18]
port 52 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[19]
port 53 nsew default input
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_in[1]
port 54 nsew default input
rlabel metal2 s 1950 0 2006 480 6 chany_bottom_in[2]
port 55 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[3]
port 56 nsew default input
rlabel metal2 s 3054 0 3110 480 6 chany_bottom_in[4]
port 57 nsew default input
rlabel metal2 s 3606 0 3662 480 6 chany_bottom_in[5]
port 58 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[6]
port 59 nsew default input
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[7]
port 60 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[8]
port 61 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[9]
port 62 nsew default input
rlabel metal2 s 12070 0 12126 480 6 chany_bottom_out[0]
port 63 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[10]
port 64 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[11]
port 65 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[12]
port 66 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[13]
port 67 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[14]
port 68 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[15]
port 69 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[16]
port 70 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[17]
port 71 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[18]
port 72 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[19]
port 73 nsew default tristate
rlabel metal2 s 12622 0 12678 480 6 chany_bottom_out[1]
port 74 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[2]
port 75 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[3]
port 76 nsew default tristate
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_out[4]
port 77 nsew default tristate
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_out[5]
port 78 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[6]
port 79 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[7]
port 80 nsew default tristate
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[8]
port 81 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[9]
port 82 nsew default tristate
rlabel metal2 s 846 22520 902 23000 6 chany_top_in[0]
port 83 nsew default input
rlabel metal2 s 6458 22520 6514 23000 6 chany_top_in[10]
port 84 nsew default input
rlabel metal2 s 7010 22520 7066 23000 6 chany_top_in[11]
port 85 nsew default input
rlabel metal2 s 7562 22520 7618 23000 6 chany_top_in[12]
port 86 nsew default input
rlabel metal2 s 8114 22520 8170 23000 6 chany_top_in[13]
port 87 nsew default input
rlabel metal2 s 8666 22520 8722 23000 6 chany_top_in[14]
port 88 nsew default input
rlabel metal2 s 9218 22520 9274 23000 6 chany_top_in[15]
port 89 nsew default input
rlabel metal2 s 9770 22520 9826 23000 6 chany_top_in[16]
port 90 nsew default input
rlabel metal2 s 10322 22520 10378 23000 6 chany_top_in[17]
port 91 nsew default input
rlabel metal2 s 10874 22520 10930 23000 6 chany_top_in[18]
port 92 nsew default input
rlabel metal2 s 11426 22520 11482 23000 6 chany_top_in[19]
port 93 nsew default input
rlabel metal2 s 1398 22520 1454 23000 6 chany_top_in[1]
port 94 nsew default input
rlabel metal2 s 1950 22520 2006 23000 6 chany_top_in[2]
port 95 nsew default input
rlabel metal2 s 2502 22520 2558 23000 6 chany_top_in[3]
port 96 nsew default input
rlabel metal2 s 3054 22520 3110 23000 6 chany_top_in[4]
port 97 nsew default input
rlabel metal2 s 3606 22520 3662 23000 6 chany_top_in[5]
port 98 nsew default input
rlabel metal2 s 4158 22520 4214 23000 6 chany_top_in[6]
port 99 nsew default input
rlabel metal2 s 4710 22520 4766 23000 6 chany_top_in[7]
port 100 nsew default input
rlabel metal2 s 5262 22520 5318 23000 6 chany_top_in[8]
port 101 nsew default input
rlabel metal2 s 5814 22520 5870 23000 6 chany_top_in[9]
port 102 nsew default input
rlabel metal2 s 12070 22520 12126 23000 6 chany_top_out[0]
port 103 nsew default tristate
rlabel metal2 s 17682 22520 17738 23000 6 chany_top_out[10]
port 104 nsew default tristate
rlabel metal2 s 18234 22520 18290 23000 6 chany_top_out[11]
port 105 nsew default tristate
rlabel metal2 s 18786 22520 18842 23000 6 chany_top_out[12]
port 106 nsew default tristate
rlabel metal2 s 19338 22520 19394 23000 6 chany_top_out[13]
port 107 nsew default tristate
rlabel metal2 s 19890 22520 19946 23000 6 chany_top_out[14]
port 108 nsew default tristate
rlabel metal2 s 20442 22520 20498 23000 6 chany_top_out[15]
port 109 nsew default tristate
rlabel metal2 s 20994 22520 21050 23000 6 chany_top_out[16]
port 110 nsew default tristate
rlabel metal2 s 21546 22520 21602 23000 6 chany_top_out[17]
port 111 nsew default tristate
rlabel metal2 s 22098 22520 22154 23000 6 chany_top_out[18]
port 112 nsew default tristate
rlabel metal2 s 22650 22520 22706 23000 6 chany_top_out[19]
port 113 nsew default tristate
rlabel metal2 s 12622 22520 12678 23000 6 chany_top_out[1]
port 114 nsew default tristate
rlabel metal2 s 13174 22520 13230 23000 6 chany_top_out[2]
port 115 nsew default tristate
rlabel metal2 s 13726 22520 13782 23000 6 chany_top_out[3]
port 116 nsew default tristate
rlabel metal2 s 14278 22520 14334 23000 6 chany_top_out[4]
port 117 nsew default tristate
rlabel metal2 s 14830 22520 14886 23000 6 chany_top_out[5]
port 118 nsew default tristate
rlabel metal2 s 15382 22520 15438 23000 6 chany_top_out[6]
port 119 nsew default tristate
rlabel metal2 s 15934 22520 15990 23000 6 chany_top_out[7]
port 120 nsew default tristate
rlabel metal2 s 16486 22520 16542 23000 6 chany_top_out[8]
port 121 nsew default tristate
rlabel metal2 s 17038 22520 17094 23000 6 chany_top_out[9]
port 122 nsew default tristate
rlabel metal3 s 22520 22584 23000 22704 6 prog_clk
port 123 nsew default input
rlabel metal3 s 22520 144 23000 264 6 right_bottom_grid_pin_34_
port 124 nsew default input
rlabel metal3 s 22520 552 23000 672 6 right_bottom_grid_pin_35_
port 125 nsew default input
rlabel metal3 s 22520 960 23000 1080 6 right_bottom_grid_pin_36_
port 126 nsew default input
rlabel metal3 s 22520 1504 23000 1624 6 right_bottom_grid_pin_37_
port 127 nsew default input
rlabel metal3 s 22520 1912 23000 2032 6 right_bottom_grid_pin_38_
port 128 nsew default input
rlabel metal3 s 22520 2456 23000 2576 6 right_bottom_grid_pin_39_
port 129 nsew default input
rlabel metal3 s 22520 2864 23000 2984 6 right_bottom_grid_pin_40_
port 130 nsew default input
rlabel metal3 s 22520 3408 23000 3528 6 right_bottom_grid_pin_41_
port 131 nsew default input
rlabel metal2 s 294 22520 350 23000 6 top_left_grid_pin_1_
port 132 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 133 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 134 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
