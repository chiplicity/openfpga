VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__0_
  CLASS BLOCK ;
  FOREIGN sb_2__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 138.395 BY 140.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 2.400 33.280 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 2.400 41.440 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 2.400 44.840 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 2.400 16.280 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 2.400 19.000 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 2.400 27.160 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 2.400 30.560 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 2.400 90.400 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 2.400 93.120 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 2.400 95.840 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 2.400 98.560 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 2.400 104.680 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 2.400 107.400 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 2.400 110.120 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 2.400 116.240 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 2.400 70.000 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 2.400 76.120 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 2.400 78.840 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 2.400 81.560 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 2.400 84.280 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.400 87.680 ;
    END
  END chanx_left_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.530 137.600 52.810 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 137.600 55.570 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.510 137.600 58.790 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.030 137.600 64.310 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 137.600 67.070 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 137.600 69.830 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 137.600 73.050 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.530 137.600 75.810 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 137.600 78.570 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 137.600 27.050 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 137.600 30.270 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 137.600 33.030 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 137.600 35.790 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 137.600 41.310 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 137.600 44.530 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 137.600 47.290 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 137.600 50.050 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 137.600 109.850 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.330 137.600 112.610 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.550 137.600 115.830 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.310 137.600 118.590 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.830 137.600 124.110 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.590 137.600 126.870 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 137.600 130.090 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 137.600 132.850 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.330 137.600 135.610 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 137.600 84.090 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 137.600 90.070 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 137.600 92.830 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.310 137.600 95.590 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.070 137.600 98.350 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 137.600 101.570 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.050 137.600 104.330 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 106.810 137.600 107.090 140.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 2.400 118.960 ;
    END
  END left_top_grid_pin_42_
  PIN left_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 2.400 121.680 ;
    END
  END left_top_grid_pin_43_
  PIN left_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 2.400 124.400 ;
    END
  END left_top_grid_pin_44_
  PIN left_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 2.400 127.120 ;
    END
  END left_top_grid_pin_45_
  PIN left_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 2.400 130.520 ;
    END
  END left_top_grid_pin_46_
  PIN left_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 2.400 133.240 ;
    END
  END left_top_grid_pin_47_
  PIN left_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 135.360 2.400 135.960 ;
    END
  END left_top_grid_pin_48_
  PIN left_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 2.400 138.680 ;
    END
  END left_top_grid_pin_49_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 2.400 ;
    END
  END prog_clk
  PIN top_left_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_34_
  PIN top_left_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 137.600 4.510 140.000 ;
    END
  END top_left_grid_pin_35_
  PIN top_left_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 137.600 7.270 140.000 ;
    END
  END top_left_grid_pin_36_
  PIN top_left_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 137.600 10.030 140.000 ;
    END
  END top_left_grid_pin_37_
  PIN top_left_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 137.600 12.790 140.000 ;
    END
  END top_left_grid_pin_38_
  PIN top_left_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 137.600 16.010 140.000 ;
    END
  END top_left_grid_pin_39_
  PIN top_left_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 137.600 18.770 140.000 ;
    END
  END top_left_grid_pin_40_
  PIN top_left_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 137.600 21.530 140.000 ;
    END
  END top_left_grid_pin_41_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.090 137.600 138.370 140.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 2.830 10.640 134.320 128.080 ;
      LAYER met2 ;
        RECT 1.010 137.320 1.190 138.565 ;
        RECT 2.030 137.320 3.950 138.565 ;
        RECT 4.790 137.320 6.710 138.565 ;
        RECT 7.550 137.320 9.470 138.565 ;
        RECT 10.310 137.320 12.230 138.565 ;
        RECT 13.070 137.320 15.450 138.565 ;
        RECT 16.290 137.320 18.210 138.565 ;
        RECT 19.050 137.320 20.970 138.565 ;
        RECT 21.810 137.320 23.730 138.565 ;
        RECT 24.570 137.320 26.490 138.565 ;
        RECT 27.330 137.320 29.710 138.565 ;
        RECT 30.550 137.320 32.470 138.565 ;
        RECT 33.310 137.320 35.230 138.565 ;
        RECT 36.070 137.320 37.990 138.565 ;
        RECT 38.830 137.320 40.750 138.565 ;
        RECT 41.590 137.320 43.970 138.565 ;
        RECT 44.810 137.320 46.730 138.565 ;
        RECT 47.570 137.320 49.490 138.565 ;
        RECT 50.330 137.320 52.250 138.565 ;
        RECT 53.090 137.320 55.010 138.565 ;
        RECT 55.850 137.320 58.230 138.565 ;
        RECT 59.070 137.320 60.990 138.565 ;
        RECT 61.830 137.320 63.750 138.565 ;
        RECT 64.590 137.320 66.510 138.565 ;
        RECT 67.350 137.320 69.270 138.565 ;
        RECT 70.110 137.320 72.490 138.565 ;
        RECT 73.330 137.320 75.250 138.565 ;
        RECT 76.090 137.320 78.010 138.565 ;
        RECT 78.850 137.320 80.770 138.565 ;
        RECT 81.610 137.320 83.530 138.565 ;
        RECT 84.370 137.320 86.750 138.565 ;
        RECT 87.590 137.320 89.510 138.565 ;
        RECT 90.350 137.320 92.270 138.565 ;
        RECT 93.110 137.320 95.030 138.565 ;
        RECT 95.870 137.320 97.790 138.565 ;
        RECT 98.630 137.320 101.010 138.565 ;
        RECT 101.850 137.320 103.770 138.565 ;
        RECT 104.610 137.320 106.530 138.565 ;
        RECT 107.370 137.320 109.290 138.565 ;
        RECT 110.130 137.320 112.050 138.565 ;
        RECT 112.890 137.320 115.270 138.565 ;
        RECT 116.110 137.320 118.030 138.565 ;
        RECT 118.870 137.320 120.790 138.565 ;
        RECT 121.630 137.320 123.550 138.565 ;
        RECT 124.390 137.320 126.310 138.565 ;
        RECT 127.150 137.320 129.530 138.565 ;
        RECT 130.370 137.320 132.290 138.565 ;
        RECT 133.130 137.320 135.050 138.565 ;
        RECT 135.890 137.320 137.810 138.565 ;
        RECT 1.010 2.680 138.370 137.320 ;
        RECT 1.010 1.515 22.810 2.680 ;
        RECT 23.650 1.515 69.270 2.680 ;
        RECT 70.110 1.515 115.730 2.680 ;
        RECT 116.570 1.515 138.370 2.680 ;
      LAYER met3 ;
        RECT 2.800 137.680 138.395 138.545 ;
        RECT 0.985 136.360 138.395 137.680 ;
        RECT 2.800 134.960 138.395 136.360 ;
        RECT 0.985 133.640 138.395 134.960 ;
        RECT 2.800 132.240 138.395 133.640 ;
        RECT 0.985 130.920 138.395 132.240 ;
        RECT 2.800 129.520 138.395 130.920 ;
        RECT 0.985 127.520 138.395 129.520 ;
        RECT 2.800 126.120 138.395 127.520 ;
        RECT 0.985 124.800 138.395 126.120 ;
        RECT 2.800 123.400 138.395 124.800 ;
        RECT 0.985 122.080 138.395 123.400 ;
        RECT 2.800 120.680 138.395 122.080 ;
        RECT 0.985 119.360 138.395 120.680 ;
        RECT 2.800 117.960 138.395 119.360 ;
        RECT 0.985 116.640 138.395 117.960 ;
        RECT 2.800 115.240 138.395 116.640 ;
        RECT 0.985 113.240 138.395 115.240 ;
        RECT 2.800 111.840 138.395 113.240 ;
        RECT 0.985 110.520 138.395 111.840 ;
        RECT 2.800 109.120 138.395 110.520 ;
        RECT 0.985 107.800 138.395 109.120 ;
        RECT 2.800 106.400 138.395 107.800 ;
        RECT 0.985 105.080 138.395 106.400 ;
        RECT 2.800 103.680 138.395 105.080 ;
        RECT 0.985 102.360 138.395 103.680 ;
        RECT 2.800 100.960 138.395 102.360 ;
        RECT 0.985 98.960 138.395 100.960 ;
        RECT 2.800 97.560 138.395 98.960 ;
        RECT 0.985 96.240 138.395 97.560 ;
        RECT 2.800 94.840 138.395 96.240 ;
        RECT 0.985 93.520 138.395 94.840 ;
        RECT 2.800 92.120 138.395 93.520 ;
        RECT 0.985 90.800 138.395 92.120 ;
        RECT 2.800 89.400 138.395 90.800 ;
        RECT 0.985 88.080 138.395 89.400 ;
        RECT 2.800 86.680 138.395 88.080 ;
        RECT 0.985 84.680 138.395 86.680 ;
        RECT 2.800 83.280 138.395 84.680 ;
        RECT 0.985 81.960 138.395 83.280 ;
        RECT 2.800 80.560 138.395 81.960 ;
        RECT 0.985 79.240 138.395 80.560 ;
        RECT 2.800 77.840 138.395 79.240 ;
        RECT 0.985 76.520 138.395 77.840 ;
        RECT 2.800 75.120 138.395 76.520 ;
        RECT 0.985 73.800 138.395 75.120 ;
        RECT 2.800 72.400 138.395 73.800 ;
        RECT 0.985 70.400 138.395 72.400 ;
        RECT 2.800 69.000 138.395 70.400 ;
        RECT 0.985 67.680 138.395 69.000 ;
        RECT 2.800 66.280 138.395 67.680 ;
        RECT 0.985 64.960 138.395 66.280 ;
        RECT 2.800 63.560 138.395 64.960 ;
        RECT 0.985 62.240 138.395 63.560 ;
        RECT 2.800 60.840 138.395 62.240 ;
        RECT 0.985 59.520 138.395 60.840 ;
        RECT 2.800 58.120 138.395 59.520 ;
        RECT 0.985 56.120 138.395 58.120 ;
        RECT 2.800 54.720 138.395 56.120 ;
        RECT 0.985 53.400 138.395 54.720 ;
        RECT 2.800 52.000 138.395 53.400 ;
        RECT 0.985 50.680 138.395 52.000 ;
        RECT 2.800 49.280 138.395 50.680 ;
        RECT 0.985 47.960 138.395 49.280 ;
        RECT 2.800 46.560 138.395 47.960 ;
        RECT 0.985 45.240 138.395 46.560 ;
        RECT 2.800 43.840 138.395 45.240 ;
        RECT 0.985 41.840 138.395 43.840 ;
        RECT 2.800 40.440 138.395 41.840 ;
        RECT 0.985 39.120 138.395 40.440 ;
        RECT 2.800 37.720 138.395 39.120 ;
        RECT 0.985 36.400 138.395 37.720 ;
        RECT 2.800 35.000 138.395 36.400 ;
        RECT 0.985 33.680 138.395 35.000 ;
        RECT 2.800 32.280 138.395 33.680 ;
        RECT 0.985 30.960 138.395 32.280 ;
        RECT 2.800 29.560 138.395 30.960 ;
        RECT 0.985 27.560 138.395 29.560 ;
        RECT 2.800 26.160 138.395 27.560 ;
        RECT 0.985 24.840 138.395 26.160 ;
        RECT 2.800 23.440 138.395 24.840 ;
        RECT 0.985 22.120 138.395 23.440 ;
        RECT 2.800 20.720 138.395 22.120 ;
        RECT 0.985 19.400 138.395 20.720 ;
        RECT 2.800 18.000 138.395 19.400 ;
        RECT 0.985 16.680 138.395 18.000 ;
        RECT 2.800 15.280 138.395 16.680 ;
        RECT 0.985 13.280 138.395 15.280 ;
        RECT 2.800 11.880 138.395 13.280 ;
        RECT 0.985 10.560 138.395 11.880 ;
        RECT 2.800 9.160 138.395 10.560 ;
        RECT 0.985 7.840 138.395 9.160 ;
        RECT 2.800 6.440 138.395 7.840 ;
        RECT 0.985 5.120 138.395 6.440 ;
        RECT 2.800 3.720 138.395 5.120 ;
        RECT 0.985 2.400 138.395 3.720 ;
        RECT 2.800 1.535 138.395 2.400 ;
      LAYER met4 ;
        RECT 26.550 10.640 27.655 128.080 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
      LAYER met5 ;
        RECT 26.340 79.100 78.540 80.700 ;
  END
END sb_2__0_
END LIBRARY

