VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_1__1_
  CLASS BLOCK ;
  FOREIGN cby_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 200.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 2.400 8.800 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 197.600 3.590 200.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 2.400 25.120 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.400 ;
    END
  END address[5]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 8.880 80.000 9.480 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 2.400 42.120 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 197.600 10.490 200.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.570 197.600 17.850 200.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 26.560 80.000 27.160 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 44.920 80.000 45.520 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 197.600 25.210 200.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.400 108.760 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 63.280 80.000 63.880 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 80.960 80.000 81.560 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.400 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 197.600 32.570 200.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.400 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 197.600 39.930 200.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 99.320 80.000 99.920 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 197.600 46.830 200.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 2.400 125.080 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 77.600 117.680 80.000 118.280 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 2.400 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 197.600 54.190 200.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 2.400 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.270 197.600 61.550 200.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 136.040 80.000 136.640 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 2.400 142.080 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 2.400 158.400 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 2.400 175.400 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 153.720 80.000 154.320 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END enable
  PIN left_grid_pin_1_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 172.080 80.000 172.680 ;
    END
  END left_grid_pin_1_
  PIN left_grid_pin_5_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 77.600 190.440 80.000 191.040 ;
    END
  END left_grid_pin_5_
  PIN left_grid_pin_9_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.630 197.600 68.910 200.000 ;
    END
  END left_grid_pin_9_
  PIN right_grid_pin_3_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 2.400 191.720 ;
    END
  END right_grid_pin_3_
  PIN right_grid_pin_7_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 197.600 76.270 200.000 ;
    END
  END right_grid_pin_7_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 18.055 10.640 19.655 187.920 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 31.385 10.640 32.985 187.920 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 74.060 187.765 ;
      LAYER met1 ;
        RECT 0.070 0.380 76.290 198.520 ;
      LAYER met2 ;
        RECT 0.100 197.320 3.030 198.550 ;
        RECT 3.870 197.320 9.930 198.550 ;
        RECT 10.770 197.320 17.290 198.550 ;
        RECT 18.130 197.320 24.650 198.550 ;
        RECT 25.490 197.320 32.010 198.550 ;
        RECT 32.850 197.320 39.370 198.550 ;
        RECT 40.210 197.320 46.270 198.550 ;
        RECT 47.110 197.320 53.630 198.550 ;
        RECT 54.470 197.320 60.990 198.550 ;
        RECT 61.830 197.320 68.350 198.550 ;
        RECT 69.190 197.320 75.710 198.550 ;
        RECT 76.550 197.320 77.650 198.550 ;
        RECT 0.100 2.680 77.650 197.320 ;
        RECT 0.100 0.270 2.110 2.680 ;
        RECT 2.950 0.270 7.170 2.680 ;
        RECT 8.010 0.270 12.690 2.680 ;
        RECT 13.530 0.270 17.750 2.680 ;
        RECT 18.590 0.270 23.270 2.680 ;
        RECT 24.110 0.270 28.790 2.680 ;
        RECT 29.630 0.270 33.850 2.680 ;
        RECT 34.690 0.270 39.370 2.680 ;
        RECT 40.210 0.270 44.430 2.680 ;
        RECT 45.270 0.270 49.950 2.680 ;
        RECT 50.790 0.270 55.470 2.680 ;
        RECT 56.310 0.270 60.530 2.680 ;
        RECT 61.370 0.270 66.050 2.680 ;
        RECT 66.890 0.270 71.110 2.680 ;
        RECT 71.950 0.270 76.630 2.680 ;
        RECT 77.470 0.270 77.650 2.680 ;
      LAYER met3 ;
        RECT 2.800 190.720 77.200 191.120 ;
        RECT 0.270 190.040 77.200 190.720 ;
        RECT 0.270 175.800 77.890 190.040 ;
        RECT 2.800 174.400 77.890 175.800 ;
        RECT 0.270 173.080 77.890 174.400 ;
        RECT 0.270 171.680 77.200 173.080 ;
        RECT 0.270 158.800 77.890 171.680 ;
        RECT 2.800 157.400 77.890 158.800 ;
        RECT 0.270 154.720 77.890 157.400 ;
        RECT 0.270 153.320 77.200 154.720 ;
        RECT 0.270 142.480 77.890 153.320 ;
        RECT 2.800 141.080 77.890 142.480 ;
        RECT 0.270 137.040 77.890 141.080 ;
        RECT 0.270 135.640 77.200 137.040 ;
        RECT 0.270 125.480 77.890 135.640 ;
        RECT 2.800 124.080 77.890 125.480 ;
        RECT 0.270 118.680 77.890 124.080 ;
        RECT 0.270 117.280 77.200 118.680 ;
        RECT 0.270 109.160 77.890 117.280 ;
        RECT 2.800 107.760 77.890 109.160 ;
        RECT 0.270 100.320 77.890 107.760 ;
        RECT 0.270 98.920 77.200 100.320 ;
        RECT 0.270 92.160 77.890 98.920 ;
        RECT 2.800 90.760 77.890 92.160 ;
        RECT 0.270 81.960 77.890 90.760 ;
        RECT 0.270 80.560 77.200 81.960 ;
        RECT 0.270 75.840 77.890 80.560 ;
        RECT 2.800 74.440 77.890 75.840 ;
        RECT 0.270 64.280 77.890 74.440 ;
        RECT 0.270 62.880 77.200 64.280 ;
        RECT 0.270 58.840 77.890 62.880 ;
        RECT 2.800 57.440 77.890 58.840 ;
        RECT 0.270 45.920 77.890 57.440 ;
        RECT 0.270 44.520 77.200 45.920 ;
        RECT 0.270 42.520 77.890 44.520 ;
        RECT 2.800 41.120 77.890 42.520 ;
        RECT 0.270 27.560 77.890 41.120 ;
        RECT 0.270 26.160 77.200 27.560 ;
        RECT 0.270 25.520 77.890 26.160 ;
        RECT 2.800 24.120 77.890 25.520 ;
        RECT 0.270 9.880 77.890 24.120 ;
        RECT 0.270 9.200 77.200 9.880 ;
        RECT 2.800 8.800 77.200 9.200 ;
      LAYER met4 ;
        RECT 0.295 10.640 17.655 187.920 ;
        RECT 20.055 10.640 30.985 187.920 ;
        RECT 33.385 10.640 72.985 187.920 ;
  END
END cby_1__1_
END LIBRARY

