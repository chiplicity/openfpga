magic
tech sky130A
magscale 1 2
timestamp 1605123025
<< locali >>
rect 3893 21335 3927 21505
rect 6101 14467 6135 14569
rect 6377 11679 6411 11781
rect 2881 11067 2915 11305
<< viali >>
rect 5641 25449 5675 25483
rect 7389 25449 7423 25483
rect 8677 25449 8711 25483
rect 11069 25449 11103 25483
rect 13645 25449 13679 25483
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4905 25313 4939 25347
rect 4997 25313 5031 25347
rect 7297 25313 7331 25347
rect 8493 25313 8527 25347
rect 9781 25313 9815 25347
rect 10885 25313 10919 25347
rect 5089 25245 5123 25279
rect 7573 25245 7607 25279
rect 12633 25245 12667 25279
rect 3249 25177 3283 25211
rect 5917 25177 5951 25211
rect 6745 25177 6779 25211
rect 9965 25177 9999 25211
rect 1593 25109 1627 25143
rect 2697 25109 2731 25143
rect 4537 25109 4571 25143
rect 6929 25109 6963 25143
rect 10425 25109 10459 25143
rect 4629 24905 4663 24939
rect 9689 24905 9723 24939
rect 10885 24905 10919 24939
rect 8585 24837 8619 24871
rect 3617 24769 3651 24803
rect 3801 24769 3835 24803
rect 5733 24769 5767 24803
rect 6653 24769 6687 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 9045 24769 9079 24803
rect 10425 24769 10459 24803
rect 12265 24769 12299 24803
rect 13001 24769 13035 24803
rect 1409 24701 1443 24735
rect 3065 24701 3099 24735
rect 3525 24701 3559 24735
rect 5641 24701 5675 24735
rect 6285 24701 6319 24735
rect 8401 24701 8435 24735
rect 9413 24701 9447 24735
rect 7941 24633 7975 24667
rect 10241 24633 10275 24667
rect 11897 24633 11931 24667
rect 12909 24633 12943 24667
rect 14013 24633 14047 24667
rect 1593 24565 1627 24599
rect 1961 24565 1995 24599
rect 2329 24565 2363 24599
rect 3157 24565 3191 24599
rect 4169 24565 4203 24599
rect 4905 24565 4939 24599
rect 5181 24565 5215 24599
rect 5549 24565 5583 24599
rect 6837 24565 6871 24599
rect 7205 24565 7239 24599
rect 8309 24565 8343 24599
rect 9873 24565 9907 24599
rect 10333 24565 10367 24599
rect 12449 24565 12483 24599
rect 12817 24565 12851 24599
rect 3433 24361 3467 24395
rect 4629 24361 4663 24395
rect 9045 24361 9079 24395
rect 11529 24361 11563 24395
rect 11989 24361 12023 24395
rect 13093 24361 13127 24395
rect 15485 24361 15519 24395
rect 16589 24361 16623 24395
rect 18981 24361 19015 24395
rect 21097 24361 21131 24395
rect 4988 24293 5022 24327
rect 7288 24293 7322 24327
rect 10425 24293 10459 24327
rect 13553 24293 13587 24327
rect 1501 24225 1535 24259
rect 2789 24225 2823 24259
rect 4721 24225 4755 24259
rect 10333 24225 10367 24259
rect 11897 24225 11931 24259
rect 13461 24225 13495 24259
rect 15301 24225 15335 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 18797 24225 18831 24259
rect 20913 24225 20947 24259
rect 1777 24157 1811 24191
rect 6561 24157 6595 24191
rect 7021 24157 7055 24191
rect 9505 24157 9539 24191
rect 10517 24157 10551 24191
rect 12173 24157 12207 24191
rect 13737 24157 13771 24191
rect 11069 24089 11103 24123
rect 17693 24089 17727 24123
rect 2513 24021 2547 24055
rect 2973 24021 3007 24055
rect 6101 24021 6135 24055
rect 6929 24021 6963 24055
rect 8401 24021 8435 24055
rect 8677 24021 8711 24055
rect 9965 24021 9999 24055
rect 12633 24021 12667 24055
rect 13001 24021 13035 24055
rect 2513 23817 2547 23851
rect 2881 23817 2915 23851
rect 5365 23817 5399 23851
rect 5733 23817 5767 23851
rect 6653 23817 6687 23851
rect 9965 23817 9999 23851
rect 11805 23817 11839 23851
rect 12817 23817 12851 23851
rect 14289 23817 14323 23851
rect 15301 23817 15335 23851
rect 16405 23817 16439 23851
rect 18245 23817 18279 23851
rect 19349 23817 19383 23851
rect 20453 23817 20487 23851
rect 21557 23817 21591 23851
rect 22661 23817 22695 23851
rect 5089 23749 5123 23783
rect 8493 23749 8527 23783
rect 12173 23749 12207 23783
rect 9229 23681 9263 23715
rect 1685 23613 1719 23647
rect 3341 23613 3375 23647
rect 5549 23613 5583 23647
rect 7113 23613 7147 23647
rect 8769 23613 8803 23647
rect 10057 23613 10091 23647
rect 10324 23613 10358 23647
rect 12909 23613 12943 23647
rect 15117 23613 15151 23647
rect 16221 23613 16255 23647
rect 16773 23613 16807 23647
rect 18061 23613 18095 23647
rect 18613 23613 18647 23647
rect 19165 23613 19199 23647
rect 20269 23613 20303 23647
rect 20821 23613 20855 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 1961 23545 1995 23579
rect 3249 23545 3283 23579
rect 3586 23545 3620 23579
rect 6285 23545 6319 23579
rect 7358 23545 7392 23579
rect 13176 23545 13210 23579
rect 15669 23545 15703 23579
rect 17509 23545 17543 23579
rect 19717 23545 19751 23579
rect 4721 23477 4755 23511
rect 9505 23477 9539 23511
rect 11437 23477 11471 23511
rect 14565 23477 14599 23511
rect 16037 23477 16071 23511
rect 17141 23477 17175 23511
rect 18981 23477 19015 23511
rect 21189 23477 21223 23511
rect 2421 23273 2455 23307
rect 7021 23273 7055 23307
rect 8493 23273 8527 23307
rect 11253 23273 11287 23307
rect 11621 23273 11655 23307
rect 11989 23273 12023 23307
rect 14289 23273 14323 23307
rect 16773 23273 16807 23307
rect 19533 23273 19567 23307
rect 1869 23205 1903 23239
rect 4344 23205 4378 23239
rect 10140 23205 10174 23239
rect 15577 23205 15611 23239
rect 21189 23205 21223 23239
rect 1593 23137 1627 23171
rect 2881 23137 2915 23171
rect 3525 23137 3559 23171
rect 3893 23137 3927 23171
rect 4077 23137 4111 23171
rect 7113 23137 7147 23171
rect 7380 23137 7414 23171
rect 9137 23137 9171 23171
rect 9873 23137 9907 23171
rect 13165 23137 13199 23171
rect 15301 23137 15335 23171
rect 16589 23137 16623 23171
rect 19349 23137 19383 23171
rect 20913 23137 20947 23171
rect 12909 23069 12943 23103
rect 3065 22933 3099 22967
rect 5457 22933 5491 22967
rect 6469 22933 6503 22967
rect 9505 22933 9539 22967
rect 12449 22933 12483 22967
rect 12817 22933 12851 22967
rect 5825 22729 5859 22763
rect 6377 22729 6411 22763
rect 7297 22729 7331 22763
rect 10425 22729 10459 22763
rect 11897 22729 11931 22763
rect 14473 22729 14507 22763
rect 15761 22729 15795 22763
rect 3249 22661 3283 22695
rect 4813 22661 4847 22695
rect 12265 22661 12299 22695
rect 1777 22593 1811 22627
rect 3709 22593 3743 22627
rect 3801 22593 3835 22627
rect 4721 22593 4755 22627
rect 5273 22593 5307 22627
rect 5457 22593 5491 22627
rect 6285 22593 6319 22627
rect 7849 22593 7883 22627
rect 8677 22593 8711 22627
rect 9965 22593 9999 22627
rect 13093 22593 13127 22627
rect 15301 22593 15335 22627
rect 1501 22525 1535 22559
rect 2789 22525 2823 22559
rect 4353 22525 4387 22559
rect 5181 22525 5215 22559
rect 6561 22525 6595 22559
rect 7205 22525 7239 22559
rect 7757 22525 7791 22559
rect 9873 22525 9907 22559
rect 10793 22525 10827 22559
rect 11069 22525 11103 22559
rect 3157 22457 3191 22491
rect 3617 22457 3651 22491
rect 7665 22457 7699 22491
rect 8309 22457 8343 22491
rect 9321 22457 9355 22491
rect 11345 22457 11379 22491
rect 13001 22457 13035 22491
rect 13338 22457 13372 22491
rect 2421 22389 2455 22423
rect 9413 22389 9447 22423
rect 9781 22389 9815 22423
rect 14749 22389 14783 22423
rect 16589 22389 16623 22423
rect 19349 22389 19383 22423
rect 20913 22389 20947 22423
rect 2421 22185 2455 22219
rect 2697 22185 2731 22219
rect 3525 22185 3559 22219
rect 5825 22185 5859 22219
rect 6193 22185 6227 22219
rect 16313 22185 16347 22219
rect 3893 22117 3927 22151
rect 15301 22117 15335 22151
rect 1593 22049 1627 22083
rect 1869 22049 1903 22083
rect 2881 22049 2915 22083
rect 4344 22049 4378 22083
rect 6837 22049 6871 22083
rect 8309 22049 8343 22083
rect 9965 22049 9999 22083
rect 10232 22049 10266 22083
rect 12081 22049 12115 22083
rect 12357 22049 12391 22083
rect 12909 22049 12943 22083
rect 13257 22049 13291 22083
rect 4077 21981 4111 22015
rect 6929 21981 6963 22015
rect 7021 21981 7055 22015
rect 8493 21981 8527 22015
rect 13001 21981 13035 22015
rect 3065 21913 3099 21947
rect 12173 21913 12207 21947
rect 5457 21845 5491 21879
rect 6469 21845 6503 21879
rect 7665 21845 7699 21879
rect 8033 21845 8067 21879
rect 9413 21845 9447 21879
rect 11345 21845 11379 21879
rect 14381 21845 14415 21879
rect 2421 21641 2455 21675
rect 3709 21641 3743 21675
rect 4077 21641 4111 21675
rect 4905 21641 4939 21675
rect 5917 21641 5951 21675
rect 10425 21641 10459 21675
rect 13553 21641 13587 21675
rect 13921 21641 13955 21675
rect 2697 21573 2731 21607
rect 10977 21573 11011 21607
rect 12541 21573 12575 21607
rect 14105 21573 14139 21607
rect 3065 21505 3099 21539
rect 3893 21505 3927 21539
rect 7481 21505 7515 21539
rect 8033 21505 8067 21539
rect 8217 21505 8251 21539
rect 8861 21505 8895 21539
rect 9873 21505 9907 21539
rect 13001 21505 13035 21539
rect 13093 21505 13127 21539
rect 14565 21505 14599 21539
rect 14657 21505 14691 21539
rect 15117 21505 15151 21539
rect 15669 21505 15703 21539
rect 1593 21437 1627 21471
rect 2881 21437 2915 21471
rect 1869 21369 1903 21403
rect 4157 21437 4191 21471
rect 5273 21437 5307 21471
rect 7941 21437 7975 21471
rect 9229 21437 9263 21471
rect 9781 21437 9815 21471
rect 11069 21437 11103 21471
rect 12265 21437 12299 21471
rect 12909 21437 12943 21471
rect 14473 21437 14507 21471
rect 11345 21369 11379 21403
rect 11897 21369 11931 21403
rect 3893 21301 3927 21335
rect 4353 21301 4387 21335
rect 5457 21301 5491 21335
rect 6469 21301 6503 21335
rect 7021 21301 7055 21335
rect 7573 21301 7607 21335
rect 9321 21301 9355 21335
rect 9689 21301 9723 21335
rect 2973 21097 3007 21131
rect 3525 21097 3559 21131
rect 5733 21097 5767 21131
rect 6561 21097 6595 21131
rect 8125 21097 8159 21131
rect 8401 21097 8435 21131
rect 9321 21097 9355 21131
rect 11069 21097 11103 21131
rect 12081 21097 12115 21131
rect 12633 21097 12667 21131
rect 14381 21097 14415 21131
rect 4344 21029 4378 21063
rect 8769 21029 8803 21063
rect 9137 21029 9171 21063
rect 9934 21029 9968 21063
rect 1685 20961 1719 20995
rect 1961 20961 1995 20995
rect 4077 20961 4111 20995
rect 6745 20961 6779 20995
rect 7012 20961 7046 20995
rect 9505 20961 9539 20995
rect 11897 20961 11931 20995
rect 13257 20961 13291 20995
rect 9689 20893 9723 20927
rect 13001 20893 13035 20927
rect 2421 20757 2455 20791
rect 2789 20757 2823 20791
rect 3893 20757 3927 20791
rect 5457 20757 5491 20791
rect 6101 20757 6135 20791
rect 11437 20757 11471 20791
rect 14749 20757 14783 20791
rect 4445 20553 4479 20587
rect 6653 20553 6687 20587
rect 8217 20553 8251 20587
rect 8585 20553 8619 20587
rect 8953 20553 8987 20587
rect 10425 20553 10459 20587
rect 11161 20553 11195 20587
rect 11897 20553 11931 20587
rect 13001 20553 13035 20587
rect 14473 20553 14507 20587
rect 14749 20553 14783 20587
rect 2421 20485 2455 20519
rect 1409 20417 1443 20451
rect 2881 20417 2915 20451
rect 3065 20417 3099 20451
rect 5549 20417 5583 20451
rect 6009 20417 6043 20451
rect 6837 20417 6871 20451
rect 2329 20349 2363 20383
rect 4905 20349 4939 20383
rect 7104 20349 7138 20383
rect 9045 20349 9079 20383
rect 13093 20349 13127 20383
rect 2789 20281 2823 20315
rect 5457 20281 5491 20315
rect 9312 20281 9346 20315
rect 11253 20281 11287 20315
rect 12265 20281 12299 20315
rect 13338 20281 13372 20315
rect 1961 20213 1995 20247
rect 3525 20213 3559 20247
rect 3893 20213 3927 20247
rect 3985 20213 4019 20247
rect 4997 20213 5031 20247
rect 5365 20213 5399 20247
rect 10701 20213 10735 20247
rect 15301 20213 15335 20247
rect 2329 20009 2363 20043
rect 4721 20009 4755 20043
rect 6929 20009 6963 20043
rect 8033 20009 8067 20043
rect 8493 20009 8527 20043
rect 9137 20009 9171 20043
rect 11069 20009 11103 20043
rect 11713 20009 11747 20043
rect 13369 20009 13403 20043
rect 5448 19941 5482 19975
rect 9956 19941 9990 19975
rect 11345 19941 11379 19975
rect 15577 19941 15611 19975
rect 2697 19873 2731 19907
rect 4077 19873 4111 19907
rect 7573 19873 7607 19907
rect 8401 19873 8435 19907
rect 13277 19873 13311 19907
rect 15301 19873 15335 19907
rect 2789 19805 2823 19839
rect 2881 19805 2915 19839
rect 3893 19805 3927 19839
rect 5181 19805 5215 19839
rect 8677 19805 8711 19839
rect 9689 19805 9723 19839
rect 11897 19805 11931 19839
rect 13461 19805 13495 19839
rect 4997 19737 5031 19771
rect 7389 19737 7423 19771
rect 12909 19737 12943 19771
rect 14657 19737 14691 19771
rect 1685 19669 1719 19703
rect 2237 19669 2271 19703
rect 3433 19669 3467 19703
rect 4261 19669 4295 19703
rect 6561 19669 6595 19703
rect 7297 19669 7331 19703
rect 7941 19669 7975 19703
rect 9413 19669 9447 19703
rect 12449 19669 12483 19703
rect 13921 19669 13955 19703
rect 5641 19465 5675 19499
rect 8401 19465 8435 19499
rect 8953 19465 8987 19499
rect 13829 19465 13863 19499
rect 15669 19465 15703 19499
rect 5089 19329 5123 19363
rect 5273 19329 5307 19363
rect 7297 19329 7331 19363
rect 7389 19329 7423 19363
rect 9597 19329 9631 19363
rect 11253 19329 11287 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 2329 19261 2363 19295
rect 4169 19261 4203 19295
rect 4537 19261 4571 19295
rect 8125 19261 8159 19295
rect 8585 19261 8619 19295
rect 9413 19261 9447 19295
rect 10057 19261 10091 19295
rect 11621 19261 11655 19295
rect 12265 19261 12299 19295
rect 12449 19261 12483 19295
rect 14473 19261 14507 19295
rect 15025 19261 15059 19295
rect 2574 19193 2608 19227
rect 4997 19193 5031 19227
rect 6285 19193 6319 19227
rect 10425 19193 10459 19227
rect 12694 19193 12728 19227
rect 1869 19125 1903 19159
rect 2145 19125 2179 19159
rect 3709 19125 3743 19159
rect 4629 19125 4663 19159
rect 6561 19125 6595 19159
rect 6837 19125 6871 19159
rect 7205 19125 7239 19159
rect 9045 19125 9079 19159
rect 9505 19125 9539 19159
rect 10609 19125 10643 19159
rect 10977 19125 11011 19159
rect 11069 19125 11103 19159
rect 14105 19125 14139 19159
rect 14657 19125 14691 19159
rect 2329 18921 2363 18955
rect 2421 18921 2455 18955
rect 4721 18921 4755 18955
rect 7573 18921 7607 18955
rect 8125 18921 8159 18955
rect 9137 18921 9171 18955
rect 11897 18921 11931 18955
rect 12541 18921 12575 18955
rect 13185 18921 13219 18955
rect 13829 18921 13863 18955
rect 14657 18921 14691 18955
rect 2789 18853 2823 18887
rect 5816 18853 5850 18887
rect 9965 18853 9999 18887
rect 10333 18853 10367 18887
rect 13093 18853 13127 18887
rect 2881 18785 2915 18819
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 5457 18785 5491 18819
rect 5549 18785 5583 18819
rect 8309 18785 8343 18819
rect 10784 18785 10818 18819
rect 1409 18717 1443 18751
rect 2973 18717 3007 18751
rect 8493 18717 8527 18751
rect 10517 18717 10551 18751
rect 13277 18717 13311 18751
rect 5273 18649 5307 18683
rect 1869 18581 1903 18615
rect 3433 18581 3467 18615
rect 3801 18581 3835 18615
rect 4261 18581 4295 18615
rect 6929 18581 6963 18615
rect 7297 18581 7331 18615
rect 9505 18581 9539 18615
rect 12725 18581 12759 18615
rect 3341 18377 3375 18411
rect 6837 18377 6871 18411
rect 7941 18377 7975 18411
rect 8401 18377 8435 18411
rect 10793 18377 10827 18411
rect 14289 18377 14323 18411
rect 5273 18309 5307 18343
rect 10425 18309 10459 18343
rect 12265 18309 12299 18343
rect 12817 18309 12851 18343
rect 5641 18241 5675 18275
rect 7389 18241 7423 18275
rect 8953 18241 8987 18275
rect 10057 18241 10091 18275
rect 11345 18241 11379 18275
rect 1685 18173 1719 18207
rect 3893 18173 3927 18207
rect 8769 18173 8803 18207
rect 9413 18173 9447 18207
rect 10701 18173 10735 18207
rect 11253 18173 11287 18207
rect 12909 18173 12943 18207
rect 1952 18105 1986 18139
rect 3709 18105 3743 18139
rect 4160 18105 4194 18139
rect 6285 18105 6319 18139
rect 7297 18105 7331 18139
rect 11897 18105 11931 18139
rect 13176 18105 13210 18139
rect 3065 18037 3099 18071
rect 6561 18037 6595 18071
rect 7205 18037 7239 18071
rect 8309 18037 8343 18071
rect 8861 18037 8895 18071
rect 10517 18037 10551 18071
rect 11161 18037 11195 18071
rect 14565 18037 14599 18071
rect 2421 17833 2455 17867
rect 2881 17833 2915 17867
rect 4261 17833 4295 17867
rect 4629 17833 4663 17867
rect 5825 17833 5859 17867
rect 11161 17833 11195 17867
rect 11529 17833 11563 17867
rect 13001 17833 13035 17867
rect 13277 17833 13311 17867
rect 13737 17833 13771 17867
rect 5181 17765 5215 17799
rect 7174 17765 7208 17799
rect 2789 17697 2823 17731
rect 4077 17697 4111 17731
rect 5733 17697 5767 17731
rect 9505 17697 9539 17731
rect 10425 17697 10459 17731
rect 11877 17697 11911 17731
rect 13829 17697 13863 17731
rect 1409 17629 1443 17663
rect 2973 17629 3007 17663
rect 3893 17629 3927 17663
rect 6009 17629 6043 17663
rect 6929 17629 6963 17663
rect 10517 17629 10551 17663
rect 10701 17629 10735 17663
rect 11621 17629 11655 17663
rect 14013 17629 14047 17663
rect 1961 17561 1995 17595
rect 2329 17561 2363 17595
rect 3525 17561 3559 17595
rect 10057 17561 10091 17595
rect 5365 17493 5399 17527
rect 6469 17493 6503 17527
rect 6837 17493 6871 17527
rect 8309 17493 8343 17527
rect 8585 17493 8619 17527
rect 9045 17493 9079 17527
rect 9965 17493 9999 17527
rect 1593 17289 1627 17323
rect 2421 17289 2455 17323
rect 4169 17289 4203 17323
rect 6285 17289 6319 17323
rect 9321 17289 9355 17323
rect 11437 17289 11471 17323
rect 11713 17289 11747 17323
rect 12081 17289 12115 17323
rect 13093 17289 13127 17323
rect 7481 17221 7515 17255
rect 4721 17153 4755 17187
rect 5825 17153 5859 17187
rect 10057 17153 10091 17187
rect 1409 17085 1443 17119
rect 2513 17085 2547 17119
rect 4997 17085 5031 17119
rect 5549 17085 5583 17119
rect 10313 17085 10347 17119
rect 13553 17085 13587 17119
rect 2780 17017 2814 17051
rect 5641 17017 5675 17051
rect 8033 17017 8067 17051
rect 13820 17017 13854 17051
rect 2053 16949 2087 16983
rect 3893 16949 3927 16983
rect 5181 16949 5215 16983
rect 6561 16949 6595 16983
rect 7021 16949 7055 16983
rect 7849 16949 7883 16983
rect 12725 16949 12759 16983
rect 13461 16949 13495 16983
rect 14933 16949 14967 16983
rect 15209 16949 15243 16983
rect 2053 16745 2087 16779
rect 2789 16745 2823 16779
rect 3525 16745 3559 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 6285 16745 6319 16779
rect 9505 16745 9539 16779
rect 9965 16745 9999 16779
rect 11621 16745 11655 16779
rect 11989 16745 12023 16779
rect 13185 16745 13219 16779
rect 13645 16745 13679 16779
rect 14657 16745 14691 16779
rect 4537 16677 4571 16711
rect 5273 16677 5307 16711
rect 6377 16677 6411 16711
rect 6929 16677 6963 16711
rect 14197 16677 14231 16711
rect 15577 16677 15611 16711
rect 3801 16609 3835 16643
rect 5641 16609 5675 16643
rect 7113 16609 7147 16643
rect 7665 16609 7699 16643
rect 7921 16609 7955 16643
rect 10333 16609 10367 16643
rect 12633 16609 12667 16643
rect 13553 16609 13587 16643
rect 15301 16609 15335 16643
rect 2145 16541 2179 16575
rect 2329 16541 2363 16575
rect 4721 16541 4755 16575
rect 6469 16541 6503 16575
rect 7297 16541 7331 16575
rect 10425 16541 10459 16575
rect 10517 16541 10551 16575
rect 12081 16541 12115 16575
rect 12173 16541 12207 16575
rect 13737 16541 13771 16575
rect 1685 16473 1719 16507
rect 5917 16473 5951 16507
rect 3157 16405 3191 16439
rect 9045 16405 9079 16439
rect 11069 16405 11103 16439
rect 11345 16405 11379 16439
rect 13093 16405 13127 16439
rect 2605 16201 2639 16235
rect 4537 16201 4571 16235
rect 5641 16201 5675 16235
rect 6285 16201 6319 16235
rect 8585 16201 8619 16235
rect 10333 16201 10367 16235
rect 11897 16201 11931 16235
rect 12265 16201 12299 16235
rect 14381 16201 14415 16235
rect 4813 16133 4847 16167
rect 9965 16133 9999 16167
rect 2053 16065 2087 16099
rect 2237 16065 2271 16099
rect 2973 16065 3007 16099
rect 5181 16065 5215 16099
rect 5733 16065 5767 16099
rect 9321 16065 9355 16099
rect 11345 16065 11379 16099
rect 15761 16065 15795 16099
rect 3157 15997 3191 16031
rect 3424 15997 3458 16031
rect 6929 15997 6963 16031
rect 9137 15997 9171 16031
rect 10701 15997 10735 16031
rect 11253 15997 11287 16031
rect 13001 15997 13035 16031
rect 14657 15997 14691 16031
rect 15301 15997 15335 16031
rect 15485 15997 15519 16031
rect 16221 15997 16255 16031
rect 7174 15929 7208 15963
rect 11161 15929 11195 15963
rect 13268 15929 13302 15963
rect 1593 15861 1627 15895
rect 1961 15861 1995 15895
rect 6653 15861 6687 15895
rect 8309 15861 8343 15895
rect 9045 15861 9079 15895
rect 10517 15861 10551 15895
rect 10793 15861 10827 15895
rect 12909 15861 12943 15895
rect 2329 15657 2363 15691
rect 3801 15657 3835 15691
rect 4445 15657 4479 15691
rect 5089 15657 5123 15691
rect 7757 15657 7791 15691
rect 8125 15657 8159 15691
rect 9505 15657 9539 15691
rect 9873 15657 9907 15691
rect 10333 15657 10367 15691
rect 10885 15657 10919 15691
rect 12265 15657 12299 15691
rect 13829 15657 13863 15691
rect 3433 15589 3467 15623
rect 11989 15589 12023 15623
rect 16405 15589 16439 15623
rect 2789 15521 2823 15555
rect 5733 15521 5767 15555
rect 6000 15521 6034 15555
rect 8309 15521 8343 15555
rect 11253 15521 11287 15555
rect 12705 15521 12739 15555
rect 16129 15521 16163 15555
rect 1409 15453 1443 15487
rect 1869 15453 1903 15487
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 4537 15453 4571 15487
rect 4629 15453 4663 15487
rect 8493 15453 8527 15487
rect 11345 15453 11379 15487
rect 11529 15453 11563 15487
rect 12449 15453 12483 15487
rect 4077 15385 4111 15419
rect 10793 15385 10827 15419
rect 2421 15317 2455 15351
rect 5549 15317 5583 15351
rect 7113 15317 7147 15351
rect 9137 15317 9171 15351
rect 14197 15317 14231 15351
rect 1593 15113 1627 15147
rect 2789 15113 2823 15147
rect 9045 15113 9079 15147
rect 10701 15113 10735 15147
rect 10793 15113 10827 15147
rect 13829 15113 13863 15147
rect 14105 15113 14139 15147
rect 14473 15113 14507 15147
rect 8585 15045 8619 15079
rect 16129 15045 16163 15079
rect 3249 14977 3283 15011
rect 3433 14977 3467 15011
rect 4445 14977 4479 15011
rect 8953 14977 8987 15011
rect 9597 14977 9631 15011
rect 11437 14977 11471 15011
rect 1409 14909 1443 14943
rect 3157 14909 3191 14943
rect 4712 14909 4746 14943
rect 6837 14909 6871 14943
rect 9413 14909 9447 14943
rect 12449 14909 12483 14943
rect 2145 14841 2179 14875
rect 6653 14841 6687 14875
rect 7104 14841 7138 14875
rect 12265 14841 12299 14875
rect 12694 14841 12728 14875
rect 2421 14773 2455 14807
rect 4169 14773 4203 14807
rect 5825 14773 5859 14807
rect 6193 14773 6227 14807
rect 8217 14773 8251 14807
rect 9505 14773 9539 14807
rect 10241 14773 10275 14807
rect 11161 14773 11195 14807
rect 11253 14773 11287 14807
rect 11897 14773 11931 14807
rect 3157 14569 3191 14603
rect 3525 14569 3559 14603
rect 3709 14569 3743 14603
rect 4077 14569 4111 14603
rect 4445 14569 4479 14603
rect 5733 14569 5767 14603
rect 6101 14569 6135 14603
rect 7757 14569 7791 14603
rect 8033 14569 8067 14603
rect 9137 14569 9171 14603
rect 11069 14569 11103 14603
rect 11437 14569 11471 14603
rect 13277 14569 13311 14603
rect 14105 14569 14139 14603
rect 6561 14501 6595 14535
rect 12142 14501 12176 14535
rect 13645 14501 13679 14535
rect 14013 14501 14047 14535
rect 1409 14433 1443 14467
rect 1676 14433 1710 14467
rect 3893 14433 3927 14467
rect 4537 14433 4571 14467
rect 5917 14433 5951 14467
rect 6101 14433 6135 14467
rect 7941 14433 7975 14467
rect 8401 14433 8435 14467
rect 9945 14433 9979 14467
rect 4629 14365 4663 14399
rect 5641 14365 5675 14399
rect 6653 14365 6687 14399
rect 6745 14365 6779 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 9689 14365 9723 14399
rect 11897 14365 11931 14399
rect 2789 14297 2823 14331
rect 7573 14297 7607 14331
rect 5273 14229 5307 14263
rect 6193 14229 6227 14263
rect 7297 14229 7331 14263
rect 9413 14229 9447 14263
rect 11713 14229 11747 14263
rect 3709 14025 3743 14059
rect 4353 14025 4387 14059
rect 4629 14025 4663 14059
rect 6285 14025 6319 14059
rect 8125 14025 8159 14059
rect 8769 14025 8803 14059
rect 11161 14025 11195 14059
rect 12449 14025 12483 14059
rect 13553 14025 13587 14059
rect 3341 13957 3375 13991
rect 6561 13957 6595 13991
rect 6837 13957 6871 13991
rect 11805 13957 11839 13991
rect 5641 13889 5675 13923
rect 5733 13889 5767 13923
rect 7389 13889 7423 13923
rect 9045 13889 9079 13923
rect 12265 13889 12299 13923
rect 12909 13889 12943 13923
rect 13093 13889 13127 13923
rect 14289 13889 14323 13923
rect 16957 13889 16991 13923
rect 1593 13821 1627 13855
rect 5089 13821 5123 13855
rect 7297 13821 7331 13855
rect 8953 13821 8987 13855
rect 14013 13821 14047 13855
rect 14749 13821 14783 13855
rect 16681 13821 16715 13855
rect 17417 13821 17451 13855
rect 1860 13753 1894 13787
rect 7205 13753 7239 13787
rect 8677 13753 8711 13787
rect 9312 13753 9346 13787
rect 12817 13753 12851 13787
rect 2973 13685 3007 13719
rect 3801 13685 3835 13719
rect 5181 13685 5215 13719
rect 5549 13685 5583 13719
rect 10425 13685 10459 13719
rect 10701 13685 10735 13719
rect 11253 13685 11287 13719
rect 2513 13481 2547 13515
rect 3893 13481 3927 13515
rect 4537 13481 4571 13515
rect 5273 13481 5307 13515
rect 5733 13481 5767 13515
rect 6193 13481 6227 13515
rect 6929 13481 6963 13515
rect 8677 13481 8711 13515
rect 9689 13481 9723 13515
rect 10057 13481 10091 13515
rect 11989 13481 12023 13515
rect 12541 13481 12575 13515
rect 12909 13481 12943 13515
rect 2881 13413 2915 13447
rect 3525 13413 3559 13447
rect 9413 13413 9447 13447
rect 10149 13413 10183 13447
rect 17693 13413 17727 13447
rect 1777 13345 1811 13379
rect 6101 13345 6135 13379
rect 7665 13345 7699 13379
rect 8401 13345 8435 13379
rect 17417 13345 17451 13379
rect 1869 13277 1903 13311
rect 1961 13277 1995 13311
rect 2973 13277 3007 13311
rect 4629 13277 4663 13311
rect 4813 13277 4847 13311
rect 6377 13277 6411 13311
rect 7757 13277 7791 13311
rect 7849 13277 7883 13311
rect 10241 13277 10275 13311
rect 11529 13277 11563 13311
rect 1409 13209 1443 13243
rect 4169 13209 4203 13243
rect 7297 13209 7331 13243
rect 9137 13209 9171 13243
rect 5549 13141 5583 13175
rect 10701 13141 10735 13175
rect 11161 13141 11195 13175
rect 1593 12937 1627 12971
rect 1961 12937 1995 12971
rect 4721 12937 4755 12971
rect 5181 12937 5215 12971
rect 6561 12937 6595 12971
rect 9045 12937 9079 12971
rect 10057 12937 10091 12971
rect 11713 12937 11747 12971
rect 14565 12937 14599 12971
rect 17417 12937 17451 12971
rect 4813 12869 4847 12903
rect 6285 12869 6319 12903
rect 8217 12869 8251 12903
rect 13829 12869 13863 12903
rect 2513 12801 2547 12835
rect 5733 12801 5767 12835
rect 9597 12801 9631 12835
rect 11161 12801 11195 12835
rect 1409 12733 1443 12767
rect 2780 12733 2814 12767
rect 4261 12733 4295 12767
rect 4997 12733 5031 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 7093 12733 7127 12767
rect 8861 12733 8895 12767
rect 9505 12733 9539 12767
rect 11069 12733 11103 12767
rect 12449 12733 12483 12767
rect 14657 12733 14691 12767
rect 14913 12733 14947 12767
rect 5549 12665 5583 12699
rect 8493 12665 8527 12699
rect 9413 12665 9447 12699
rect 10517 12665 10551 12699
rect 10977 12665 11011 12699
rect 12265 12665 12299 12699
rect 12694 12665 12728 12699
rect 2421 12597 2455 12631
rect 3893 12597 3927 12631
rect 10609 12597 10643 12631
rect 16037 12597 16071 12631
rect 3893 12393 3927 12427
rect 4537 12393 4571 12427
rect 6009 12393 6043 12427
rect 7481 12393 7515 12427
rect 7757 12393 7791 12427
rect 9413 12393 9447 12427
rect 9965 12393 9999 12427
rect 10241 12393 10275 12427
rect 12265 12393 12299 12427
rect 13461 12393 13495 12427
rect 14657 12393 14691 12427
rect 4997 12325 5031 12359
rect 8309 12325 8343 12359
rect 11152 12325 11186 12359
rect 13553 12325 13587 12359
rect 21189 12325 21223 12359
rect 2044 12257 2078 12291
rect 4905 12257 4939 12291
rect 5641 12257 5675 12291
rect 6368 12257 6402 12291
rect 10609 12257 10643 12291
rect 20913 12257 20947 12291
rect 1777 12189 1811 12223
rect 4353 12189 4387 12223
rect 5181 12189 5215 12223
rect 6101 12189 6135 12223
rect 10885 12189 10919 12223
rect 12633 12189 12667 12223
rect 13645 12189 13679 12223
rect 3433 12121 3467 12155
rect 8125 12121 8159 12155
rect 1685 12053 1719 12087
rect 3157 12053 3191 12087
rect 9045 12053 9079 12087
rect 10425 12053 10459 12087
rect 13093 12053 13127 12087
rect 5181 11849 5215 11883
rect 6285 11849 6319 11883
rect 8125 11849 8159 11883
rect 9321 11849 9355 11883
rect 11253 11849 11287 11883
rect 11529 11849 11563 11883
rect 11897 11849 11931 11883
rect 13093 11849 13127 11883
rect 13461 11849 13495 11883
rect 13829 11849 13863 11883
rect 4997 11781 5031 11815
rect 6377 11781 6411 11815
rect 7757 11781 7791 11815
rect 1961 11713 1995 11747
rect 2513 11713 2547 11747
rect 2973 11713 3007 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 6837 11713 6871 11747
rect 7481 11713 7515 11747
rect 8861 11713 8895 11747
rect 9873 11713 9907 11747
rect 18337 11713 18371 11747
rect 1869 11645 1903 11679
rect 5549 11645 5583 11679
rect 6377 11645 6411 11679
rect 6653 11645 6687 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 18061 11645 18095 11679
rect 18797 11645 18831 11679
rect 2881 11577 2915 11611
rect 3240 11577 3274 11611
rect 9781 11577 9815 11611
rect 10118 11577 10152 11611
rect 1409 11509 1443 11543
rect 1777 11509 1811 11543
rect 4353 11509 4387 11543
rect 4629 11509 4663 11543
rect 8309 11509 8343 11543
rect 20913 11509 20947 11543
rect 2881 11305 2915 11339
rect 4077 11305 4111 11339
rect 5273 11305 5307 11339
rect 5641 11305 5675 11339
rect 6745 11305 6779 11339
rect 11069 11305 11103 11339
rect 11345 11305 11379 11339
rect 1409 11169 1443 11203
rect 1676 11169 1710 11203
rect 3065 11237 3099 11271
rect 9934 11237 9968 11271
rect 19809 11237 19843 11271
rect 4445 11169 4479 11203
rect 6009 11169 6043 11203
rect 8217 11169 8251 11203
rect 8953 11169 8987 11203
rect 9505 11169 9539 11203
rect 9689 11169 9723 11203
rect 19533 11169 19567 11203
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 8309 11101 8343 11135
rect 8493 11101 8527 11135
rect 2789 11033 2823 11067
rect 2881 11033 2915 11067
rect 3433 11033 3467 11067
rect 7021 11033 7055 11067
rect 7389 11033 7423 11067
rect 7849 11033 7883 11067
rect 3893 10965 3927 10999
rect 3893 10761 3927 10795
rect 7113 10761 7147 10795
rect 7941 10761 7975 10795
rect 9597 10761 9631 10795
rect 19533 10761 19567 10795
rect 10425 10693 10459 10727
rect 1961 10625 1995 10659
rect 2145 10625 2179 10659
rect 7205 10625 7239 10659
rect 10977 10625 11011 10659
rect 11437 10625 11471 10659
rect 18613 10625 18647 10659
rect 19901 10625 19935 10659
rect 3249 10557 3283 10591
rect 3985 10557 4019 10591
rect 8217 10557 8251 10591
rect 8484 10557 8518 10591
rect 10241 10557 10275 10591
rect 10885 10557 10919 10591
rect 18337 10557 18371 10591
rect 19073 10557 19107 10591
rect 19625 10557 19659 10591
rect 20361 10557 20395 10591
rect 2513 10489 2547 10523
rect 4230 10489 4264 10523
rect 6377 10489 6411 10523
rect 10793 10489 10827 10523
rect 1501 10421 1535 10455
rect 1869 10421 1903 10455
rect 2973 10421 3007 10455
rect 5365 10421 5399 10455
rect 5641 10421 5675 10455
rect 6101 10421 6135 10455
rect 9873 10421 9907 10455
rect 2789 10217 2823 10251
rect 3525 10217 3559 10251
rect 4077 10217 4111 10251
rect 4537 10217 4571 10251
rect 5089 10217 5123 10251
rect 5457 10217 5491 10251
rect 7941 10217 7975 10251
rect 8309 10217 8343 10251
rect 8585 10217 8619 10251
rect 10057 10217 10091 10251
rect 10701 10217 10735 10251
rect 3065 10149 3099 10183
rect 6254 10149 6288 10183
rect 9505 10149 9539 10183
rect 10149 10149 10183 10183
rect 1676 10081 1710 10115
rect 4445 10081 4479 10115
rect 1409 10013 1443 10047
rect 4721 10013 4755 10047
rect 6009 10013 6043 10047
rect 10241 10013 10275 10047
rect 9689 9945 9723 9979
rect 3893 9877 3927 9911
rect 5825 9877 5859 9911
rect 7389 9877 7423 9911
rect 1777 9673 1811 9707
rect 5457 9673 5491 9707
rect 6469 9673 6503 9707
rect 8493 9673 8527 9707
rect 9781 9673 9815 9707
rect 10425 9673 10459 9707
rect 3617 9605 3651 9639
rect 5733 9605 5767 9639
rect 3893 9537 3927 9571
rect 7113 9537 7147 9571
rect 10057 9537 10091 9571
rect 1869 9469 1903 9503
rect 2125 9469 2159 9503
rect 4077 9469 4111 9503
rect 4344 9469 4378 9503
rect 8769 9469 8803 9503
rect 7380 9401 7414 9435
rect 3249 9333 3283 9367
rect 6193 9333 6227 9367
rect 1685 9129 1719 9163
rect 1961 9129 1995 9163
rect 2605 9129 2639 9163
rect 3249 9129 3283 9163
rect 4077 9129 4111 9163
rect 4813 9129 4847 9163
rect 6469 9129 6503 9163
rect 7297 9129 7331 9163
rect 7757 9129 7791 9163
rect 2513 9061 2547 9095
rect 3893 9061 3927 9095
rect 5356 9061 5390 9095
rect 6745 9061 6779 9095
rect 7665 9061 7699 9095
rect 5089 8993 5123 9027
rect 2697 8925 2731 8959
rect 7941 8925 7975 8959
rect 7205 8857 7239 8891
rect 2145 8789 2179 8823
rect 2237 8585 2271 8619
rect 2605 8585 2639 8619
rect 2973 8585 3007 8619
rect 4537 8585 4571 8619
rect 4721 8585 4755 8619
rect 7757 8585 7791 8619
rect 8033 8585 8067 8619
rect 7389 8517 7423 8551
rect 1593 8449 1627 8483
rect 3433 8449 3467 8483
rect 3617 8449 3651 8483
rect 4261 8449 4295 8483
rect 5365 8449 5399 8483
rect 5733 8449 5767 8483
rect 3341 8381 3375 8415
rect 5089 8381 5123 8415
rect 5181 8381 5215 8415
rect 1685 8041 1719 8075
rect 2237 8041 2271 8075
rect 2881 8041 2915 8075
rect 3801 8041 3835 8075
rect 4537 8041 4571 8075
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 5733 8041 5767 8075
rect 4445 7973 4479 8007
rect 2789 7905 2823 7939
rect 3525 7905 3559 7939
rect 3065 7837 3099 7871
rect 4629 7837 4663 7871
rect 4077 7769 4111 7803
rect 2421 7701 2455 7735
rect 1685 7497 1719 7531
rect 1961 7497 1995 7531
rect 2513 7497 2547 7531
rect 2881 7497 2915 7531
rect 3157 7497 3191 7531
rect 4169 7497 4203 7531
rect 4537 7497 4571 7531
rect 22385 7497 22419 7531
rect 4813 7429 4847 7463
rect 22201 7293 22235 7327
rect 22753 7293 22787 7327
rect 22753 6817 22787 6851
rect 22937 6681 22971 6715
rect 22753 6409 22787 6443
rect 23857 6409 23891 6443
rect 23673 6205 23707 6239
rect 24225 6205 24259 6239
rect 24133 5865 24167 5899
rect 23949 5729 23983 5763
rect 23949 5321 23983 5355
rect 24685 5321 24719 5355
rect 24501 5117 24535 5151
rect 25053 5117 25087 5151
rect 24777 4777 24811 4811
rect 24593 4641 24627 4675
rect 24685 4233 24719 4267
<< metal1 >>
rect 4062 26800 4068 26852
rect 4120 26840 4126 26852
rect 7374 26840 7380 26852
rect 4120 26812 7380 26840
rect 4120 26800 4126 26812
rect 7374 26800 7380 26812
rect 7432 26800 7438 26852
rect 4062 26392 4068 26444
rect 4120 26432 4126 26444
rect 12066 26432 12072 26444
rect 4120 26404 12072 26432
rect 4120 26392 4126 26404
rect 12066 26392 12072 26404
rect 12124 26392 12130 26444
rect 3510 26324 3516 26376
rect 3568 26364 3574 26376
rect 11146 26364 11152 26376
rect 3568 26336 11152 26364
rect 3568 26324 3574 26336
rect 11146 26324 11152 26336
rect 11204 26324 11210 26376
rect 2038 25712 2044 25764
rect 2096 25752 2102 25764
rect 8478 25752 8484 25764
rect 2096 25724 8484 25752
rect 2096 25712 2102 25724
rect 8478 25712 8484 25724
rect 8536 25712 8542 25764
rect 3510 25644 3516 25696
rect 3568 25684 3574 25696
rect 13630 25684 13636 25696
rect 3568 25656 13636 25684
rect 3568 25644 3574 25656
rect 13630 25644 13636 25656
rect 13688 25644 13694 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 5629 25483 5687 25489
rect 5629 25449 5641 25483
rect 5675 25480 5687 25483
rect 6178 25480 6184 25492
rect 5675 25452 6184 25480
rect 5675 25449 5687 25452
rect 5629 25443 5687 25449
rect 6178 25440 6184 25452
rect 6236 25440 6242 25492
rect 6638 25440 6644 25492
rect 6696 25480 6702 25492
rect 7377 25483 7435 25489
rect 7377 25480 7389 25483
rect 6696 25452 7389 25480
rect 6696 25440 6702 25452
rect 7377 25449 7389 25452
rect 7423 25480 7435 25483
rect 8202 25480 8208 25492
rect 7423 25452 8208 25480
rect 7423 25449 7435 25452
rect 7377 25443 7435 25449
rect 8202 25440 8208 25452
rect 8260 25440 8266 25492
rect 8665 25483 8723 25489
rect 8665 25449 8677 25483
rect 8711 25449 8723 25483
rect 8665 25443 8723 25449
rect 11057 25483 11115 25489
rect 11057 25449 11069 25483
rect 11103 25480 11115 25483
rect 11146 25480 11152 25492
rect 11103 25452 11152 25480
rect 11103 25449 11115 25452
rect 11057 25443 11115 25449
rect 4062 25372 4068 25424
rect 4120 25412 4126 25424
rect 8680 25412 8708 25443
rect 11146 25440 11152 25452
rect 11204 25440 11210 25492
rect 13630 25480 13636 25492
rect 13591 25452 13636 25480
rect 13630 25440 13636 25452
rect 13688 25440 13694 25492
rect 4120 25384 8708 25412
rect 4120 25372 4126 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2314 25344 2320 25356
rect 1443 25316 2320 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2314 25304 2320 25316
rect 2372 25304 2378 25356
rect 2498 25344 2504 25356
rect 2459 25316 2504 25344
rect 2498 25304 2504 25316
rect 2556 25304 2562 25356
rect 4890 25344 4896 25356
rect 4851 25316 4896 25344
rect 4890 25304 4896 25316
rect 4948 25304 4954 25356
rect 4982 25304 4988 25356
rect 5040 25344 5046 25356
rect 5040 25316 5764 25344
rect 5040 25304 5046 25316
rect 4154 25236 4160 25288
rect 4212 25276 4218 25288
rect 5077 25279 5135 25285
rect 5077 25276 5089 25279
rect 4212 25248 5089 25276
rect 4212 25236 4218 25248
rect 5077 25245 5089 25248
rect 5123 25245 5135 25279
rect 5736 25276 5764 25316
rect 6914 25304 6920 25356
rect 6972 25344 6978 25356
rect 7285 25347 7343 25353
rect 7285 25344 7297 25347
rect 6972 25316 7297 25344
rect 6972 25304 6978 25316
rect 7285 25313 7297 25316
rect 7331 25313 7343 25347
rect 7650 25344 7656 25356
rect 7285 25307 7343 25313
rect 7392 25316 7656 25344
rect 7392 25276 7420 25316
rect 7650 25304 7656 25316
rect 7708 25304 7714 25356
rect 8478 25344 8484 25356
rect 8439 25316 8484 25344
rect 8478 25304 8484 25316
rect 8536 25304 8542 25356
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 9769 25347 9827 25353
rect 9769 25344 9781 25347
rect 9732 25316 9781 25344
rect 9732 25304 9738 25316
rect 9769 25313 9781 25316
rect 9815 25313 9827 25347
rect 9769 25307 9827 25313
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 10870 25344 10876 25356
rect 10100 25316 10876 25344
rect 10100 25304 10106 25316
rect 10870 25304 10876 25316
rect 10928 25304 10934 25356
rect 7558 25276 7564 25288
rect 5736 25248 7420 25276
rect 7519 25248 7564 25276
rect 5077 25239 5135 25245
rect 7558 25236 7564 25248
rect 7616 25236 7622 25288
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 12621 25279 12679 25285
rect 12621 25276 12633 25279
rect 12400 25248 12633 25276
rect 12400 25236 12406 25248
rect 12621 25245 12633 25248
rect 12667 25245 12679 25279
rect 12621 25239 12679 25245
rect 3237 25211 3295 25217
rect 3237 25177 3249 25211
rect 3283 25208 3295 25211
rect 4706 25208 4712 25220
rect 3283 25180 4712 25208
rect 3283 25177 3295 25180
rect 3237 25171 3295 25177
rect 4706 25168 4712 25180
rect 4764 25168 4770 25220
rect 5626 25168 5632 25220
rect 5684 25208 5690 25220
rect 5905 25211 5963 25217
rect 5905 25208 5917 25211
rect 5684 25180 5917 25208
rect 5684 25168 5690 25180
rect 5905 25177 5917 25180
rect 5951 25177 5963 25211
rect 5905 25171 5963 25177
rect 6733 25211 6791 25217
rect 6733 25177 6745 25211
rect 6779 25208 6791 25211
rect 7282 25208 7288 25220
rect 6779 25180 7288 25208
rect 6779 25177 6791 25180
rect 6733 25171 6791 25177
rect 7282 25168 7288 25180
rect 7340 25168 7346 25220
rect 7374 25168 7380 25220
rect 7432 25208 7438 25220
rect 9953 25211 10011 25217
rect 9953 25208 9965 25211
rect 7432 25180 9965 25208
rect 7432 25168 7438 25180
rect 9953 25177 9965 25180
rect 9999 25177 10011 25211
rect 9953 25171 10011 25177
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2774 25140 2780 25152
rect 2731 25112 2780 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 3602 25100 3608 25152
rect 3660 25140 3666 25152
rect 4525 25143 4583 25149
rect 4525 25140 4537 25143
rect 3660 25112 4537 25140
rect 3660 25100 3666 25112
rect 4525 25109 4537 25112
rect 4571 25109 4583 25143
rect 4525 25103 4583 25109
rect 5994 25100 6000 25152
rect 6052 25140 6058 25152
rect 6917 25143 6975 25149
rect 6917 25140 6929 25143
rect 6052 25112 6929 25140
rect 6052 25100 6058 25112
rect 6917 25109 6929 25112
rect 6963 25109 6975 25143
rect 6917 25103 6975 25109
rect 10413 25143 10471 25149
rect 10413 25109 10425 25143
rect 10459 25140 10471 25143
rect 10686 25140 10692 25152
rect 10459 25112 10692 25140
rect 10459 25109 10471 25112
rect 10413 25103 10471 25109
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 4617 24939 4675 24945
rect 4617 24905 4629 24939
rect 4663 24936 4675 24939
rect 4982 24936 4988 24948
rect 4663 24908 4988 24936
rect 4663 24905 4675 24908
rect 4617 24899 4675 24905
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 9674 24936 9680 24948
rect 9635 24908 9680 24936
rect 9674 24896 9680 24908
rect 9732 24896 9738 24948
rect 10870 24936 10876 24948
rect 10831 24908 10876 24936
rect 10870 24896 10876 24908
rect 10928 24896 10934 24948
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 8573 24871 8631 24877
rect 8573 24868 8585 24871
rect 4120 24840 8585 24868
rect 4120 24828 4126 24840
rect 8573 24837 8585 24840
rect 8619 24837 8631 24871
rect 10134 24868 10140 24880
rect 8573 24831 8631 24837
rect 9600 24840 10140 24868
rect 3602 24800 3608 24812
rect 3563 24772 3608 24800
rect 3602 24760 3608 24772
rect 3660 24760 3666 24812
rect 3789 24803 3847 24809
rect 3789 24769 3801 24803
rect 3835 24800 3847 24803
rect 4706 24800 4712 24812
rect 3835 24772 4712 24800
rect 3835 24769 3847 24772
rect 3789 24763 3847 24769
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 5074 24760 5080 24812
rect 5132 24800 5138 24812
rect 5534 24800 5540 24812
rect 5132 24772 5540 24800
rect 5132 24760 5138 24772
rect 5534 24760 5540 24772
rect 5592 24800 5598 24812
rect 5721 24803 5779 24809
rect 5721 24800 5733 24803
rect 5592 24772 5733 24800
rect 5592 24760 5598 24772
rect 5721 24769 5733 24772
rect 5767 24769 5779 24803
rect 6638 24800 6644 24812
rect 6599 24772 6644 24800
rect 5721 24763 5779 24769
rect 6638 24760 6644 24772
rect 6696 24760 6702 24812
rect 7282 24800 7288 24812
rect 7243 24772 7288 24800
rect 7282 24760 7288 24772
rect 7340 24760 7346 24812
rect 7466 24760 7472 24812
rect 7524 24800 7530 24812
rect 9033 24803 9091 24809
rect 7524 24772 7972 24800
rect 7524 24760 7530 24772
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 3053 24735 3111 24741
rect 1443 24704 1900 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1872 24608 1900 24704
rect 3053 24701 3065 24735
rect 3099 24732 3111 24735
rect 3510 24732 3516 24744
rect 3099 24704 3516 24732
rect 3099 24701 3111 24704
rect 3053 24695 3111 24701
rect 3510 24692 3516 24704
rect 3568 24692 3574 24744
rect 4614 24692 4620 24744
rect 4672 24732 4678 24744
rect 5629 24735 5687 24741
rect 5629 24732 5641 24735
rect 4672 24704 5641 24732
rect 4672 24692 4678 24704
rect 5629 24701 5641 24704
rect 5675 24732 5687 24735
rect 5994 24732 6000 24744
rect 5675 24704 6000 24732
rect 5675 24701 5687 24704
rect 5629 24695 5687 24701
rect 5994 24692 6000 24704
rect 6052 24692 6058 24744
rect 6273 24735 6331 24741
rect 6273 24701 6285 24735
rect 6319 24732 6331 24735
rect 6914 24732 6920 24744
rect 6319 24704 6920 24732
rect 6319 24701 6331 24704
rect 6273 24695 6331 24701
rect 6914 24692 6920 24704
rect 6972 24692 6978 24744
rect 2406 24624 2412 24676
rect 2464 24664 2470 24676
rect 7944 24673 7972 24772
rect 9033 24769 9045 24803
rect 9079 24800 9091 24803
rect 9600 24800 9628 24840
rect 10134 24828 10140 24840
rect 10192 24868 10198 24880
rect 10192 24840 10456 24868
rect 10192 24828 10198 24840
rect 10428 24809 10456 24840
rect 9079 24772 9628 24800
rect 10413 24803 10471 24809
rect 9079 24769 9091 24772
rect 9033 24763 9091 24769
rect 10413 24769 10425 24803
rect 10459 24769 10471 24803
rect 10413 24763 10471 24769
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12342 24800 12348 24812
rect 12299 24772 12348 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12342 24760 12348 24772
rect 12400 24800 12406 24812
rect 12618 24800 12624 24812
rect 12400 24772 12624 24800
rect 12400 24760 12406 24772
rect 12618 24760 12624 24772
rect 12676 24760 12682 24812
rect 12986 24800 12992 24812
rect 12947 24772 12992 24800
rect 12986 24760 12992 24772
rect 13044 24760 13050 24812
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13814 24800 13820 24812
rect 13412 24772 13820 24800
rect 13412 24760 13418 24772
rect 13814 24760 13820 24772
rect 13872 24760 13878 24812
rect 8389 24735 8447 24741
rect 8389 24701 8401 24735
rect 8435 24732 8447 24735
rect 8662 24732 8668 24744
rect 8435 24704 8668 24732
rect 8435 24701 8447 24704
rect 8389 24695 8447 24701
rect 8662 24692 8668 24704
rect 8720 24692 8726 24744
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24732 9459 24735
rect 9447 24704 10272 24732
rect 9447 24701 9459 24704
rect 9401 24695 9459 24701
rect 10244 24676 10272 24704
rect 7929 24667 7987 24673
rect 2464 24636 3188 24664
rect 2464 24624 2470 24636
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 1854 24556 1860 24608
rect 1912 24596 1918 24608
rect 1949 24599 2007 24605
rect 1949 24596 1961 24599
rect 1912 24568 1961 24596
rect 1912 24556 1918 24568
rect 1949 24565 1961 24568
rect 1995 24565 2007 24599
rect 2314 24596 2320 24608
rect 2227 24568 2320 24596
rect 1949 24559 2007 24565
rect 2314 24556 2320 24568
rect 2372 24596 2378 24608
rect 2682 24596 2688 24608
rect 2372 24568 2688 24596
rect 2372 24556 2378 24568
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 3160 24605 3188 24636
rect 7929 24633 7941 24667
rect 7975 24664 7987 24667
rect 8202 24664 8208 24676
rect 7975 24636 8208 24664
rect 7975 24633 7987 24636
rect 7929 24627 7987 24633
rect 8202 24624 8208 24636
rect 8260 24624 8266 24676
rect 9582 24624 9588 24676
rect 9640 24664 9646 24676
rect 10226 24664 10232 24676
rect 9640 24636 9904 24664
rect 10187 24636 10232 24664
rect 9640 24624 9646 24636
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24565 3203 24599
rect 4154 24596 4160 24608
rect 4115 24568 4160 24596
rect 3145 24559 3203 24565
rect 4154 24556 4160 24568
rect 4212 24556 4218 24608
rect 4890 24596 4896 24608
rect 4851 24568 4896 24596
rect 4890 24556 4896 24568
rect 4948 24556 4954 24608
rect 5166 24596 5172 24608
rect 5127 24568 5172 24596
rect 5166 24556 5172 24568
rect 5224 24556 5230 24608
rect 5537 24599 5595 24605
rect 5537 24565 5549 24599
rect 5583 24596 5595 24599
rect 5994 24596 6000 24608
rect 5583 24568 6000 24596
rect 5583 24565 5595 24568
rect 5537 24559 5595 24565
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 6822 24596 6828 24608
rect 6783 24568 6828 24596
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 6914 24556 6920 24608
rect 6972 24596 6978 24608
rect 7193 24599 7251 24605
rect 7193 24596 7205 24599
rect 6972 24568 7205 24596
rect 6972 24556 6978 24568
rect 7193 24565 7205 24568
rect 7239 24565 7251 24599
rect 7193 24559 7251 24565
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 8297 24599 8355 24605
rect 8297 24596 8309 24599
rect 7616 24568 8309 24596
rect 7616 24556 7622 24568
rect 8297 24565 8309 24568
rect 8343 24596 8355 24599
rect 8386 24596 8392 24608
rect 8343 24568 8392 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 9876 24605 9904 24636
rect 10226 24624 10232 24636
rect 10284 24624 10290 24676
rect 11885 24667 11943 24673
rect 11885 24633 11897 24667
rect 11931 24664 11943 24667
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 11931 24636 12909 24664
rect 11931 24633 11943 24636
rect 11885 24627 11943 24633
rect 12897 24633 12909 24636
rect 12943 24664 12955 24667
rect 13078 24664 13084 24676
rect 12943 24636 13084 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 13078 24624 13084 24636
rect 13136 24624 13142 24676
rect 13998 24664 14004 24676
rect 13959 24636 14004 24664
rect 13998 24624 14004 24636
rect 14056 24624 14062 24676
rect 9861 24599 9919 24605
rect 9861 24565 9873 24599
rect 9907 24565 9919 24599
rect 9861 24559 9919 24565
rect 10321 24599 10379 24605
rect 10321 24565 10333 24599
rect 10367 24596 10379 24599
rect 10686 24596 10692 24608
rect 10367 24568 10692 24596
rect 10367 24565 10379 24568
rect 10321 24559 10379 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 12158 24556 12164 24608
rect 12216 24596 12222 24608
rect 12437 24599 12495 24605
rect 12437 24596 12449 24599
rect 12216 24568 12449 24596
rect 12216 24556 12222 24568
rect 12437 24565 12449 24568
rect 12483 24565 12495 24599
rect 12437 24559 12495 24565
rect 12618 24556 12624 24608
rect 12676 24596 12682 24608
rect 12805 24599 12863 24605
rect 12805 24596 12817 24599
rect 12676 24568 12817 24596
rect 12676 24556 12682 24568
rect 12805 24565 12817 24568
rect 12851 24565 12863 24599
rect 12805 24559 12863 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 3421 24395 3479 24401
rect 3421 24361 3433 24395
rect 3467 24392 3479 24395
rect 3602 24392 3608 24404
rect 3467 24364 3608 24392
rect 3467 24361 3479 24364
rect 3421 24355 3479 24361
rect 3602 24352 3608 24364
rect 3660 24352 3666 24404
rect 4614 24392 4620 24404
rect 4575 24364 4620 24392
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 8478 24352 8484 24404
rect 8536 24392 8542 24404
rect 9033 24395 9091 24401
rect 9033 24392 9045 24395
rect 8536 24364 9045 24392
rect 8536 24352 8542 24364
rect 9033 24361 9045 24364
rect 9079 24361 9091 24395
rect 9033 24355 9091 24361
rect 10686 24352 10692 24404
rect 10744 24392 10750 24404
rect 11517 24395 11575 24401
rect 11517 24392 11529 24395
rect 10744 24364 11529 24392
rect 10744 24352 10750 24364
rect 11517 24361 11529 24364
rect 11563 24361 11575 24395
rect 11517 24355 11575 24361
rect 11977 24395 12035 24401
rect 11977 24361 11989 24395
rect 12023 24392 12035 24395
rect 12250 24392 12256 24404
rect 12023 24364 12256 24392
rect 12023 24361 12035 24364
rect 11977 24355 12035 24361
rect 12250 24352 12256 24364
rect 12308 24352 12314 24404
rect 13078 24392 13084 24404
rect 13039 24364 13084 24392
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 16482 24392 16488 24404
rect 15519 24364 16488 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 16482 24352 16488 24364
rect 16540 24352 16546 24404
rect 16577 24395 16635 24401
rect 16577 24361 16589 24395
rect 16623 24392 16635 24395
rect 17862 24392 17868 24404
rect 16623 24364 17868 24392
rect 16623 24361 16635 24364
rect 16577 24355 16635 24361
rect 17862 24352 17868 24364
rect 17920 24352 17926 24404
rect 18966 24392 18972 24404
rect 18927 24364 18972 24392
rect 18966 24352 18972 24364
rect 19024 24352 19030 24404
rect 21085 24395 21143 24401
rect 21085 24361 21097 24395
rect 21131 24392 21143 24395
rect 22462 24392 22468 24404
rect 21131 24364 22468 24392
rect 21131 24361 21143 24364
rect 21085 24355 21143 24361
rect 22462 24352 22468 24364
rect 22520 24352 22526 24404
rect 4976 24327 5034 24333
rect 4976 24293 4988 24327
rect 5022 24324 5034 24327
rect 5074 24324 5080 24336
rect 5022 24296 5080 24324
rect 5022 24293 5034 24296
rect 4976 24287 5034 24293
rect 5074 24284 5080 24296
rect 5132 24284 5138 24336
rect 7276 24327 7334 24333
rect 7276 24293 7288 24327
rect 7322 24324 7334 24327
rect 7466 24324 7472 24336
rect 7322 24296 7472 24324
rect 7322 24293 7334 24296
rect 7276 24287 7334 24293
rect 7466 24284 7472 24296
rect 7524 24284 7530 24336
rect 9950 24284 9956 24336
rect 10008 24324 10014 24336
rect 10413 24327 10471 24333
rect 10413 24324 10425 24327
rect 10008 24296 10425 24324
rect 10008 24284 10014 24296
rect 10413 24293 10425 24296
rect 10459 24324 10471 24327
rect 11698 24324 11704 24336
rect 10459 24296 11704 24324
rect 10459 24293 10471 24296
rect 10413 24287 10471 24293
rect 11698 24284 11704 24296
rect 11756 24284 11762 24336
rect 12802 24284 12808 24336
rect 12860 24324 12866 24336
rect 13541 24327 13599 24333
rect 13541 24324 13553 24327
rect 12860 24296 13553 24324
rect 12860 24284 12866 24296
rect 13541 24293 13553 24296
rect 13587 24293 13599 24327
rect 13541 24287 13599 24293
rect 1489 24259 1547 24265
rect 1489 24225 1501 24259
rect 1535 24256 1547 24259
rect 2590 24256 2596 24268
rect 1535 24228 2596 24256
rect 1535 24225 1547 24228
rect 1489 24219 1547 24225
rect 2590 24216 2596 24228
rect 2648 24216 2654 24268
rect 2777 24259 2835 24265
rect 2777 24225 2789 24259
rect 2823 24256 2835 24259
rect 2866 24256 2872 24268
rect 2823 24228 2872 24256
rect 2823 24225 2835 24228
rect 2777 24219 2835 24225
rect 2866 24216 2872 24228
rect 2924 24216 2930 24268
rect 4062 24216 4068 24268
rect 4120 24256 4126 24268
rect 4709 24259 4767 24265
rect 4709 24256 4721 24259
rect 4120 24228 4721 24256
rect 4120 24216 4126 24228
rect 4709 24225 4721 24228
rect 4755 24256 4767 24259
rect 4755 24228 6592 24256
rect 4755 24225 4767 24228
rect 4709 24219 4767 24225
rect 1762 24188 1768 24200
rect 1723 24160 1768 24188
rect 1762 24148 1768 24160
rect 1820 24148 1826 24200
rect 6564 24197 6592 24228
rect 9306 24216 9312 24268
rect 9364 24256 9370 24268
rect 10321 24259 10379 24265
rect 10321 24256 10333 24259
rect 9364 24228 10333 24256
rect 9364 24216 9370 24228
rect 10321 24225 10333 24228
rect 10367 24225 10379 24259
rect 11882 24256 11888 24268
rect 11843 24228 11888 24256
rect 10321 24219 10379 24225
rect 11882 24216 11888 24228
rect 11940 24216 11946 24268
rect 11974 24216 11980 24268
rect 12032 24256 12038 24268
rect 13449 24259 13507 24265
rect 13449 24256 13461 24259
rect 12032 24228 13461 24256
rect 12032 24216 12038 24228
rect 13449 24225 13461 24228
rect 13495 24225 13507 24259
rect 13449 24219 13507 24225
rect 15289 24259 15347 24265
rect 15289 24225 15301 24259
rect 15335 24256 15347 24259
rect 16022 24256 16028 24268
rect 15335 24228 16028 24256
rect 15335 24225 15347 24228
rect 15289 24219 15347 24225
rect 16022 24216 16028 24228
rect 16080 24216 16086 24268
rect 16114 24216 16120 24268
rect 16172 24256 16178 24268
rect 16393 24259 16451 24265
rect 16393 24256 16405 24259
rect 16172 24228 16405 24256
rect 16172 24216 16178 24228
rect 16393 24225 16405 24228
rect 16439 24225 16451 24259
rect 17494 24256 17500 24268
rect 17455 24228 17500 24256
rect 16393 24219 16451 24225
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 18782 24256 18788 24268
rect 18743 24228 18788 24256
rect 18782 24216 18788 24228
rect 18840 24216 18846 24268
rect 20901 24259 20959 24265
rect 20901 24225 20913 24259
rect 20947 24256 20959 24259
rect 21174 24256 21180 24268
rect 20947 24228 21180 24256
rect 20947 24225 20959 24228
rect 20901 24219 20959 24225
rect 21174 24216 21180 24228
rect 21232 24216 21238 24268
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24188 6607 24191
rect 7006 24188 7012 24200
rect 6595 24160 7012 24188
rect 6595 24157 6607 24160
rect 6549 24151 6607 24157
rect 7006 24148 7012 24160
rect 7064 24148 7070 24200
rect 9493 24191 9551 24197
rect 9493 24157 9505 24191
rect 9539 24188 9551 24191
rect 10505 24191 10563 24197
rect 10505 24188 10517 24191
rect 9539 24160 10517 24188
rect 9539 24157 9551 24160
rect 9493 24151 9551 24157
rect 10505 24157 10517 24160
rect 10551 24188 10563 24191
rect 10962 24188 10968 24200
rect 10551 24160 10968 24188
rect 10551 24157 10563 24160
rect 10505 24151 10563 24157
rect 10962 24148 10968 24160
rect 11020 24148 11026 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24188 12219 24191
rect 12342 24188 12348 24200
rect 12207 24160 12348 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 13725 24191 13783 24197
rect 13725 24157 13737 24191
rect 13771 24188 13783 24191
rect 14550 24188 14556 24200
rect 13771 24160 14556 24188
rect 13771 24157 13783 24160
rect 13725 24151 13783 24157
rect 14550 24148 14556 24160
rect 14608 24148 14614 24200
rect 10042 24080 10048 24132
rect 10100 24120 10106 24132
rect 11057 24123 11115 24129
rect 11057 24120 11069 24123
rect 10100 24092 11069 24120
rect 10100 24080 10106 24092
rect 11057 24089 11069 24092
rect 11103 24120 11115 24123
rect 12894 24120 12900 24132
rect 11103 24092 12900 24120
rect 11103 24089 11115 24092
rect 11057 24083 11115 24089
rect 12894 24080 12900 24092
rect 12952 24080 12958 24132
rect 17678 24120 17684 24132
rect 17639 24092 17684 24120
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 1762 24012 1768 24064
rect 1820 24052 1826 24064
rect 2498 24052 2504 24064
rect 1820 24024 2504 24052
rect 1820 24012 1826 24024
rect 2498 24012 2504 24024
rect 2556 24012 2562 24064
rect 2958 24052 2964 24064
rect 2919 24024 2964 24052
rect 2958 24012 2964 24024
rect 3016 24012 3022 24064
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 6089 24055 6147 24061
rect 6089 24052 6101 24055
rect 4212 24024 6101 24052
rect 4212 24012 4218 24024
rect 6089 24021 6101 24024
rect 6135 24021 6147 24055
rect 6914 24052 6920 24064
rect 6875 24024 6920 24052
rect 6089 24015 6147 24021
rect 6914 24012 6920 24024
rect 6972 24012 6978 24064
rect 8386 24052 8392 24064
rect 8347 24024 8392 24052
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 9858 24012 9864 24064
rect 9916 24052 9922 24064
rect 9953 24055 10011 24061
rect 9953 24052 9965 24055
rect 9916 24024 9965 24052
rect 9916 24012 9922 24024
rect 9953 24021 9965 24024
rect 9999 24021 10011 24055
rect 9953 24015 10011 24021
rect 12621 24055 12679 24061
rect 12621 24021 12633 24055
rect 12667 24052 12679 24055
rect 12986 24052 12992 24064
rect 12667 24024 12992 24052
rect 12667 24021 12679 24024
rect 12621 24015 12679 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2498 23848 2504 23860
rect 2459 23820 2504 23848
rect 2498 23808 2504 23820
rect 2556 23808 2562 23860
rect 2866 23848 2872 23860
rect 2827 23820 2872 23848
rect 2866 23808 2872 23820
rect 2924 23808 2930 23860
rect 5350 23848 5356 23860
rect 5311 23820 5356 23848
rect 5350 23808 5356 23820
rect 5408 23808 5414 23860
rect 5534 23808 5540 23860
rect 5592 23848 5598 23860
rect 5721 23851 5779 23857
rect 5721 23848 5733 23851
rect 5592 23820 5733 23848
rect 5592 23808 5598 23820
rect 5721 23817 5733 23820
rect 5767 23817 5779 23851
rect 5721 23811 5779 23817
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 7466 23848 7472 23860
rect 6687 23820 7472 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 7466 23808 7472 23820
rect 7524 23808 7530 23860
rect 9950 23848 9956 23860
rect 9911 23820 9956 23848
rect 9950 23808 9956 23820
rect 10008 23808 10014 23860
rect 11793 23851 11851 23857
rect 11793 23817 11805 23851
rect 11839 23848 11851 23851
rect 12250 23848 12256 23860
rect 11839 23820 12256 23848
rect 11839 23817 11851 23820
rect 11793 23811 11851 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12802 23848 12808 23860
rect 12763 23820 12808 23848
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 14274 23848 14280 23860
rect 14235 23820 14280 23848
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 15289 23851 15347 23857
rect 15289 23817 15301 23851
rect 15335 23848 15347 23851
rect 16206 23848 16212 23860
rect 15335 23820 16212 23848
rect 15335 23817 15347 23820
rect 15289 23811 15347 23817
rect 16206 23808 16212 23820
rect 16264 23808 16270 23860
rect 16390 23848 16396 23860
rect 16351 23820 16396 23848
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19242 23848 19248 23860
rect 18279 23820 19248 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 20254 23848 20260 23860
rect 19383 23820 20260 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20438 23848 20444 23860
rect 20399 23820 20444 23848
rect 20438 23808 20444 23820
rect 20496 23808 20502 23860
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 23382 23848 23388 23860
rect 22695 23820 23388 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 23382 23808 23388 23820
rect 23440 23808 23446 23860
rect 5074 23780 5080 23792
rect 5035 23752 5080 23780
rect 5074 23740 5080 23752
rect 5132 23740 5138 23792
rect 8478 23780 8484 23792
rect 8439 23752 8484 23780
rect 8478 23740 8484 23752
rect 8536 23740 8542 23792
rect 11974 23740 11980 23792
rect 12032 23780 12038 23792
rect 12161 23783 12219 23789
rect 12161 23780 12173 23783
rect 12032 23752 12173 23780
rect 12032 23740 12038 23752
rect 12161 23749 12173 23752
rect 12207 23749 12219 23783
rect 12161 23743 12219 23749
rect 4614 23672 4620 23724
rect 4672 23712 4678 23724
rect 5258 23712 5264 23724
rect 4672 23684 5264 23712
rect 4672 23672 4678 23684
rect 5258 23672 5264 23684
rect 5316 23672 5322 23724
rect 9217 23715 9275 23721
rect 9217 23681 9229 23715
rect 9263 23712 9275 23715
rect 9263 23684 10180 23712
rect 9263 23681 9275 23684
rect 9217 23675 9275 23681
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23644 1731 23647
rect 2406 23644 2412 23656
rect 1719 23616 2412 23644
rect 1719 23613 1731 23616
rect 1673 23607 1731 23613
rect 2406 23604 2412 23616
rect 2464 23604 2470 23656
rect 3329 23647 3387 23653
rect 3329 23613 3341 23647
rect 3375 23644 3387 23647
rect 4062 23644 4068 23656
rect 3375 23616 4068 23644
rect 3375 23613 3387 23616
rect 3329 23607 3387 23613
rect 4062 23604 4068 23616
rect 4120 23604 4126 23656
rect 5350 23604 5356 23656
rect 5408 23644 5414 23656
rect 5537 23647 5595 23653
rect 5537 23644 5549 23647
rect 5408 23616 5549 23644
rect 5408 23604 5414 23616
rect 5537 23613 5549 23616
rect 5583 23613 5595 23647
rect 5537 23607 5595 23613
rect 7006 23604 7012 23656
rect 7064 23644 7070 23656
rect 7101 23647 7159 23653
rect 7101 23644 7113 23647
rect 7064 23616 7113 23644
rect 7064 23604 7070 23616
rect 7101 23613 7113 23616
rect 7147 23644 7159 23647
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 7147 23616 8769 23644
rect 7147 23613 7159 23616
rect 7101 23607 7159 23613
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 10042 23644 10048 23656
rect 10003 23616 10048 23644
rect 8757 23607 8815 23613
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 10152 23644 10180 23684
rect 10312 23647 10370 23653
rect 10312 23644 10324 23647
rect 10152 23616 10324 23644
rect 10312 23613 10324 23616
rect 10358 23644 10370 23647
rect 12342 23644 12348 23656
rect 10358 23616 12348 23644
rect 10358 23613 10370 23616
rect 10312 23607 10370 23613
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12894 23644 12900 23656
rect 12855 23616 12900 23644
rect 12894 23604 12900 23616
rect 12952 23604 12958 23656
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 15105 23647 15163 23653
rect 15105 23644 15117 23647
rect 14424 23616 15117 23644
rect 14424 23604 14430 23616
rect 15105 23613 15117 23616
rect 15151 23613 15163 23647
rect 15105 23607 15163 23613
rect 1946 23576 1952 23588
rect 1907 23548 1952 23576
rect 1946 23536 1952 23548
rect 2004 23536 2010 23588
rect 3237 23579 3295 23585
rect 3237 23545 3249 23579
rect 3283 23576 3295 23579
rect 3574 23579 3632 23585
rect 3574 23576 3586 23579
rect 3283 23548 3586 23576
rect 3283 23545 3295 23548
rect 3237 23539 3295 23545
rect 3574 23545 3586 23548
rect 3620 23576 3632 23579
rect 4154 23576 4160 23588
rect 3620 23548 4160 23576
rect 3620 23545 3632 23548
rect 3574 23539 3632 23545
rect 4154 23536 4160 23548
rect 4212 23536 4218 23588
rect 6273 23579 6331 23585
rect 6273 23545 6285 23579
rect 6319 23576 6331 23579
rect 7346 23579 7404 23585
rect 7346 23576 7358 23579
rect 6319 23548 7358 23576
rect 6319 23545 6331 23548
rect 6273 23539 6331 23545
rect 7346 23545 7358 23548
rect 7392 23576 7404 23579
rect 8386 23576 8392 23588
rect 7392 23548 8392 23576
rect 7392 23545 7404 23548
rect 7346 23539 7404 23545
rect 8386 23536 8392 23548
rect 8444 23536 8450 23588
rect 12986 23536 12992 23588
rect 13044 23576 13050 23588
rect 13164 23579 13222 23585
rect 13164 23576 13176 23579
rect 13044 23548 13176 23576
rect 13044 23536 13050 23548
rect 13164 23545 13176 23548
rect 13210 23576 13222 23579
rect 13722 23576 13728 23588
rect 13210 23548 13728 23576
rect 13210 23545 13222 23548
rect 13164 23539 13222 23545
rect 13722 23536 13728 23548
rect 13780 23536 13786 23588
rect 15120 23576 15148 23607
rect 15562 23604 15568 23656
rect 15620 23644 15626 23656
rect 16209 23647 16267 23653
rect 16209 23644 16221 23647
rect 15620 23616 16221 23644
rect 15620 23604 15626 23616
rect 16209 23613 16221 23616
rect 16255 23644 16267 23647
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16255 23616 16773 23644
rect 16255 23613 16267 23616
rect 16209 23607 16267 23613
rect 16761 23613 16773 23616
rect 16807 23613 16819 23647
rect 18046 23644 18052 23656
rect 18007 23616 18052 23644
rect 16761 23607 16819 23613
rect 18046 23604 18052 23616
rect 18104 23644 18110 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18104 23616 18613 23644
rect 18104 23604 18110 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18601 23607 18659 23613
rect 19153 23647 19211 23653
rect 19153 23613 19165 23647
rect 19199 23613 19211 23647
rect 19153 23607 19211 23613
rect 15657 23579 15715 23585
rect 15657 23576 15669 23579
rect 15120 23548 15669 23576
rect 15657 23545 15669 23548
rect 15703 23545 15715 23579
rect 15657 23539 15715 23545
rect 16574 23536 16580 23588
rect 16632 23576 16638 23588
rect 17494 23576 17500 23588
rect 16632 23548 17500 23576
rect 16632 23536 16638 23548
rect 17494 23536 17500 23548
rect 17552 23536 17558 23588
rect 17586 23536 17592 23588
rect 17644 23576 17650 23588
rect 19168 23576 19196 23607
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20036 23616 20269 23644
rect 20036 23604 20042 23616
rect 20257 23613 20269 23616
rect 20303 23644 20315 23647
rect 20809 23647 20867 23653
rect 20809 23644 20821 23647
rect 20303 23616 20821 23644
rect 20303 23613 20315 23616
rect 20257 23607 20315 23613
rect 20809 23613 20821 23616
rect 20855 23613 20867 23647
rect 20809 23607 20867 23613
rect 20990 23604 20996 23656
rect 21048 23644 21054 23656
rect 21361 23647 21419 23653
rect 21361 23644 21373 23647
rect 21048 23616 21373 23644
rect 21048 23604 21054 23616
rect 21361 23613 21373 23616
rect 21407 23644 21419 23647
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21407 23616 21925 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 21913 23607 21971 23613
rect 22094 23604 22100 23656
rect 22152 23644 22158 23656
rect 22465 23647 22523 23653
rect 22465 23644 22477 23647
rect 22152 23616 22477 23644
rect 22152 23604 22158 23616
rect 22465 23613 22477 23616
rect 22511 23644 22523 23647
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22511 23616 23029 23644
rect 22511 23613 22523 23616
rect 22465 23607 22523 23613
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23017 23607 23075 23613
rect 19705 23579 19763 23585
rect 19705 23576 19717 23579
rect 17644 23548 19717 23576
rect 17644 23536 17650 23548
rect 19705 23545 19717 23548
rect 19751 23545 19763 23579
rect 19705 23539 19763 23545
rect 4706 23508 4712 23520
rect 4667 23480 4712 23508
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 9306 23468 9312 23520
rect 9364 23508 9370 23520
rect 9493 23511 9551 23517
rect 9493 23508 9505 23511
rect 9364 23480 9505 23508
rect 9364 23468 9370 23480
rect 9493 23477 9505 23480
rect 9539 23477 9551 23511
rect 9493 23471 9551 23477
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 11425 23511 11483 23517
rect 11425 23508 11437 23511
rect 10928 23480 11437 23508
rect 10928 23468 10934 23480
rect 11425 23477 11437 23480
rect 11471 23477 11483 23511
rect 14550 23508 14556 23520
rect 14511 23480 14556 23508
rect 11425 23471 11483 23477
rect 14550 23468 14556 23480
rect 14608 23468 14614 23520
rect 16022 23508 16028 23520
rect 15983 23480 16028 23508
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 16114 23468 16120 23520
rect 16172 23508 16178 23520
rect 17129 23511 17187 23517
rect 17129 23508 17141 23511
rect 16172 23480 17141 23508
rect 16172 23468 16178 23480
rect 17129 23477 17141 23480
rect 17175 23477 17187 23511
rect 17129 23471 17187 23477
rect 18322 23468 18328 23520
rect 18380 23508 18386 23520
rect 18782 23508 18788 23520
rect 18380 23480 18788 23508
rect 18380 23468 18386 23480
rect 18782 23468 18788 23480
rect 18840 23508 18846 23520
rect 18969 23511 19027 23517
rect 18969 23508 18981 23511
rect 18840 23480 18981 23508
rect 18840 23468 18846 23480
rect 18969 23477 18981 23480
rect 19015 23477 19027 23511
rect 21174 23508 21180 23520
rect 21135 23480 21180 23508
rect 18969 23471 19027 23477
rect 21174 23468 21180 23480
rect 21232 23468 21238 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 2406 23304 2412 23316
rect 2367 23276 2412 23304
rect 2406 23264 2412 23276
rect 2464 23264 2470 23316
rect 7006 23304 7012 23316
rect 6967 23276 7012 23304
rect 7006 23264 7012 23276
rect 7064 23264 7070 23316
rect 8294 23264 8300 23316
rect 8352 23304 8358 23316
rect 8481 23307 8539 23313
rect 8481 23304 8493 23307
rect 8352 23276 8493 23304
rect 8352 23264 8358 23276
rect 8481 23273 8493 23276
rect 8527 23273 8539 23307
rect 8481 23267 8539 23273
rect 10962 23264 10968 23316
rect 11020 23304 11026 23316
rect 11241 23307 11299 23313
rect 11241 23304 11253 23307
rect 11020 23276 11253 23304
rect 11020 23264 11026 23276
rect 11241 23273 11253 23276
rect 11287 23273 11299 23307
rect 11241 23267 11299 23273
rect 11422 23264 11428 23316
rect 11480 23304 11486 23316
rect 11609 23307 11667 23313
rect 11609 23304 11621 23307
rect 11480 23276 11621 23304
rect 11480 23264 11486 23276
rect 11609 23273 11621 23276
rect 11655 23304 11667 23307
rect 11882 23304 11888 23316
rect 11655 23276 11888 23304
rect 11655 23273 11667 23276
rect 11609 23267 11667 23273
rect 11882 23264 11888 23276
rect 11940 23264 11946 23316
rect 11977 23307 12035 23313
rect 11977 23273 11989 23307
rect 12023 23304 12035 23307
rect 12342 23304 12348 23316
rect 12023 23276 12348 23304
rect 12023 23273 12035 23276
rect 11977 23267 12035 23273
rect 12342 23264 12348 23276
rect 12400 23264 12406 23316
rect 13722 23264 13728 23316
rect 13780 23304 13786 23316
rect 14277 23307 14335 23313
rect 14277 23304 14289 23307
rect 13780 23276 14289 23304
rect 13780 23264 13786 23276
rect 14277 23273 14289 23276
rect 14323 23273 14335 23307
rect 16758 23304 16764 23316
rect 16719 23276 16764 23304
rect 14277 23267 14335 23273
rect 16758 23264 16764 23276
rect 16816 23264 16822 23316
rect 19518 23304 19524 23316
rect 19479 23276 19524 23304
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 1857 23239 1915 23245
rect 1857 23205 1869 23239
rect 1903 23236 1915 23239
rect 2038 23236 2044 23248
rect 1903 23208 2044 23236
rect 1903 23205 1915 23208
rect 1857 23199 1915 23205
rect 2038 23196 2044 23208
rect 2096 23196 2102 23248
rect 4332 23239 4390 23245
rect 4332 23205 4344 23239
rect 4378 23236 4390 23239
rect 4706 23236 4712 23248
rect 4378 23208 4712 23236
rect 4378 23205 4390 23208
rect 4332 23199 4390 23205
rect 4706 23196 4712 23208
rect 4764 23196 4770 23248
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 2682 23168 2688 23180
rect 1627 23140 2688 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2682 23128 2688 23140
rect 2740 23128 2746 23180
rect 2869 23171 2927 23177
rect 2869 23137 2881 23171
rect 2915 23137 2927 23171
rect 2869 23131 2927 23137
rect 3513 23171 3571 23177
rect 3513 23137 3525 23171
rect 3559 23168 3571 23171
rect 3881 23171 3939 23177
rect 3881 23168 3893 23171
rect 3559 23140 3893 23168
rect 3559 23137 3571 23140
rect 3513 23131 3571 23137
rect 3881 23137 3893 23140
rect 3927 23168 3939 23171
rect 4062 23168 4068 23180
rect 3927 23140 4068 23168
rect 3927 23137 3939 23140
rect 3881 23131 3939 23137
rect 2406 23060 2412 23112
rect 2464 23100 2470 23112
rect 2884 23100 2912 23131
rect 4062 23128 4068 23140
rect 4120 23128 4126 23180
rect 7024 23168 7052 23264
rect 10134 23245 10140 23248
rect 10128 23236 10140 23245
rect 10095 23208 10140 23236
rect 10128 23199 10140 23208
rect 10192 23236 10198 23248
rect 10870 23236 10876 23248
rect 10192 23208 10876 23236
rect 10134 23196 10140 23199
rect 10192 23196 10198 23208
rect 10870 23196 10876 23208
rect 10928 23196 10934 23248
rect 15562 23236 15568 23248
rect 15523 23208 15568 23236
rect 15562 23196 15568 23208
rect 15620 23196 15626 23248
rect 21177 23239 21235 23245
rect 21177 23205 21189 23239
rect 21223 23236 21235 23239
rect 22002 23236 22008 23248
rect 21223 23208 22008 23236
rect 21223 23205 21235 23208
rect 21177 23199 21235 23205
rect 22002 23196 22008 23208
rect 22060 23196 22066 23248
rect 7374 23177 7380 23180
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 7024 23140 7113 23168
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7368 23168 7380 23177
rect 7335 23140 7380 23168
rect 7101 23131 7159 23137
rect 7368 23131 7380 23140
rect 7374 23128 7380 23131
rect 7432 23128 7438 23180
rect 9125 23171 9183 23177
rect 9125 23137 9137 23171
rect 9171 23168 9183 23171
rect 9861 23171 9919 23177
rect 9861 23168 9873 23171
rect 9171 23140 9873 23168
rect 9171 23137 9183 23140
rect 9125 23131 9183 23137
rect 9861 23137 9873 23140
rect 9907 23168 9919 23171
rect 9950 23168 9956 23180
rect 9907 23140 9956 23168
rect 9907 23137 9919 23140
rect 9861 23131 9919 23137
rect 9950 23128 9956 23140
rect 10008 23128 10014 23180
rect 12342 23128 12348 23180
rect 12400 23168 12406 23180
rect 13153 23171 13211 23177
rect 13153 23168 13165 23171
rect 12400 23140 13165 23168
rect 12400 23128 12406 23140
rect 13153 23137 13165 23140
rect 13199 23137 13211 23171
rect 15286 23168 15292 23180
rect 15247 23140 15292 23168
rect 13153 23131 13211 23137
rect 15286 23128 15292 23140
rect 15344 23128 15350 23180
rect 16574 23168 16580 23180
rect 16535 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 19334 23168 19340 23180
rect 19295 23140 19340 23168
rect 19334 23128 19340 23140
rect 19392 23128 19398 23180
rect 20898 23168 20904 23180
rect 20859 23140 20904 23168
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 2464 23072 2912 23100
rect 12897 23103 12955 23109
rect 2464 23060 2470 23072
rect 12897 23069 12909 23103
rect 12943 23069 12955 23103
rect 12897 23063 12955 23069
rect 12912 22976 12940 23063
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 3053 22967 3111 22973
rect 3053 22964 3065 22967
rect 2924 22936 3065 22964
rect 2924 22924 2930 22936
rect 3053 22933 3065 22936
rect 3099 22933 3111 22967
rect 5442 22964 5448 22976
rect 5403 22936 5448 22964
rect 3053 22927 3111 22933
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 6457 22967 6515 22973
rect 6457 22933 6469 22967
rect 6503 22964 6515 22967
rect 6638 22964 6644 22976
rect 6503 22936 6644 22964
rect 6503 22933 6515 22936
rect 6457 22927 6515 22933
rect 6638 22924 6644 22936
rect 6696 22924 6702 22976
rect 9490 22964 9496 22976
rect 9451 22936 9496 22964
rect 9490 22924 9496 22936
rect 9548 22924 9554 22976
rect 12437 22967 12495 22973
rect 12437 22933 12449 22967
rect 12483 22964 12495 22967
rect 12805 22967 12863 22973
rect 12805 22964 12817 22967
rect 12483 22936 12817 22964
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 12805 22933 12817 22936
rect 12851 22964 12863 22967
rect 12894 22964 12900 22976
rect 12851 22936 12900 22964
rect 12851 22933 12863 22936
rect 12805 22927 12863 22933
rect 12894 22924 12900 22936
rect 12952 22924 12958 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 4706 22720 4712 22772
rect 4764 22760 4770 22772
rect 5813 22763 5871 22769
rect 5813 22760 5825 22763
rect 4764 22732 5825 22760
rect 4764 22720 4770 22732
rect 5813 22729 5825 22732
rect 5859 22729 5871 22763
rect 6362 22760 6368 22772
rect 6275 22732 6368 22760
rect 5813 22723 5871 22729
rect 6362 22720 6368 22732
rect 6420 22760 6426 22772
rect 7006 22760 7012 22772
rect 6420 22732 7012 22760
rect 6420 22720 6426 22732
rect 7006 22720 7012 22732
rect 7064 22720 7070 22772
rect 7282 22760 7288 22772
rect 7243 22732 7288 22760
rect 7282 22720 7288 22732
rect 7340 22720 7346 22772
rect 10134 22720 10140 22772
rect 10192 22760 10198 22772
rect 10413 22763 10471 22769
rect 10413 22760 10425 22763
rect 10192 22732 10425 22760
rect 10192 22720 10198 22732
rect 10413 22729 10425 22732
rect 10459 22729 10471 22763
rect 10413 22723 10471 22729
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12158 22760 12164 22772
rect 11931 22732 12164 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 2682 22652 2688 22704
rect 2740 22692 2746 22704
rect 3237 22695 3295 22701
rect 3237 22692 3249 22695
rect 2740 22664 3249 22692
rect 2740 22652 2746 22664
rect 3237 22661 3249 22664
rect 3283 22661 3295 22695
rect 4801 22695 4859 22701
rect 4801 22692 4813 22695
rect 3237 22655 3295 22661
rect 3712 22664 4813 22692
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3712 22633 3740 22664
rect 4801 22661 4813 22664
rect 4847 22661 4859 22695
rect 4801 22655 4859 22661
rect 3697 22627 3755 22633
rect 3697 22624 3709 22627
rect 3568 22596 3709 22624
rect 3568 22584 3574 22596
rect 3697 22593 3709 22596
rect 3743 22593 3755 22627
rect 3697 22587 3755 22593
rect 3789 22627 3847 22633
rect 3789 22593 3801 22627
rect 3835 22593 3847 22627
rect 3789 22587 3847 22593
rect 4709 22627 4767 22633
rect 4709 22593 4721 22627
rect 4755 22624 4767 22627
rect 5258 22624 5264 22636
rect 4755 22596 5264 22624
rect 4755 22593 4767 22596
rect 4709 22587 4767 22593
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22556 1547 22559
rect 2498 22556 2504 22568
rect 1535 22528 2504 22556
rect 1535 22525 1547 22528
rect 1489 22519 1547 22525
rect 2498 22516 2504 22528
rect 2556 22516 2562 22568
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 3804 22556 3832 22587
rect 5258 22584 5264 22596
rect 5316 22584 5322 22636
rect 5442 22624 5448 22636
rect 5403 22596 5448 22624
rect 5442 22584 5448 22596
rect 5500 22584 5506 22636
rect 6273 22627 6331 22633
rect 6273 22593 6285 22627
rect 6319 22624 6331 22627
rect 7374 22624 7380 22636
rect 6319 22596 7380 22624
rect 6319 22593 6331 22596
rect 6273 22587 6331 22593
rect 7374 22584 7380 22596
rect 7432 22624 7438 22636
rect 7837 22627 7895 22633
rect 7837 22624 7849 22627
rect 7432 22596 7849 22624
rect 7432 22584 7438 22596
rect 7837 22593 7849 22596
rect 7883 22624 7895 22627
rect 8110 22624 8116 22636
rect 7883 22596 8116 22624
rect 7883 22593 7895 22596
rect 7837 22587 7895 22593
rect 8110 22584 8116 22596
rect 8168 22624 8174 22636
rect 8665 22627 8723 22633
rect 8665 22624 8677 22627
rect 8168 22596 8677 22624
rect 8168 22584 8174 22596
rect 8665 22593 8677 22596
rect 8711 22593 8723 22627
rect 8665 22587 8723 22593
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 9950 22624 9956 22636
rect 9548 22596 9956 22624
rect 9548 22584 9554 22596
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 4246 22556 4252 22568
rect 2823 22528 4252 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 4246 22516 4252 22528
rect 4304 22516 4310 22568
rect 4341 22559 4399 22565
rect 4341 22525 4353 22559
rect 4387 22556 4399 22559
rect 5166 22556 5172 22568
rect 4387 22528 5172 22556
rect 4387 22525 4399 22528
rect 4341 22519 4399 22525
rect 5166 22516 5172 22528
rect 5224 22516 5230 22568
rect 6549 22559 6607 22565
rect 6549 22525 6561 22559
rect 6595 22556 6607 22559
rect 6638 22556 6644 22568
rect 6595 22528 6644 22556
rect 6595 22525 6607 22528
rect 6549 22519 6607 22525
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7193 22559 7251 22565
rect 7193 22525 7205 22559
rect 7239 22556 7251 22559
rect 7742 22556 7748 22568
rect 7239 22528 7748 22556
rect 7239 22525 7251 22528
rect 7193 22519 7251 22525
rect 7742 22516 7748 22528
rect 7800 22516 7806 22568
rect 9858 22556 9864 22568
rect 9819 22528 9864 22556
rect 9858 22516 9864 22528
rect 9916 22556 9922 22568
rect 10781 22559 10839 22565
rect 10781 22556 10793 22559
rect 9916 22528 10793 22556
rect 9916 22516 9922 22528
rect 10781 22525 10793 22528
rect 10827 22525 10839 22559
rect 10781 22519 10839 22525
rect 11057 22559 11115 22565
rect 11057 22525 11069 22559
rect 11103 22556 11115 22559
rect 11900 22556 11928 22723
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 14461 22763 14519 22769
rect 14461 22760 14473 22763
rect 13096 22732 14473 22760
rect 12253 22695 12311 22701
rect 12253 22661 12265 22695
rect 12299 22692 12311 22695
rect 12342 22692 12348 22704
rect 12299 22664 12348 22692
rect 12299 22661 12311 22664
rect 12253 22655 12311 22661
rect 12342 22652 12348 22664
rect 12400 22692 12406 22704
rect 13096 22692 13124 22732
rect 14461 22729 14473 22732
rect 14507 22760 14519 22763
rect 14550 22760 14556 22772
rect 14507 22732 14556 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 14550 22720 14556 22732
rect 14608 22720 14614 22772
rect 15286 22720 15292 22772
rect 15344 22760 15350 22772
rect 15746 22760 15752 22772
rect 15344 22732 15752 22760
rect 15344 22720 15350 22732
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 12400 22664 13124 22692
rect 12400 22652 12406 22664
rect 12986 22584 12992 22636
rect 13044 22624 13050 22636
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 13044 22596 13093 22624
rect 13044 22584 13050 22596
rect 13081 22593 13093 22596
rect 13127 22593 13139 22627
rect 13081 22587 13139 22593
rect 15289 22627 15347 22633
rect 15289 22593 15301 22627
rect 15335 22624 15347 22627
rect 15378 22624 15384 22636
rect 15335 22596 15384 22624
rect 15335 22593 15347 22596
rect 15289 22587 15347 22593
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 11103 22528 11928 22556
rect 11103 22525 11115 22528
rect 11057 22519 11115 22525
rect 3145 22491 3203 22497
rect 3145 22457 3157 22491
rect 3191 22488 3203 22491
rect 3605 22491 3663 22497
rect 3605 22488 3617 22491
rect 3191 22460 3617 22488
rect 3191 22457 3203 22460
rect 3145 22451 3203 22457
rect 3605 22457 3617 22460
rect 3651 22488 3663 22491
rect 3694 22488 3700 22500
rect 3651 22460 3700 22488
rect 3651 22457 3663 22460
rect 3605 22451 3663 22457
rect 3694 22448 3700 22460
rect 3752 22448 3758 22500
rect 7653 22491 7711 22497
rect 7653 22457 7665 22491
rect 7699 22488 7711 22491
rect 8294 22488 8300 22500
rect 7699 22460 8300 22488
rect 7699 22457 7711 22460
rect 7653 22451 7711 22457
rect 8294 22448 8300 22460
rect 8352 22448 8358 22500
rect 9309 22491 9367 22497
rect 9309 22457 9321 22491
rect 9355 22488 9367 22491
rect 11330 22488 11336 22500
rect 9355 22460 9812 22488
rect 11291 22460 11336 22488
rect 9355 22457 9367 22460
rect 9309 22451 9367 22457
rect 9784 22432 9812 22460
rect 11330 22448 11336 22460
rect 11388 22448 11394 22500
rect 12989 22491 13047 22497
rect 12989 22457 13001 22491
rect 13035 22488 13047 22491
rect 13326 22491 13384 22497
rect 13326 22488 13338 22491
rect 13035 22460 13338 22488
rect 13035 22457 13047 22460
rect 12989 22451 13047 22457
rect 13096 22432 13124 22460
rect 13326 22457 13338 22460
rect 13372 22457 13384 22491
rect 13326 22451 13384 22457
rect 2406 22420 2412 22432
rect 2367 22392 2412 22420
rect 2406 22380 2412 22392
rect 2464 22380 2470 22432
rect 9398 22420 9404 22432
rect 9359 22392 9404 22420
rect 9398 22380 9404 22392
rect 9456 22380 9462 22432
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 13078 22380 13084 22432
rect 13136 22380 13142 22432
rect 14734 22420 14740 22432
rect 14695 22392 14740 22420
rect 14734 22380 14740 22392
rect 14792 22380 14798 22432
rect 16574 22420 16580 22432
rect 16535 22392 16580 22420
rect 16574 22380 16580 22392
rect 16632 22380 16638 22432
rect 19334 22420 19340 22432
rect 19295 22392 19340 22420
rect 19334 22380 19340 22392
rect 19392 22380 19398 22432
rect 20898 22420 20904 22432
rect 20859 22392 20904 22420
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2409 22219 2467 22225
rect 2409 22185 2421 22219
rect 2455 22216 2467 22219
rect 2498 22216 2504 22228
rect 2455 22188 2504 22216
rect 2455 22185 2467 22188
rect 2409 22179 2467 22185
rect 2498 22176 2504 22188
rect 2556 22176 2562 22228
rect 2682 22216 2688 22228
rect 2643 22188 2688 22216
rect 2682 22176 2688 22188
rect 2740 22176 2746 22228
rect 3510 22216 3516 22228
rect 3471 22188 3516 22216
rect 3510 22176 3516 22188
rect 3568 22176 3574 22228
rect 5813 22219 5871 22225
rect 5813 22185 5825 22219
rect 5859 22216 5871 22219
rect 6181 22219 6239 22225
rect 6181 22216 6193 22219
rect 5859 22188 6193 22216
rect 5859 22185 5871 22188
rect 5813 22179 5871 22185
rect 6181 22185 6193 22188
rect 6227 22216 6239 22219
rect 6362 22216 6368 22228
rect 6227 22188 6368 22216
rect 6227 22185 6239 22188
rect 6181 22179 6239 22185
rect 6362 22176 6368 22188
rect 6420 22176 6426 22228
rect 16298 22216 16304 22228
rect 16259 22188 16304 22216
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 3881 22151 3939 22157
rect 3881 22148 3893 22151
rect 3791 22120 3893 22148
rect 3881 22117 3893 22120
rect 3927 22148 3939 22151
rect 4062 22148 4068 22160
rect 3927 22120 4068 22148
rect 3927 22117 3939 22120
rect 3881 22111 3939 22117
rect 1578 22080 1584 22092
rect 1539 22052 1584 22080
rect 1578 22040 1584 22052
rect 1636 22040 1642 22092
rect 1854 22080 1860 22092
rect 1815 22052 1860 22080
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 2869 22083 2927 22089
rect 2869 22049 2881 22083
rect 2915 22080 2927 22083
rect 3694 22080 3700 22092
rect 2915 22052 3700 22080
rect 2915 22049 2927 22052
rect 2869 22043 2927 22049
rect 3694 22040 3700 22052
rect 3752 22040 3758 22092
rect 3896 22012 3924 22111
rect 4062 22108 4068 22120
rect 4120 22108 4126 22160
rect 10042 22148 10048 22160
rect 9968 22120 10048 22148
rect 4338 22089 4344 22092
rect 4332 22080 4344 22089
rect 4299 22052 4344 22080
rect 4332 22043 4344 22052
rect 4338 22040 4344 22043
rect 4396 22040 4402 22092
rect 6454 22040 6460 22092
rect 6512 22080 6518 22092
rect 6825 22083 6883 22089
rect 6825 22080 6837 22083
rect 6512 22052 6837 22080
rect 6512 22040 6518 22052
rect 6825 22049 6837 22052
rect 6871 22049 6883 22083
rect 6825 22043 6883 22049
rect 8297 22083 8355 22089
rect 8297 22049 8309 22083
rect 8343 22080 8355 22083
rect 8386 22080 8392 22092
rect 8343 22052 8392 22080
rect 8343 22049 8355 22052
rect 8297 22043 8355 22049
rect 8386 22040 8392 22052
rect 8444 22080 8450 22092
rect 9582 22080 9588 22092
rect 8444 22052 9588 22080
rect 8444 22040 8450 22052
rect 9582 22040 9588 22052
rect 9640 22040 9646 22092
rect 9968 22089 9996 22120
rect 10042 22108 10048 22120
rect 10100 22108 10106 22160
rect 15286 22148 15292 22160
rect 15247 22120 15292 22148
rect 15286 22108 15292 22120
rect 15344 22108 15350 22160
rect 9953 22083 10011 22089
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10220 22083 10278 22089
rect 9999 22052 10033 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10220 22049 10232 22083
rect 10266 22080 10278 22083
rect 10502 22080 10508 22092
rect 10266 22052 10508 22080
rect 10266 22049 10278 22052
rect 10220 22043 10278 22049
rect 10502 22040 10508 22052
rect 10560 22080 10566 22092
rect 10962 22080 10968 22092
rect 10560 22052 10968 22080
rect 10560 22040 10566 22052
rect 10962 22040 10968 22052
rect 11020 22040 11026 22092
rect 11238 22040 11244 22092
rect 11296 22080 11302 22092
rect 12069 22083 12127 22089
rect 12069 22080 12081 22083
rect 11296 22052 12081 22080
rect 11296 22040 11302 22052
rect 12069 22049 12081 22052
rect 12115 22080 12127 22083
rect 12345 22083 12403 22089
rect 12345 22080 12357 22083
rect 12115 22052 12357 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 12345 22049 12357 22052
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12897 22083 12955 22089
rect 12897 22049 12909 22083
rect 12943 22080 12955 22083
rect 13245 22083 13303 22089
rect 13245 22080 13257 22083
rect 12943 22052 13257 22080
rect 12943 22049 12955 22052
rect 12897 22043 12955 22049
rect 13245 22049 13257 22052
rect 13291 22080 13303 22083
rect 14642 22080 14648 22092
rect 13291 22052 14648 22080
rect 13291 22049 13303 22052
rect 13245 22043 13303 22049
rect 14642 22040 14648 22052
rect 14700 22040 14706 22092
rect 4062 22012 4068 22024
rect 3896 21984 4068 22012
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 6914 22012 6920 22024
rect 6875 21984 6920 22012
rect 6914 21972 6920 21984
rect 6972 21972 6978 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 8478 22012 8484 22024
rect 7064 21984 7109 22012
rect 8439 21984 8484 22012
rect 7064 21972 7070 21984
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 12986 22012 12992 22024
rect 12176 21984 12992 22012
rect 3050 21944 3056 21956
rect 3011 21916 3056 21944
rect 3050 21904 3056 21916
rect 3108 21904 3114 21956
rect 12176 21953 12204 21984
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 12161 21947 12219 21953
rect 12161 21913 12173 21947
rect 12207 21913 12219 21947
rect 12161 21907 12219 21913
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 4430 21876 4436 21888
rect 4304 21848 4436 21876
rect 4304 21836 4310 21848
rect 4430 21836 4436 21848
rect 4488 21876 4494 21888
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 4488 21848 5457 21876
rect 4488 21836 4494 21848
rect 5445 21845 5457 21848
rect 5491 21845 5503 21879
rect 5445 21839 5503 21845
rect 5534 21836 5540 21888
rect 5592 21876 5598 21888
rect 6457 21879 6515 21885
rect 6457 21876 6469 21879
rect 5592 21848 6469 21876
rect 5592 21836 5598 21848
rect 6457 21845 6469 21848
rect 6503 21845 6515 21879
rect 7650 21876 7656 21888
rect 7611 21848 7656 21876
rect 6457 21839 6515 21845
rect 7650 21836 7656 21848
rect 7708 21836 7714 21888
rect 8021 21879 8079 21885
rect 8021 21845 8033 21879
rect 8067 21876 8079 21879
rect 8202 21876 8208 21888
rect 8067 21848 8208 21876
rect 8067 21845 8079 21848
rect 8021 21839 8079 21845
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 9398 21876 9404 21888
rect 9359 21848 9404 21876
rect 9398 21836 9404 21848
rect 9456 21836 9462 21888
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 11333 21879 11391 21885
rect 11333 21876 11345 21879
rect 10008 21848 11345 21876
rect 10008 21836 10014 21848
rect 11333 21845 11345 21848
rect 11379 21845 11391 21879
rect 11333 21839 11391 21845
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 14369 21879 14427 21885
rect 14369 21876 14381 21879
rect 13228 21848 14381 21876
rect 13228 21836 13234 21848
rect 14369 21845 14381 21848
rect 14415 21845 14427 21879
rect 14369 21839 14427 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2406 21672 2412 21684
rect 2367 21644 2412 21672
rect 2406 21632 2412 21644
rect 2464 21632 2470 21684
rect 3694 21672 3700 21684
rect 3655 21644 3700 21672
rect 3694 21632 3700 21644
rect 3752 21632 3758 21684
rect 4065 21675 4123 21681
rect 4065 21641 4077 21675
rect 4111 21672 4123 21675
rect 4338 21672 4344 21684
rect 4111 21644 4344 21672
rect 4111 21641 4123 21644
rect 4065 21635 4123 21641
rect 4338 21632 4344 21644
rect 4396 21672 4402 21684
rect 4893 21675 4951 21681
rect 4893 21672 4905 21675
rect 4396 21644 4905 21672
rect 4396 21632 4402 21644
rect 4893 21641 4905 21644
rect 4939 21672 4951 21675
rect 5442 21672 5448 21684
rect 4939 21644 5448 21672
rect 4939 21641 4951 21644
rect 4893 21635 4951 21641
rect 5442 21632 5448 21644
rect 5500 21632 5506 21684
rect 5905 21675 5963 21681
rect 5905 21641 5917 21675
rect 5951 21672 5963 21675
rect 5994 21672 6000 21684
rect 5951 21644 6000 21672
rect 5951 21641 5963 21644
rect 5905 21635 5963 21641
rect 1578 21564 1584 21616
rect 1636 21604 1642 21616
rect 2682 21604 2688 21616
rect 1636 21576 2688 21604
rect 1636 21564 1642 21576
rect 2682 21564 2688 21576
rect 2740 21564 2746 21616
rect 2774 21564 2780 21616
rect 2832 21604 2838 21616
rect 2832 21576 3096 21604
rect 2832 21564 2838 21576
rect 3068 21545 3096 21576
rect 4154 21564 4160 21616
rect 4212 21604 4218 21616
rect 5920 21604 5948 21635
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 10413 21675 10471 21681
rect 10413 21641 10425 21675
rect 10459 21672 10471 21675
rect 10502 21672 10508 21684
rect 10459 21644 10508 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 13446 21632 13452 21684
rect 13504 21672 13510 21684
rect 13541 21675 13599 21681
rect 13541 21672 13553 21675
rect 13504 21644 13553 21672
rect 13504 21632 13510 21644
rect 13541 21641 13553 21644
rect 13587 21641 13599 21675
rect 13541 21635 13599 21641
rect 13814 21632 13820 21684
rect 13872 21672 13878 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 13872 21644 13921 21672
rect 13872 21632 13878 21644
rect 13909 21641 13921 21644
rect 13955 21672 13967 21675
rect 13955 21644 14596 21672
rect 13955 21641 13967 21644
rect 13909 21635 13967 21641
rect 4212 21576 5948 21604
rect 10965 21607 11023 21613
rect 4212 21564 4218 21576
rect 10965 21573 10977 21607
rect 11011 21604 11023 21607
rect 12529 21607 12587 21613
rect 12529 21604 12541 21607
rect 11011 21576 12541 21604
rect 11011 21573 11023 21576
rect 10965 21567 11023 21573
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 3053 21499 3111 21505
rect 3881 21539 3939 21545
rect 3881 21505 3893 21539
rect 3927 21536 3939 21539
rect 7469 21539 7527 21545
rect 3927 21508 5304 21536
rect 3927 21505 3939 21508
rect 3881 21499 3939 21505
rect 1581 21471 1639 21477
rect 1581 21437 1593 21471
rect 1627 21468 1639 21471
rect 2406 21468 2412 21480
rect 1627 21440 2412 21468
rect 1627 21437 1639 21440
rect 1581 21431 1639 21437
rect 2406 21428 2412 21440
rect 2464 21428 2470 21480
rect 2869 21471 2927 21477
rect 2869 21437 2881 21471
rect 2915 21468 2927 21471
rect 3510 21468 3516 21480
rect 2915 21440 3516 21468
rect 2915 21437 2927 21440
rect 2869 21431 2927 21437
rect 3510 21428 3516 21440
rect 3568 21428 3574 21480
rect 4154 21477 4160 21480
rect 4145 21471 4160 21477
rect 4145 21437 4157 21471
rect 4145 21431 4160 21437
rect 4154 21428 4160 21431
rect 4212 21428 4218 21480
rect 5276 21477 5304 21508
rect 7469 21505 7481 21539
rect 7515 21536 7527 21539
rect 8018 21536 8024 21548
rect 7515 21508 8024 21536
rect 7515 21505 7527 21508
rect 7469 21499 7527 21505
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 8202 21536 8208 21548
rect 8163 21508 8208 21536
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 8849 21539 8907 21545
rect 8849 21505 8861 21539
rect 8895 21536 8907 21539
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 8895 21508 9873 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 9861 21505 9873 21508
rect 9907 21536 9919 21539
rect 10778 21536 10784 21548
rect 9907 21508 10784 21536
rect 9907 21505 9919 21508
rect 9861 21499 9919 21505
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21468 5319 21471
rect 5718 21468 5724 21480
rect 5307 21440 5724 21468
rect 5307 21437 5319 21440
rect 5261 21431 5319 21437
rect 5718 21428 5724 21440
rect 5776 21428 5782 21480
rect 7650 21428 7656 21480
rect 7708 21468 7714 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7708 21440 7941 21468
rect 7708 21428 7714 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 7929 21431 7987 21437
rect 9217 21471 9275 21477
rect 9217 21437 9229 21471
rect 9263 21468 9275 21471
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9263 21440 9781 21468
rect 9263 21437 9275 21440
rect 9217 21431 9275 21437
rect 9769 21437 9781 21440
rect 9815 21468 9827 21471
rect 10962 21468 10968 21480
rect 9815 21440 10968 21468
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 10962 21428 10968 21440
rect 11020 21428 11026 21480
rect 11072 21477 11100 21576
rect 12529 21573 12541 21576
rect 12575 21573 12587 21607
rect 14093 21607 14151 21613
rect 14093 21604 14105 21607
rect 12529 21567 12587 21573
rect 13004 21576 14105 21604
rect 13004 21545 13032 21576
rect 14093 21573 14105 21576
rect 14139 21573 14151 21607
rect 14093 21567 14151 21573
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21437 11115 21471
rect 11057 21431 11115 21437
rect 12253 21471 12311 21477
rect 12253 21437 12265 21471
rect 12299 21468 12311 21471
rect 12894 21468 12900 21480
rect 12299 21440 12900 21468
rect 12299 21437 12311 21440
rect 12253 21431 12311 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 1857 21403 1915 21409
rect 1857 21369 1869 21403
rect 1903 21369 1915 21403
rect 1857 21363 1915 21369
rect 11333 21403 11391 21409
rect 11333 21369 11345 21403
rect 11379 21369 11391 21403
rect 11333 21363 11391 21369
rect 11885 21403 11943 21409
rect 11885 21369 11897 21403
rect 11931 21400 11943 21403
rect 13004 21400 13032 21499
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 14568 21545 14596 21644
rect 14553 21539 14611 21545
rect 13136 21508 13181 21536
rect 13136 21496 13142 21508
rect 14553 21505 14565 21539
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 14642 21496 14648 21548
rect 14700 21536 14706 21548
rect 15105 21539 15163 21545
rect 15105 21536 15117 21539
rect 14700 21508 15117 21536
rect 14700 21496 14706 21508
rect 15105 21505 15117 21508
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 15657 21539 15715 21545
rect 15657 21536 15669 21539
rect 15436 21508 15669 21536
rect 15436 21496 15442 21508
rect 15657 21505 15669 21508
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 13446 21428 13452 21480
rect 13504 21468 13510 21480
rect 14461 21471 14519 21477
rect 14461 21468 14473 21471
rect 13504 21440 14473 21468
rect 13504 21428 13510 21440
rect 14461 21437 14473 21440
rect 14507 21437 14519 21471
rect 14461 21431 14519 21437
rect 11931 21372 13032 21400
rect 11931 21369 11943 21372
rect 11885 21363 11943 21369
rect 1872 21332 1900 21363
rect 3881 21335 3939 21341
rect 3881 21332 3893 21335
rect 1872 21304 3893 21332
rect 3881 21301 3893 21304
rect 3927 21301 3939 21335
rect 3881 21295 3939 21301
rect 3970 21292 3976 21344
rect 4028 21332 4034 21344
rect 4341 21335 4399 21341
rect 4341 21332 4353 21335
rect 4028 21304 4353 21332
rect 4028 21292 4034 21304
rect 4341 21301 4353 21304
rect 4387 21301 4399 21335
rect 5442 21332 5448 21344
rect 5403 21304 5448 21332
rect 4341 21295 4399 21301
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 6454 21332 6460 21344
rect 6415 21304 6460 21332
rect 6454 21292 6460 21304
rect 6512 21292 6518 21344
rect 7006 21332 7012 21344
rect 6967 21304 7012 21332
rect 7006 21292 7012 21304
rect 7064 21292 7070 21344
rect 7558 21332 7564 21344
rect 7519 21304 7564 21332
rect 7558 21292 7564 21304
rect 7616 21292 7622 21344
rect 8846 21292 8852 21344
rect 8904 21332 8910 21344
rect 9309 21335 9367 21341
rect 9309 21332 9321 21335
rect 8904 21304 9321 21332
rect 8904 21292 8910 21304
rect 9309 21301 9321 21304
rect 9355 21301 9367 21335
rect 9309 21295 9367 21301
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 9677 21335 9735 21341
rect 9677 21332 9689 21335
rect 9456 21304 9689 21332
rect 9456 21292 9462 21304
rect 9677 21301 9689 21304
rect 9723 21332 9735 21335
rect 10042 21332 10048 21344
rect 9723 21304 10048 21332
rect 9723 21301 9735 21304
rect 9677 21295 9735 21301
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11348 21332 11376 21363
rect 11112 21304 11376 21332
rect 11112 21292 11118 21304
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 2958 21128 2964 21140
rect 2919 21100 2964 21128
rect 2958 21088 2964 21100
rect 3016 21088 3022 21140
rect 3510 21128 3516 21140
rect 3471 21100 3516 21128
rect 3510 21088 3516 21100
rect 3568 21088 3574 21140
rect 5718 21128 5724 21140
rect 5679 21100 5724 21128
rect 5718 21088 5724 21100
rect 5776 21088 5782 21140
rect 6549 21131 6607 21137
rect 6549 21097 6561 21131
rect 6595 21128 6607 21131
rect 6914 21128 6920 21140
rect 6595 21100 6920 21128
rect 6595 21097 6607 21100
rect 6549 21091 6607 21097
rect 6914 21088 6920 21100
rect 6972 21128 6978 21140
rect 7558 21128 7564 21140
rect 6972 21100 7564 21128
rect 6972 21088 6978 21100
rect 7558 21088 7564 21100
rect 7616 21088 7622 21140
rect 8110 21128 8116 21140
rect 8071 21100 8116 21128
rect 8110 21088 8116 21100
rect 8168 21088 8174 21140
rect 8386 21128 8392 21140
rect 8347 21100 8392 21128
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 9306 21128 9312 21140
rect 9267 21100 9312 21128
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 10778 21088 10784 21140
rect 10836 21128 10842 21140
rect 11057 21131 11115 21137
rect 11057 21128 11069 21131
rect 10836 21100 11069 21128
rect 10836 21088 10842 21100
rect 11057 21097 11069 21100
rect 11103 21097 11115 21131
rect 12066 21128 12072 21140
rect 12027 21100 12072 21128
rect 11057 21091 11115 21097
rect 12066 21088 12072 21100
rect 12124 21088 12130 21140
rect 12621 21131 12679 21137
rect 12621 21097 12633 21131
rect 12667 21128 12679 21131
rect 13078 21128 13084 21140
rect 12667 21100 13084 21128
rect 12667 21097 12679 21100
rect 12621 21091 12679 21097
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 14369 21131 14427 21137
rect 14369 21097 14381 21131
rect 14415 21128 14427 21131
rect 14642 21128 14648 21140
rect 14415 21100 14648 21128
rect 14415 21097 14427 21100
rect 14369 21091 14427 21097
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 4332 21063 4390 21069
rect 4332 21029 4344 21063
rect 4378 21060 4390 21063
rect 4430 21060 4436 21072
rect 4378 21032 4436 21060
rect 4378 21029 4390 21032
rect 4332 21023 4390 21029
rect 4430 21020 4436 21032
rect 4488 21020 4494 21072
rect 8757 21063 8815 21069
rect 8757 21060 8769 21063
rect 6840 21032 8769 21060
rect 6840 21004 6868 21032
rect 8757 21029 8769 21032
rect 8803 21060 8815 21063
rect 9125 21063 9183 21069
rect 9125 21060 9137 21063
rect 8803 21032 9137 21060
rect 8803 21029 8815 21032
rect 8757 21023 8815 21029
rect 9125 21029 9137 21032
rect 9171 21029 9183 21063
rect 9125 21023 9183 21029
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 9950 21069 9956 21072
rect 9922 21063 9956 21069
rect 9922 21060 9934 21063
rect 9732 21032 9934 21060
rect 9732 21020 9738 21032
rect 9922 21029 9934 21032
rect 10008 21060 10014 21072
rect 10008 21032 10070 21060
rect 9922 21023 9956 21029
rect 9950 21020 9956 21023
rect 10008 21020 10014 21032
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20961 1731 20995
rect 1946 20992 1952 21004
rect 1907 20964 1952 20992
rect 1673 20955 1731 20961
rect 1688 20924 1716 20955
rect 1946 20952 1952 20964
rect 2004 20952 2010 21004
rect 4062 20992 4068 21004
rect 4023 20964 4068 20992
rect 4062 20952 4068 20964
rect 4120 20952 4126 21004
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 6733 20995 6791 21001
rect 6733 20992 6745 20995
rect 6420 20964 6745 20992
rect 6420 20952 6426 20964
rect 6733 20961 6745 20964
rect 6779 20992 6791 20995
rect 6822 20992 6828 21004
rect 6779 20964 6828 20992
rect 6779 20961 6791 20964
rect 6733 20955 6791 20961
rect 6822 20952 6828 20964
rect 6880 20952 6886 21004
rect 7006 21001 7012 21004
rect 7000 20992 7012 21001
rect 6967 20964 7012 20992
rect 7000 20955 7012 20964
rect 7006 20952 7012 20955
rect 7064 20952 7070 21004
rect 8570 20952 8576 21004
rect 8628 20992 8634 21004
rect 9493 20995 9551 21001
rect 9493 20992 9505 20995
rect 8628 20964 9505 20992
rect 8628 20952 8634 20964
rect 9493 20961 9505 20964
rect 9539 20961 9551 20995
rect 11882 20992 11888 21004
rect 11843 20964 11888 20992
rect 9493 20955 9551 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 13078 20952 13084 21004
rect 13136 20992 13142 21004
rect 13245 20995 13303 21001
rect 13245 20992 13257 20995
rect 13136 20964 13257 20992
rect 13136 20952 13142 20964
rect 13245 20961 13257 20964
rect 13291 20961 13303 20995
rect 13245 20955 13303 20961
rect 9677 20927 9735 20933
rect 1688 20896 1992 20924
rect 1964 20868 1992 20896
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 12986 20924 12992 20936
rect 12899 20896 12992 20924
rect 9677 20887 9735 20893
rect 1946 20816 1952 20868
rect 2004 20816 2010 20868
rect 2314 20748 2320 20800
rect 2372 20788 2378 20800
rect 2409 20791 2467 20797
rect 2409 20788 2421 20791
rect 2372 20760 2421 20788
rect 2372 20748 2378 20760
rect 2409 20757 2421 20760
rect 2455 20757 2467 20791
rect 2409 20751 2467 20757
rect 2774 20748 2780 20800
rect 2832 20788 2838 20800
rect 3878 20788 3884 20800
rect 2832 20760 2877 20788
rect 3839 20760 3884 20788
rect 2832 20748 2838 20760
rect 3878 20748 3884 20760
rect 3936 20748 3942 20800
rect 5442 20788 5448 20800
rect 5403 20760 5448 20788
rect 5442 20748 5448 20760
rect 5500 20748 5506 20800
rect 6086 20788 6092 20800
rect 6047 20760 6092 20788
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 9582 20748 9588 20800
rect 9640 20788 9646 20800
rect 9692 20788 9720 20887
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 10612 20828 11192 20856
rect 10612 20788 10640 20828
rect 11164 20800 11192 20828
rect 9640 20760 10640 20788
rect 9640 20748 9646 20760
rect 11146 20748 11152 20800
rect 11204 20788 11210 20800
rect 11425 20791 11483 20797
rect 11425 20788 11437 20791
rect 11204 20760 11437 20788
rect 11204 20748 11210 20760
rect 11425 20757 11437 20760
rect 11471 20788 11483 20791
rect 13004 20788 13032 20884
rect 14734 20788 14740 20800
rect 11471 20760 14740 20788
rect 11471 20757 11483 20760
rect 11425 20751 11483 20757
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 4430 20584 4436 20596
rect 4391 20556 4436 20584
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 7006 20584 7012 20596
rect 6687 20556 7012 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 7006 20544 7012 20556
rect 7064 20584 7070 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 7064 20556 8217 20584
rect 7064 20544 7070 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 8570 20584 8576 20596
rect 8531 20556 8576 20584
rect 8205 20547 8263 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 8941 20587 8999 20593
rect 8941 20553 8953 20587
rect 8987 20584 8999 20587
rect 9674 20584 9680 20596
rect 8987 20556 9680 20584
rect 8987 20553 8999 20556
rect 8941 20547 8999 20553
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 10410 20584 10416 20596
rect 10371 20556 10416 20584
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11146 20584 11152 20596
rect 11107 20556 11152 20584
rect 11146 20544 11152 20556
rect 11204 20544 11210 20596
rect 11882 20584 11888 20596
rect 11843 20556 11888 20584
rect 11882 20544 11888 20556
rect 11940 20544 11946 20596
rect 12989 20587 13047 20593
rect 12989 20553 13001 20587
rect 13035 20584 13047 20587
rect 13078 20584 13084 20596
rect 13035 20556 13084 20584
rect 13035 20553 13047 20556
rect 12989 20547 13047 20553
rect 13078 20544 13084 20556
rect 13136 20584 13142 20596
rect 14461 20587 14519 20593
rect 14461 20584 14473 20587
rect 13136 20556 14473 20584
rect 13136 20544 13142 20556
rect 14461 20553 14473 20556
rect 14507 20584 14519 20587
rect 14550 20584 14556 20596
rect 14507 20556 14556 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 14734 20584 14740 20596
rect 14695 20556 14740 20584
rect 14734 20544 14740 20556
rect 14792 20544 14798 20596
rect 2406 20516 2412 20528
rect 2367 20488 2412 20516
rect 2406 20476 2412 20488
rect 2464 20476 2470 20528
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20448 1455 20451
rect 2130 20448 2136 20460
rect 1443 20420 2136 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2222 20408 2228 20460
rect 2280 20448 2286 20460
rect 2869 20451 2927 20457
rect 2869 20448 2881 20451
rect 2280 20420 2881 20448
rect 2280 20408 2286 20420
rect 2869 20417 2881 20420
rect 2915 20417 2927 20451
rect 3050 20448 3056 20460
rect 3011 20420 3056 20448
rect 2869 20411 2927 20417
rect 3050 20408 3056 20420
rect 3108 20408 3114 20460
rect 5442 20408 5448 20460
rect 5500 20448 5506 20460
rect 5537 20451 5595 20457
rect 5537 20448 5549 20451
rect 5500 20420 5549 20448
rect 5500 20408 5506 20420
rect 5537 20417 5549 20420
rect 5583 20448 5595 20451
rect 5997 20451 6055 20457
rect 5997 20448 6009 20451
rect 5583 20420 6009 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 5997 20417 6009 20420
rect 6043 20417 6055 20451
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 5997 20411 6055 20417
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 2317 20383 2375 20389
rect 2317 20349 2329 20383
rect 2363 20380 2375 20383
rect 3068 20380 3096 20408
rect 2363 20352 3096 20380
rect 4893 20383 4951 20389
rect 2363 20349 2375 20352
rect 2317 20343 2375 20349
rect 4893 20349 4905 20383
rect 4939 20380 4951 20383
rect 5350 20380 5356 20392
rect 4939 20352 5356 20380
rect 4939 20349 4951 20352
rect 4893 20343 4951 20349
rect 5350 20340 5356 20352
rect 5408 20380 5414 20392
rect 5408 20352 5488 20380
rect 5408 20340 5414 20352
rect 2774 20272 2780 20324
rect 2832 20312 2838 20324
rect 5460 20321 5488 20352
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7092 20383 7150 20389
rect 7092 20380 7104 20383
rect 6972 20352 7104 20380
rect 6972 20340 6978 20352
rect 7092 20349 7104 20352
rect 7138 20380 7150 20383
rect 8202 20380 8208 20392
rect 7138 20352 8208 20380
rect 7138 20349 7150 20352
rect 7092 20343 7150 20349
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 9033 20383 9091 20389
rect 9033 20349 9045 20383
rect 9079 20380 9091 20383
rect 9582 20380 9588 20392
rect 9079 20352 9588 20380
rect 9079 20349 9091 20352
rect 9033 20343 9091 20349
rect 9582 20340 9588 20352
rect 9640 20340 9646 20392
rect 13078 20380 13084 20392
rect 13039 20352 13084 20380
rect 13078 20340 13084 20352
rect 13136 20340 13142 20392
rect 9306 20321 9312 20324
rect 5445 20315 5503 20321
rect 2832 20284 2877 20312
rect 2832 20272 2838 20284
rect 5445 20281 5457 20315
rect 5491 20281 5503 20315
rect 9300 20312 9312 20321
rect 9267 20284 9312 20312
rect 5445 20275 5503 20281
rect 9300 20275 9312 20284
rect 9306 20272 9312 20275
rect 9364 20272 9370 20324
rect 10962 20272 10968 20324
rect 11020 20312 11026 20324
rect 11241 20315 11299 20321
rect 11241 20312 11253 20315
rect 11020 20284 11253 20312
rect 11020 20272 11026 20284
rect 11241 20281 11253 20284
rect 11287 20281 11299 20315
rect 11241 20275 11299 20281
rect 12253 20315 12311 20321
rect 12253 20281 12265 20315
rect 12299 20312 12311 20315
rect 13326 20315 13384 20321
rect 13326 20312 13338 20315
rect 12299 20284 13338 20312
rect 12299 20281 12311 20284
rect 12253 20275 12311 20281
rect 13326 20281 13338 20284
rect 13372 20312 13384 20315
rect 13446 20312 13452 20324
rect 13372 20284 13452 20312
rect 13372 20281 13384 20284
rect 13326 20275 13384 20281
rect 13446 20272 13452 20284
rect 13504 20272 13510 20324
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 3513 20247 3571 20253
rect 3513 20213 3525 20247
rect 3559 20244 3571 20247
rect 3878 20244 3884 20256
rect 3559 20216 3884 20244
rect 3559 20213 3571 20216
rect 3513 20207 3571 20213
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 3973 20247 4031 20253
rect 3973 20213 3985 20247
rect 4019 20244 4031 20247
rect 4062 20244 4068 20256
rect 4019 20216 4068 20244
rect 4019 20213 4031 20216
rect 3973 20207 4031 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4982 20244 4988 20256
rect 4943 20216 4988 20244
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 5074 20204 5080 20256
rect 5132 20244 5138 20256
rect 5353 20247 5411 20253
rect 5353 20244 5365 20247
rect 5132 20216 5365 20244
rect 5132 20204 5138 20216
rect 5353 20213 5365 20216
rect 5399 20213 5411 20247
rect 5353 20207 5411 20213
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10689 20247 10747 20253
rect 10689 20244 10701 20247
rect 9732 20216 10701 20244
rect 9732 20204 9738 20216
rect 10689 20213 10701 20216
rect 10735 20244 10747 20247
rect 11330 20244 11336 20256
rect 10735 20216 11336 20244
rect 10735 20213 10747 20216
rect 10689 20207 10747 20213
rect 11330 20204 11336 20216
rect 11388 20204 11394 20256
rect 15286 20244 15292 20256
rect 15247 20216 15292 20244
rect 15286 20204 15292 20216
rect 15344 20204 15350 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 2314 20040 2320 20052
rect 2275 20012 2320 20040
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 4709 20043 4767 20049
rect 4709 20009 4721 20043
rect 4755 20040 4767 20043
rect 4982 20040 4988 20052
rect 4755 20012 4988 20040
rect 4755 20009 4767 20012
rect 4709 20003 4767 20009
rect 4982 20000 4988 20012
rect 5040 20000 5046 20052
rect 6914 20040 6920 20052
rect 6875 20012 6920 20040
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 8260 20012 8493 20040
rect 8260 20000 8266 20012
rect 8481 20009 8493 20012
rect 8527 20040 8539 20043
rect 8846 20040 8852 20052
rect 8527 20012 8852 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9306 20040 9312 20052
rect 9171 20012 9312 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9306 20000 9312 20012
rect 9364 20040 9370 20052
rect 11057 20043 11115 20049
rect 11057 20040 11069 20043
rect 9364 20012 11069 20040
rect 9364 20000 9370 20012
rect 11057 20009 11069 20012
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 11204 20012 11713 20040
rect 11204 20000 11210 20012
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 12342 20000 12348 20052
rect 12400 20040 12406 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 12400 20012 13369 20040
rect 12400 20000 12406 20012
rect 13357 20009 13369 20012
rect 13403 20040 13415 20043
rect 13722 20040 13728 20052
rect 13403 20012 13728 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 5258 19932 5264 19984
rect 5316 19972 5322 19984
rect 5442 19981 5448 19984
rect 5436 19972 5448 19981
rect 5316 19944 5448 19972
rect 5316 19932 5322 19944
rect 5436 19935 5448 19944
rect 5442 19932 5448 19935
rect 5500 19932 5506 19984
rect 8570 19972 8576 19984
rect 7576 19944 8576 19972
rect 7576 19916 7604 19944
rect 8570 19932 8576 19944
rect 8628 19932 8634 19984
rect 9950 19981 9956 19984
rect 9944 19972 9956 19981
rect 9863 19944 9956 19972
rect 9944 19935 9956 19944
rect 10008 19972 10014 19984
rect 10778 19972 10784 19984
rect 10008 19944 10784 19972
rect 9950 19932 9956 19935
rect 10008 19932 10014 19944
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 11330 19972 11336 19984
rect 11291 19944 11336 19972
rect 11330 19932 11336 19944
rect 11388 19932 11394 19984
rect 15565 19975 15623 19981
rect 15565 19941 15577 19975
rect 15611 19972 15623 19975
rect 16022 19972 16028 19984
rect 15611 19944 16028 19972
rect 15611 19941 15623 19944
rect 15565 19935 15623 19941
rect 16022 19932 16028 19944
rect 16080 19932 16086 19984
rect 2222 19864 2228 19916
rect 2280 19904 2286 19916
rect 2685 19907 2743 19913
rect 2685 19904 2697 19907
rect 2280 19876 2697 19904
rect 2280 19864 2286 19876
rect 2685 19873 2697 19876
rect 2731 19873 2743 19907
rect 2685 19867 2743 19873
rect 4065 19907 4123 19913
rect 4065 19873 4077 19907
rect 4111 19904 4123 19907
rect 4154 19904 4160 19916
rect 4111 19876 4160 19904
rect 4111 19873 4123 19876
rect 4065 19867 4123 19873
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 7558 19904 7564 19916
rect 7471 19876 7564 19904
rect 7558 19864 7564 19876
rect 7616 19864 7622 19916
rect 8386 19904 8392 19916
rect 8347 19876 8392 19904
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 13630 19904 13636 19916
rect 13311 19876 13636 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 15252 19876 15301 19904
rect 15252 19864 15258 19876
rect 15289 19873 15301 19876
rect 15335 19904 15347 19907
rect 15654 19904 15660 19916
rect 15335 19876 15660 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15654 19864 15660 19876
rect 15712 19864 15718 19916
rect 2406 19796 2412 19848
rect 2464 19836 2470 19848
rect 2777 19839 2835 19845
rect 2777 19836 2789 19839
rect 2464 19808 2789 19836
rect 2464 19796 2470 19808
rect 2777 19805 2789 19808
rect 2823 19805 2835 19839
rect 2777 19799 2835 19805
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 3878 19836 3884 19848
rect 3791 19808 3884 19836
rect 2869 19799 2927 19805
rect 2498 19728 2504 19780
rect 2556 19768 2562 19780
rect 2884 19768 2912 19799
rect 3878 19796 3884 19808
rect 3936 19836 3942 19848
rect 5166 19836 5172 19848
rect 3936 19808 5172 19836
rect 3936 19796 3942 19808
rect 5166 19796 5172 19808
rect 5224 19796 5230 19848
rect 8665 19839 8723 19845
rect 8665 19805 8677 19839
rect 8711 19836 8723 19839
rect 9306 19836 9312 19848
rect 8711 19808 9312 19836
rect 8711 19805 8723 19808
rect 8665 19799 8723 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9674 19836 9680 19848
rect 9635 19808 9680 19836
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 11882 19836 11888 19848
rect 11843 19808 11888 19836
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 13446 19836 13452 19848
rect 13407 19808 13452 19836
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 2556 19740 2912 19768
rect 2556 19728 2562 19740
rect 3510 19728 3516 19780
rect 3568 19768 3574 19780
rect 4985 19771 5043 19777
rect 4985 19768 4997 19771
rect 3568 19740 4997 19768
rect 3568 19728 3574 19740
rect 4985 19737 4997 19740
rect 5031 19768 5043 19771
rect 5074 19768 5080 19780
rect 5031 19740 5080 19768
rect 5031 19737 5043 19740
rect 4985 19731 5043 19737
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 6638 19768 6644 19780
rect 6380 19740 6644 19768
rect 1673 19703 1731 19709
rect 1673 19669 1685 19703
rect 1719 19700 1731 19703
rect 1854 19700 1860 19712
rect 1719 19672 1860 19700
rect 1719 19669 1731 19672
rect 1673 19663 1731 19669
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2222 19700 2228 19712
rect 2183 19672 2228 19700
rect 2222 19660 2228 19672
rect 2280 19660 2286 19712
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3786 19700 3792 19712
rect 3467 19672 3792 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4120 19672 4261 19700
rect 4120 19660 4126 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4249 19663 4307 19669
rect 5534 19660 5540 19712
rect 5592 19700 5598 19712
rect 6380 19700 6408 19740
rect 6638 19728 6644 19740
rect 6696 19768 6702 19780
rect 7377 19771 7435 19777
rect 7377 19768 7389 19771
rect 6696 19740 7389 19768
rect 6696 19728 6702 19740
rect 7377 19737 7389 19740
rect 7423 19737 7435 19771
rect 7377 19731 7435 19737
rect 12897 19771 12955 19777
rect 12897 19737 12909 19771
rect 12943 19768 12955 19771
rect 14642 19768 14648 19780
rect 12943 19740 14648 19768
rect 12943 19737 12955 19740
rect 12897 19731 12955 19737
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 6546 19700 6552 19712
rect 5592 19672 6408 19700
rect 6507 19672 6552 19700
rect 5592 19660 5598 19672
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 7282 19700 7288 19712
rect 7243 19672 7288 19700
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7926 19700 7932 19712
rect 7887 19672 7932 19700
rect 7926 19660 7932 19672
rect 7984 19660 7990 19712
rect 9398 19700 9404 19712
rect 9359 19672 9404 19700
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 12434 19700 12440 19712
rect 11388 19672 12440 19700
rect 11388 19660 11394 19672
rect 12434 19660 12440 19672
rect 12492 19700 12498 19712
rect 13078 19700 13084 19712
rect 12492 19672 13084 19700
rect 12492 19660 12498 19672
rect 13078 19660 13084 19672
rect 13136 19700 13142 19712
rect 13909 19703 13967 19709
rect 13909 19700 13921 19703
rect 13136 19672 13921 19700
rect 13136 19660 13142 19672
rect 13909 19669 13921 19672
rect 13955 19669 13967 19703
rect 13909 19663 13967 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 5258 19456 5264 19508
rect 5316 19496 5322 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 5316 19468 5641 19496
rect 5316 19456 5322 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 5629 19459 5687 19465
rect 8389 19499 8447 19505
rect 8389 19465 8401 19499
rect 8435 19496 8447 19499
rect 8570 19496 8576 19508
rect 8435 19468 8576 19496
rect 8435 19465 8447 19468
rect 8389 19459 8447 19465
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 8941 19499 8999 19505
rect 8941 19465 8953 19499
rect 8987 19496 8999 19499
rect 9306 19496 9312 19508
rect 8987 19468 9312 19496
rect 8987 19465 8999 19468
rect 8941 19459 8999 19465
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 13446 19456 13452 19508
rect 13504 19496 13510 19508
rect 13814 19496 13820 19508
rect 13504 19468 13820 19496
rect 13504 19456 13510 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 15654 19496 15660 19508
rect 15615 19468 15660 19496
rect 15654 19456 15660 19468
rect 15712 19456 15718 19508
rect 6546 19428 6552 19440
rect 5276 19400 6552 19428
rect 5276 19372 5304 19400
rect 6546 19388 6552 19400
rect 6604 19388 6610 19440
rect 7926 19388 7932 19440
rect 7984 19428 7990 19440
rect 7984 19400 8524 19428
rect 7984 19388 7990 19400
rect 4982 19320 4988 19372
rect 5040 19360 5046 19372
rect 5077 19363 5135 19369
rect 5077 19360 5089 19363
rect 5040 19332 5089 19360
rect 5040 19320 5046 19332
rect 5077 19329 5089 19332
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 7282 19360 7288 19372
rect 5316 19332 5409 19360
rect 7243 19332 7288 19360
rect 5316 19320 5322 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 8386 19360 8392 19372
rect 7377 19323 7435 19329
rect 8312 19332 8392 19360
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 4154 19292 4160 19304
rect 4115 19264 4160 19292
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4525 19295 4583 19301
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5276 19292 5304 19320
rect 7392 19292 7420 19323
rect 4571 19264 5304 19292
rect 6932 19264 7420 19292
rect 8113 19295 8171 19301
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 6932 19236 6960 19264
rect 8113 19261 8125 19295
rect 8159 19292 8171 19295
rect 8312 19292 8340 19332
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8159 19264 8340 19292
rect 8496 19292 8524 19400
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 14608 19400 15240 19428
rect 14608 19388 14614 19400
rect 9582 19360 9588 19372
rect 9543 19332 9588 19360
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19329 11299 19363
rect 11241 19323 11299 19329
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8496 19264 8585 19292
rect 8159 19261 8171 19264
rect 8113 19255 8171 19261
rect 8573 19261 8585 19264
rect 8619 19292 8631 19295
rect 9214 19292 9220 19304
rect 8619 19264 9220 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 9398 19292 9404 19304
rect 9359 19264 9404 19292
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 9824 19264 10057 19292
rect 9824 19252 9830 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10045 19255 10103 19261
rect 11146 19252 11152 19304
rect 11204 19292 11210 19304
rect 11256 19292 11284 19323
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 15212 19369 15240 19400
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 14700 19332 15117 19360
rect 14700 19320 14706 19332
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 25038 19320 25044 19372
rect 25096 19360 25102 19372
rect 25314 19360 25320 19372
rect 25096 19332 25320 19360
rect 25096 19320 25102 19332
rect 25314 19320 25320 19332
rect 25372 19320 25378 19372
rect 11609 19295 11667 19301
rect 11609 19292 11621 19295
rect 11204 19264 11621 19292
rect 11204 19252 11210 19264
rect 11609 19261 11621 19264
rect 11655 19261 11667 19295
rect 11609 19255 11667 19261
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12342 19292 12348 19304
rect 12299 19264 12348 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 14458 19292 14464 19304
rect 12492 19264 12940 19292
rect 14419 19264 14464 19292
rect 12492 19252 12498 19264
rect 2498 19224 2504 19236
rect 2148 19196 2504 19224
rect 2148 19168 2176 19196
rect 2498 19184 2504 19196
rect 2556 19233 2562 19236
rect 2556 19227 2620 19233
rect 2556 19193 2574 19227
rect 2608 19193 2620 19227
rect 4982 19224 4988 19236
rect 4943 19196 4988 19224
rect 2556 19187 2620 19193
rect 2556 19184 2562 19187
rect 4982 19184 4988 19196
rect 5040 19184 5046 19236
rect 6273 19227 6331 19233
rect 6273 19193 6285 19227
rect 6319 19224 6331 19227
rect 6914 19224 6920 19236
rect 6319 19196 6920 19224
rect 6319 19193 6331 19196
rect 6273 19187 6331 19193
rect 6914 19184 6920 19196
rect 6972 19184 6978 19236
rect 9416 19224 9444 19252
rect 12912 19236 12940 19264
rect 14458 19252 14464 19264
rect 14516 19292 14522 19304
rect 15013 19295 15071 19301
rect 15013 19292 15025 19295
rect 14516 19264 15025 19292
rect 14516 19252 14522 19264
rect 15013 19261 15025 19264
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 10226 19224 10232 19236
rect 9416 19196 10232 19224
rect 10226 19184 10232 19196
rect 10284 19184 10290 19236
rect 10413 19227 10471 19233
rect 10413 19193 10425 19227
rect 10459 19193 10471 19227
rect 10686 19224 10692 19236
rect 10413 19187 10471 19193
rect 10612 19196 10692 19224
rect 1857 19159 1915 19165
rect 1857 19125 1869 19159
rect 1903 19156 1915 19159
rect 2130 19156 2136 19168
rect 1903 19128 2136 19156
rect 1903 19125 1915 19128
rect 1857 19119 1915 19125
rect 2130 19116 2136 19128
rect 2188 19116 2194 19168
rect 3050 19116 3056 19168
rect 3108 19156 3114 19168
rect 3697 19159 3755 19165
rect 3697 19156 3709 19159
rect 3108 19128 3709 19156
rect 3108 19116 3114 19128
rect 3697 19125 3709 19128
rect 3743 19156 3755 19159
rect 3970 19156 3976 19168
rect 3743 19128 3976 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 4614 19156 4620 19168
rect 4575 19128 4620 19156
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6512 19128 6561 19156
rect 6512 19116 6518 19128
rect 6549 19125 6561 19128
rect 6595 19125 6607 19159
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 6549 19119 6607 19125
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9490 19156 9496 19168
rect 9451 19128 9496 19156
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 10042 19116 10048 19168
rect 10100 19156 10106 19168
rect 10428 19156 10456 19187
rect 10612 19165 10640 19196
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 12526 19184 12532 19236
rect 12584 19224 12590 19236
rect 12682 19227 12740 19233
rect 12682 19224 12694 19227
rect 12584 19196 12694 19224
rect 12584 19184 12590 19196
rect 12682 19193 12694 19196
rect 12728 19193 12740 19227
rect 12682 19187 12740 19193
rect 12894 19184 12900 19236
rect 12952 19184 12958 19236
rect 10100 19128 10456 19156
rect 10597 19159 10655 19165
rect 10100 19116 10106 19128
rect 10597 19125 10609 19159
rect 10643 19125 10655 19159
rect 10962 19156 10968 19168
rect 10923 19128 10968 19156
rect 10597 19119 10655 19125
rect 10962 19116 10968 19128
rect 11020 19116 11026 19168
rect 11057 19159 11115 19165
rect 11057 19125 11069 19159
rect 11103 19156 11115 19159
rect 11330 19156 11336 19168
rect 11103 19128 11336 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 11330 19116 11336 19128
rect 11388 19116 11394 19168
rect 13630 19116 13636 19168
rect 13688 19156 13694 19168
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 13688 19128 14105 19156
rect 13688 19116 13694 19128
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 14642 19156 14648 19168
rect 14603 19128 14648 19156
rect 14093 19119 14151 19125
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2317 18955 2375 18961
rect 2317 18921 2329 18955
rect 2363 18952 2375 18955
rect 2406 18952 2412 18964
rect 2363 18924 2412 18952
rect 2363 18921 2375 18924
rect 2317 18915 2375 18921
rect 2406 18912 2412 18924
rect 2464 18912 2470 18964
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 4982 18952 4988 18964
rect 4755 18924 4988 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 6454 18912 6460 18964
rect 6512 18952 6518 18964
rect 7190 18952 7196 18964
rect 6512 18924 7196 18952
rect 6512 18912 6518 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 7558 18952 7564 18964
rect 7519 18924 7564 18952
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 8113 18955 8171 18961
rect 8113 18921 8125 18955
rect 8159 18952 8171 18955
rect 8202 18952 8208 18964
rect 8159 18924 8208 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9582 18952 9588 18964
rect 9171 18924 9588 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9582 18912 9588 18924
rect 9640 18952 9646 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 9640 18924 11897 18952
rect 9640 18912 9646 18924
rect 11885 18921 11897 18924
rect 11931 18952 11943 18955
rect 12526 18952 12532 18964
rect 11931 18924 12532 18952
rect 11931 18921 11943 18924
rect 11885 18915 11943 18921
rect 12526 18912 12532 18924
rect 12584 18912 12590 18964
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13173 18955 13231 18961
rect 13173 18952 13185 18955
rect 12860 18924 13185 18952
rect 12860 18912 12866 18924
rect 13173 18921 13185 18924
rect 13219 18952 13231 18955
rect 13262 18952 13268 18964
rect 13219 18924 13268 18952
rect 13219 18921 13231 18924
rect 13173 18915 13231 18921
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 13814 18952 13820 18964
rect 13775 18924 13820 18952
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14608 18924 14657 18952
rect 14608 18912 14614 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 2777 18887 2835 18893
rect 2777 18853 2789 18887
rect 2823 18884 2835 18887
rect 2958 18884 2964 18896
rect 2823 18856 2964 18884
rect 2823 18853 2835 18856
rect 2777 18847 2835 18853
rect 2958 18844 2964 18856
rect 3016 18844 3022 18896
rect 5804 18887 5862 18893
rect 5804 18853 5816 18887
rect 5850 18884 5862 18887
rect 5994 18884 6000 18896
rect 5850 18856 6000 18884
rect 5850 18853 5862 18856
rect 5804 18847 5862 18853
rect 5994 18844 6000 18856
rect 6052 18844 6058 18896
rect 9950 18884 9956 18896
rect 9911 18856 9956 18884
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 10192 18856 10333 18884
rect 10192 18844 10198 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 11330 18884 11336 18896
rect 10321 18847 10379 18853
rect 10612 18856 11336 18884
rect 2866 18816 2872 18828
rect 2827 18788 2872 18816
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 3878 18776 3884 18828
rect 3936 18816 3942 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3936 18788 4077 18816
rect 3936 18776 3942 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5442 18816 5448 18828
rect 5215 18788 5448 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 5537 18819 5595 18825
rect 5537 18785 5549 18819
rect 5583 18816 5595 18819
rect 6086 18816 6092 18828
rect 5583 18788 6092 18816
rect 5583 18785 5595 18788
rect 5537 18779 5595 18785
rect 1394 18748 1400 18760
rect 1355 18720 1400 18748
rect 1394 18708 1400 18720
rect 1452 18708 1458 18760
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 2961 18751 3019 18757
rect 2961 18748 2973 18751
rect 2832 18720 2973 18748
rect 2832 18708 2838 18720
rect 2961 18717 2973 18720
rect 3007 18717 3019 18751
rect 2961 18711 3019 18717
rect 5166 18640 5172 18692
rect 5224 18680 5230 18692
rect 5261 18683 5319 18689
rect 5261 18680 5273 18683
rect 5224 18652 5273 18680
rect 5224 18640 5230 18652
rect 5261 18649 5273 18652
rect 5307 18680 5319 18683
rect 5552 18680 5580 18779
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 7926 18776 7932 18828
rect 7984 18816 7990 18828
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 7984 18788 8309 18816
rect 7984 18776 7990 18788
rect 8297 18785 8309 18788
rect 8343 18816 8355 18819
rect 9030 18816 9036 18828
rect 8343 18788 9036 18816
rect 8343 18785 8355 18788
rect 8297 18779 8355 18785
rect 9030 18776 9036 18788
rect 9088 18776 9094 18828
rect 10042 18776 10048 18828
rect 10100 18816 10106 18828
rect 10612 18816 10640 18856
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 13081 18887 13139 18893
rect 13081 18884 13093 18887
rect 12400 18856 13093 18884
rect 12400 18844 12406 18856
rect 13081 18853 13093 18856
rect 13127 18884 13139 18887
rect 13354 18884 13360 18896
rect 13127 18856 13360 18884
rect 13127 18853 13139 18856
rect 13081 18847 13139 18853
rect 13354 18844 13360 18856
rect 13412 18844 13418 18896
rect 10100 18788 10640 18816
rect 10772 18819 10830 18825
rect 10100 18776 10106 18788
rect 10772 18785 10784 18819
rect 10818 18816 10830 18819
rect 11146 18816 11152 18828
rect 10818 18788 11152 18816
rect 10818 18785 10830 18788
rect 10772 18779 10830 18785
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 8478 18748 8484 18760
rect 8439 18720 8484 18748
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 10410 18748 10416 18760
rect 9732 18720 10416 18748
rect 9732 18708 9738 18720
rect 10410 18708 10416 18720
rect 10468 18748 10474 18760
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 10468 18720 10517 18748
rect 10468 18708 10474 18720
rect 10505 18717 10517 18720
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 13262 18708 13268 18760
rect 13320 18748 13326 18760
rect 13320 18720 13365 18748
rect 13320 18708 13326 18720
rect 5307 18652 5580 18680
rect 5307 18649 5319 18652
rect 5261 18643 5319 18649
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 1857 18615 1915 18621
rect 1857 18612 1869 18615
rect 1728 18584 1869 18612
rect 1728 18572 1734 18584
rect 1857 18581 1869 18584
rect 1903 18581 1915 18615
rect 3418 18612 3424 18624
rect 3379 18584 3424 18612
rect 1857 18575 1915 18581
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 3786 18612 3792 18624
rect 3747 18584 3792 18612
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 4246 18612 4252 18624
rect 4207 18584 4252 18612
rect 4246 18572 4252 18584
rect 4304 18572 4310 18624
rect 6914 18612 6920 18624
rect 6875 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7285 18615 7343 18621
rect 7285 18581 7297 18615
rect 7331 18612 7343 18615
rect 7374 18612 7380 18624
rect 7331 18584 7380 18612
rect 7331 18581 7343 18584
rect 7285 18575 7343 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 9490 18612 9496 18624
rect 9451 18584 9496 18612
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 12710 18612 12716 18624
rect 12671 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 2866 18368 2872 18420
rect 2924 18408 2930 18420
rect 3050 18408 3056 18420
rect 2924 18380 3056 18408
rect 2924 18368 2930 18380
rect 3050 18368 3056 18380
rect 3108 18408 3114 18420
rect 3329 18411 3387 18417
rect 3329 18408 3341 18411
rect 3108 18380 3341 18408
rect 3108 18368 3114 18380
rect 3329 18377 3341 18380
rect 3375 18377 3387 18411
rect 3329 18371 3387 18377
rect 6825 18411 6883 18417
rect 6825 18377 6837 18411
rect 6871 18408 6883 18411
rect 7282 18408 7288 18420
rect 6871 18380 7288 18408
rect 6871 18377 6883 18380
rect 6825 18371 6883 18377
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 7926 18408 7932 18420
rect 7887 18380 7932 18408
rect 7926 18368 7932 18380
rect 7984 18368 7990 18420
rect 8386 18408 8392 18420
rect 8347 18380 8392 18408
rect 8386 18368 8392 18380
rect 8444 18368 8450 18420
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9548 18380 10793 18408
rect 9548 18368 9554 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 10781 18371 10839 18377
rect 11348 18380 14289 18408
rect 5261 18343 5319 18349
rect 5261 18309 5273 18343
rect 5307 18309 5319 18343
rect 5261 18303 5319 18309
rect 5276 18272 5304 18303
rect 9766 18300 9772 18352
rect 9824 18340 9830 18352
rect 10413 18343 10471 18349
rect 10413 18340 10425 18343
rect 9824 18312 10425 18340
rect 9824 18300 9830 18312
rect 10413 18309 10425 18312
rect 10459 18340 10471 18343
rect 11054 18340 11060 18352
rect 10459 18312 11060 18340
rect 10459 18309 10471 18312
rect 10413 18303 10471 18309
rect 11054 18300 11060 18312
rect 11112 18300 11118 18352
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5276 18244 5641 18272
rect 5629 18241 5641 18244
rect 5675 18272 5687 18275
rect 5994 18272 6000 18284
rect 5675 18244 6000 18272
rect 5675 18241 5687 18244
rect 5629 18235 5687 18241
rect 5994 18232 6000 18244
rect 6052 18272 6058 18284
rect 7374 18272 7380 18284
rect 6052 18244 7380 18272
rect 6052 18232 6058 18244
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8941 18275 8999 18281
rect 8941 18272 8953 18275
rect 8352 18244 8953 18272
rect 8352 18232 8358 18244
rect 8941 18241 8953 18244
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 11146 18272 11152 18284
rect 10091 18244 11152 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 11146 18232 11152 18244
rect 11204 18272 11210 18284
rect 11348 18281 11376 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 12253 18343 12311 18349
rect 12253 18309 12265 18343
rect 12299 18340 12311 18343
rect 12342 18340 12348 18352
rect 12299 18312 12348 18340
rect 12299 18309 12311 18312
rect 12253 18303 12311 18309
rect 12342 18300 12348 18312
rect 12400 18340 12406 18352
rect 12526 18340 12532 18352
rect 12400 18312 12532 18340
rect 12400 18300 12406 18312
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 12802 18340 12808 18352
rect 12763 18312 12808 18340
rect 12802 18300 12808 18312
rect 12860 18300 12866 18352
rect 11333 18275 11391 18281
rect 11333 18272 11345 18275
rect 11204 18244 11345 18272
rect 11204 18232 11210 18244
rect 11333 18241 11345 18244
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 2314 18204 2320 18216
rect 1719 18176 2320 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 2314 18164 2320 18176
rect 2372 18204 2378 18216
rect 3881 18207 3939 18213
rect 3881 18204 3893 18207
rect 2372 18176 3893 18204
rect 2372 18164 2378 18176
rect 3881 18173 3893 18176
rect 3927 18204 3939 18207
rect 5166 18204 5172 18216
rect 3927 18176 5172 18204
rect 3927 18173 3939 18176
rect 3881 18167 3939 18173
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 8754 18204 8760 18216
rect 8715 18176 8760 18204
rect 8754 18164 8760 18176
rect 8812 18204 8818 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 8812 18176 9413 18204
rect 8812 18164 8818 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10689 18207 10747 18213
rect 10689 18204 10701 18207
rect 10192 18176 10701 18204
rect 10192 18164 10198 18176
rect 10689 18173 10701 18176
rect 10735 18173 10747 18207
rect 10689 18167 10747 18173
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 11514 18204 11520 18216
rect 11287 18176 11520 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 11514 18164 11520 18176
rect 11572 18204 11578 18216
rect 12710 18204 12716 18216
rect 11572 18176 12716 18204
rect 11572 18164 11578 18176
rect 12710 18164 12716 18176
rect 12768 18164 12774 18216
rect 12894 18204 12900 18216
rect 12807 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18204 12958 18216
rect 13722 18204 13728 18216
rect 12952 18176 13728 18204
rect 12952 18164 12958 18176
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 1946 18145 1952 18148
rect 1940 18136 1952 18145
rect 1907 18108 1952 18136
rect 1940 18099 1952 18108
rect 1946 18096 1952 18099
rect 2004 18096 2010 18148
rect 2958 18096 2964 18148
rect 3016 18136 3022 18148
rect 3697 18139 3755 18145
rect 3697 18136 3709 18139
rect 3016 18108 3709 18136
rect 3016 18096 3022 18108
rect 3697 18105 3709 18108
rect 3743 18105 3755 18139
rect 3697 18099 3755 18105
rect 3970 18096 3976 18148
rect 4028 18136 4034 18148
rect 4148 18139 4206 18145
rect 4148 18136 4160 18139
rect 4028 18108 4160 18136
rect 4028 18096 4034 18108
rect 4148 18105 4160 18108
rect 4194 18136 4206 18139
rect 4614 18136 4620 18148
rect 4194 18108 4620 18136
rect 4194 18105 4206 18108
rect 4148 18099 4206 18105
rect 4614 18096 4620 18108
rect 4672 18096 4678 18148
rect 6273 18139 6331 18145
rect 6273 18105 6285 18139
rect 6319 18136 6331 18139
rect 6362 18136 6368 18148
rect 6319 18108 6368 18136
rect 6319 18105 6331 18108
rect 6273 18099 6331 18105
rect 6362 18096 6368 18108
rect 6420 18136 6426 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 6420 18108 7297 18136
rect 6420 18096 6426 18108
rect 7285 18105 7297 18108
rect 7331 18136 7343 18139
rect 8662 18136 8668 18148
rect 7331 18108 8668 18136
rect 7331 18105 7343 18108
rect 7285 18099 7343 18105
rect 8662 18096 8668 18108
rect 8720 18096 8726 18148
rect 10410 18096 10416 18148
rect 10468 18096 10474 18148
rect 11885 18139 11943 18145
rect 11885 18105 11897 18139
rect 11931 18136 11943 18139
rect 13164 18139 13222 18145
rect 13164 18136 13176 18139
rect 11931 18108 13176 18136
rect 11931 18105 11943 18108
rect 11885 18099 11943 18105
rect 13164 18105 13176 18108
rect 13210 18136 13222 18139
rect 13262 18136 13268 18148
rect 13210 18108 13268 18136
rect 13210 18105 13222 18108
rect 13164 18099 13222 18105
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2314 18068 2320 18080
rect 2188 18040 2320 18068
rect 2188 18028 2194 18040
rect 2314 18028 2320 18040
rect 2372 18068 2378 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 2372 18040 3065 18068
rect 2372 18028 2378 18040
rect 3053 18037 3065 18040
rect 3099 18037 3111 18071
rect 6546 18068 6552 18080
rect 6507 18040 6552 18068
rect 3053 18031 3111 18037
rect 6546 18028 6552 18040
rect 6604 18068 6610 18080
rect 7193 18071 7251 18077
rect 7193 18068 7205 18071
rect 6604 18040 7205 18068
rect 6604 18028 6610 18040
rect 7193 18037 7205 18040
rect 7239 18037 7251 18071
rect 8294 18068 8300 18080
rect 8255 18040 8300 18068
rect 7193 18031 7251 18037
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8628 18040 8861 18068
rect 8628 18028 8634 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10428 18068 10456 18096
rect 10505 18071 10563 18077
rect 10505 18068 10517 18071
rect 10100 18040 10517 18068
rect 10100 18028 10106 18040
rect 10505 18037 10517 18040
rect 10551 18037 10563 18071
rect 10505 18031 10563 18037
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11149 18071 11207 18077
rect 11149 18068 11161 18071
rect 11112 18040 11161 18068
rect 11112 18028 11118 18040
rect 11149 18037 11161 18040
rect 11195 18068 11207 18071
rect 11422 18068 11428 18080
rect 11195 18040 11428 18068
rect 11195 18037 11207 18040
rect 11149 18031 11207 18037
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 14550 18068 14556 18080
rect 14511 18040 14556 18068
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2222 17824 2228 17876
rect 2280 17864 2286 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 2280 17836 2421 17864
rect 2280 17824 2286 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 2409 17827 2467 17833
rect 2682 17824 2688 17876
rect 2740 17824 2746 17876
rect 2869 17867 2927 17873
rect 2869 17833 2881 17867
rect 2915 17864 2927 17867
rect 3142 17864 3148 17876
rect 2915 17836 3148 17864
rect 2915 17833 2927 17836
rect 2869 17827 2927 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 4246 17864 4252 17876
rect 4207 17836 4252 17864
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 5813 17867 5871 17873
rect 5813 17833 5825 17867
rect 5859 17864 5871 17867
rect 6270 17864 6276 17876
rect 5859 17836 6276 17864
rect 5859 17833 5871 17836
rect 5813 17827 5871 17833
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 11146 17864 11152 17876
rect 11107 17836 11152 17864
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11514 17864 11520 17876
rect 11475 17836 11520 17864
rect 11514 17824 11520 17836
rect 11572 17824 11578 17876
rect 12989 17867 13047 17873
rect 12989 17833 13001 17867
rect 13035 17864 13047 17867
rect 13262 17864 13268 17876
rect 13035 17836 13268 17864
rect 13035 17833 13047 17836
rect 12989 17827 13047 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 13722 17864 13728 17876
rect 13635 17836 13728 17864
rect 13722 17824 13728 17836
rect 13780 17864 13786 17876
rect 14550 17864 14556 17876
rect 13780 17836 14556 17864
rect 13780 17824 13786 17836
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2700 17796 2728 17824
rect 1820 17768 2728 17796
rect 1820 17756 1826 17768
rect 3602 17756 3608 17808
rect 3660 17796 3666 17808
rect 5169 17799 5227 17805
rect 5169 17796 5181 17799
rect 3660 17768 5181 17796
rect 3660 17756 3666 17768
rect 5169 17765 5181 17768
rect 5215 17796 5227 17799
rect 5534 17796 5540 17808
rect 5215 17768 5540 17796
rect 5215 17765 5227 17768
rect 5169 17759 5227 17765
rect 5534 17756 5540 17768
rect 5592 17756 5598 17808
rect 6914 17756 6920 17808
rect 6972 17796 6978 17808
rect 7162 17799 7220 17805
rect 7162 17796 7174 17799
rect 6972 17768 7174 17796
rect 6972 17756 6978 17768
rect 7162 17765 7174 17768
rect 7208 17765 7220 17799
rect 7162 17759 7220 17765
rect 2682 17688 2688 17740
rect 2740 17728 2746 17740
rect 2777 17731 2835 17737
rect 2777 17728 2789 17731
rect 2740 17700 2789 17728
rect 2740 17688 2746 17700
rect 2777 17697 2789 17700
rect 2823 17697 2835 17731
rect 4062 17728 4068 17740
rect 4023 17700 4068 17728
rect 2777 17691 2835 17697
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 4982 17688 4988 17740
rect 5040 17728 5046 17740
rect 5721 17731 5779 17737
rect 5721 17728 5733 17731
rect 5040 17700 5733 17728
rect 5040 17688 5046 17700
rect 5721 17697 5733 17700
rect 5767 17697 5779 17731
rect 5721 17691 5779 17697
rect 6086 17688 6092 17740
rect 6144 17728 6150 17740
rect 7650 17728 7656 17740
rect 6144 17700 7656 17728
rect 6144 17688 6150 17700
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 3878 17660 3884 17672
rect 3839 17632 3884 17660
rect 2961 17623 3019 17629
rect 1412 17524 1440 17623
rect 1946 17592 1952 17604
rect 1859 17564 1952 17592
rect 1946 17552 1952 17564
rect 2004 17592 2010 17604
rect 2317 17595 2375 17601
rect 2317 17592 2329 17595
rect 2004 17564 2329 17592
rect 2004 17552 2010 17564
rect 2317 17561 2329 17564
rect 2363 17592 2375 17595
rect 2774 17592 2780 17604
rect 2363 17564 2780 17592
rect 2363 17561 2375 17564
rect 2317 17555 2375 17561
rect 2774 17552 2780 17564
rect 2832 17592 2838 17604
rect 2976 17592 3004 17623
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 5994 17660 6000 17672
rect 5955 17632 6000 17660
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 6932 17669 6960 17700
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 9950 17728 9956 17740
rect 9539 17700 9956 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 9950 17688 9956 17700
rect 10008 17728 10014 17740
rect 10413 17731 10471 17737
rect 10413 17728 10425 17731
rect 10008 17700 10425 17728
rect 10008 17688 10014 17700
rect 10413 17697 10425 17700
rect 10459 17697 10471 17731
rect 11865 17731 11923 17737
rect 11865 17728 11877 17731
rect 10413 17691 10471 17697
rect 11440 17700 11877 17728
rect 11440 17672 11468 17700
rect 11865 17697 11877 17700
rect 11911 17697 11923 17731
rect 11865 17691 11923 17697
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13817 17731 13875 17737
rect 13817 17728 13829 17731
rect 13136 17700 13829 17728
rect 13136 17688 13142 17700
rect 13817 17697 13829 17700
rect 13863 17728 13875 17731
rect 14642 17728 14648 17740
rect 13863 17700 14648 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 14642 17688 14648 17700
rect 14700 17688 14706 17740
rect 6917 17663 6975 17669
rect 6917 17629 6929 17663
rect 6963 17629 6975 17663
rect 6917 17623 6975 17629
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 10505 17663 10563 17669
rect 10505 17660 10517 17663
rect 9824 17632 10517 17660
rect 9824 17620 9830 17632
rect 10505 17629 10517 17632
rect 10551 17629 10563 17663
rect 10505 17623 10563 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17660 10747 17663
rect 11422 17660 11428 17672
rect 10735 17632 11428 17660
rect 10735 17629 10747 17632
rect 10689 17623 10747 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17629 11667 17663
rect 13998 17660 14004 17672
rect 13959 17632 14004 17660
rect 11609 17623 11667 17629
rect 2832 17564 3004 17592
rect 3513 17595 3571 17601
rect 2832 17552 2838 17564
rect 3513 17561 3525 17595
rect 3559 17592 3571 17595
rect 4062 17592 4068 17604
rect 3559 17564 4068 17592
rect 3559 17561 3571 17564
rect 3513 17555 3571 17561
rect 4062 17552 4068 17564
rect 4120 17552 4126 17604
rect 9674 17552 9680 17604
rect 9732 17592 9738 17604
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 9732 17564 10057 17592
rect 9732 17552 9738 17564
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 3326 17524 3332 17536
rect 1412 17496 3332 17524
rect 3326 17484 3332 17496
rect 3384 17484 3390 17536
rect 5350 17524 5356 17536
rect 5311 17496 5356 17524
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 6457 17527 6515 17533
rect 6457 17493 6469 17527
rect 6503 17524 6515 17527
rect 6822 17524 6828 17536
rect 6503 17496 6828 17524
rect 6503 17493 6515 17496
rect 6457 17487 6515 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8294 17524 8300 17536
rect 7892 17496 8300 17524
rect 7892 17484 7898 17496
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 8570 17524 8576 17536
rect 8531 17496 8576 17524
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 9033 17527 9091 17533
rect 9033 17493 9045 17527
rect 9079 17524 9091 17527
rect 9122 17524 9128 17536
rect 9079 17496 9128 17524
rect 9079 17493 9091 17496
rect 9033 17487 9091 17493
rect 9122 17484 9128 17496
rect 9180 17484 9186 17536
rect 9953 17527 10011 17533
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 10134 17524 10140 17536
rect 9999 17496 10140 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10134 17484 10140 17496
rect 10192 17484 10198 17536
rect 11624 17524 11652 17623
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 12894 17524 12900 17536
rect 11624 17496 12900 17524
rect 12894 17484 12900 17496
rect 12952 17484 12958 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17320 2467 17323
rect 3142 17320 3148 17332
rect 2455 17292 3148 17320
rect 2455 17289 2467 17292
rect 2409 17283 2467 17289
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 6270 17280 6276 17292
rect 6328 17320 6334 17332
rect 6638 17320 6644 17332
rect 6328 17292 6644 17320
rect 6328 17280 6334 17292
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 9214 17320 9220 17332
rect 8260 17292 9220 17320
rect 8260 17280 8266 17292
rect 9214 17280 9220 17292
rect 9272 17320 9278 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 9272 17292 9321 17320
rect 9272 17280 9278 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 11422 17320 11428 17332
rect 11383 17292 11428 17320
rect 9309 17283 9367 17289
rect 11422 17280 11428 17292
rect 11480 17320 11486 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 11480 17292 11713 17320
rect 11480 17280 11486 17292
rect 11701 17289 11713 17292
rect 11747 17320 11759 17323
rect 12069 17323 12127 17329
rect 12069 17320 12081 17323
rect 11747 17292 12081 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 12069 17289 12081 17292
rect 12115 17289 12127 17323
rect 13078 17320 13084 17332
rect 13039 17292 13084 17320
rect 12069 17283 12127 17289
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 6822 17212 6828 17264
rect 6880 17252 6886 17264
rect 7006 17252 7012 17264
rect 6880 17224 7012 17252
rect 6880 17212 6886 17224
rect 7006 17212 7012 17224
rect 7064 17252 7070 17264
rect 7469 17255 7527 17261
rect 7469 17252 7481 17255
rect 7064 17224 7481 17252
rect 7064 17212 7070 17224
rect 7469 17221 7481 17224
rect 7515 17252 7527 17255
rect 9122 17252 9128 17264
rect 7515 17224 9128 17252
rect 7515 17221 7527 17224
rect 7469 17215 7527 17221
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 23474 17212 23480 17264
rect 23532 17252 23538 17264
rect 24762 17252 24768 17264
rect 23532 17224 24768 17252
rect 23532 17212 23538 17224
rect 24762 17212 24768 17224
rect 24820 17212 24826 17264
rect 24854 17212 24860 17264
rect 24912 17252 24918 17264
rect 25958 17252 25964 17264
rect 24912 17224 25964 17252
rect 24912 17212 24918 17224
rect 25958 17212 25964 17224
rect 26016 17212 26022 17264
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17184 4767 17187
rect 5626 17184 5632 17196
rect 4755 17156 5632 17184
rect 4755 17153 4767 17156
rect 4709 17147 4767 17153
rect 5626 17144 5632 17156
rect 5684 17184 5690 17196
rect 5813 17187 5871 17193
rect 5813 17184 5825 17187
rect 5684 17156 5825 17184
rect 5684 17144 5690 17156
rect 5813 17153 5825 17156
rect 5859 17184 5871 17187
rect 5994 17184 6000 17196
rect 5859 17156 6000 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 5994 17144 6000 17156
rect 6052 17144 6058 17196
rect 10042 17184 10048 17196
rect 10003 17156 10048 17184
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 1578 17116 1584 17128
rect 1443 17088 1584 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1578 17076 1584 17088
rect 1636 17076 1642 17128
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 2590 17116 2596 17128
rect 2547 17088 2596 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 2590 17076 2596 17088
rect 2648 17076 2654 17128
rect 4982 17116 4988 17128
rect 2700 17088 4988 17116
rect 1486 17008 1492 17060
rect 1544 17048 1550 17060
rect 2700 17048 2728 17088
rect 4982 17076 4988 17088
rect 5040 17076 5046 17128
rect 5534 17116 5540 17128
rect 5495 17088 5540 17116
rect 5534 17076 5540 17088
rect 5592 17116 5598 17128
rect 6086 17116 6092 17128
rect 5592 17088 6092 17116
rect 5592 17076 5598 17088
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 10301 17119 10359 17125
rect 10301 17116 10313 17119
rect 10192 17088 10313 17116
rect 10192 17076 10198 17088
rect 10301 17085 10313 17088
rect 10347 17085 10359 17119
rect 10301 17079 10359 17085
rect 13541 17119 13599 17125
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 14550 17116 14556 17128
rect 13587 17088 14556 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 14550 17076 14556 17088
rect 14608 17076 14614 17128
rect 1544 17020 2728 17048
rect 2768 17051 2826 17057
rect 1544 17008 1550 17020
rect 2768 17017 2780 17051
rect 2814 17048 2826 17051
rect 3142 17048 3148 17060
rect 2814 17020 3148 17048
rect 2814 17017 2826 17020
rect 2768 17011 2826 17017
rect 3142 17008 3148 17020
rect 3200 17008 3206 17060
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 5629 17051 5687 17057
rect 5629 17048 5641 17051
rect 5132 17020 5641 17048
rect 5132 17008 5138 17020
rect 5629 17017 5641 17020
rect 5675 17017 5687 17051
rect 5629 17011 5687 17017
rect 8021 17051 8079 17057
rect 8021 17017 8033 17051
rect 8067 17017 8079 17051
rect 8021 17011 8079 17017
rect 13808 17051 13866 17057
rect 13808 17017 13820 17051
rect 13854 17017 13866 17051
rect 13808 17011 13866 17017
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16980 2099 16983
rect 2682 16980 2688 16992
rect 2087 16952 2688 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 2682 16940 2688 16952
rect 2740 16940 2746 16992
rect 3878 16980 3884 16992
rect 3839 16952 3884 16980
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 5166 16980 5172 16992
rect 5127 16952 5172 16980
rect 5166 16940 5172 16952
rect 5224 16940 5230 16992
rect 6546 16980 6552 16992
rect 6507 16952 6552 16980
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 6972 16952 7021 16980
rect 6972 16940 6978 16952
rect 7009 16949 7021 16952
rect 7055 16949 7067 16983
rect 7009 16943 7067 16949
rect 7466 16940 7472 16992
rect 7524 16980 7530 16992
rect 7837 16983 7895 16989
rect 7837 16980 7849 16983
rect 7524 16952 7849 16980
rect 7524 16940 7530 16952
rect 7837 16949 7849 16952
rect 7883 16980 7895 16983
rect 8036 16980 8064 17011
rect 12710 16980 12716 16992
rect 7883 16952 8064 16980
rect 12671 16952 12716 16980
rect 7883 16949 7895 16952
rect 7837 16943 7895 16949
rect 12710 16940 12716 16952
rect 12768 16940 12774 16992
rect 13449 16983 13507 16989
rect 13449 16949 13461 16983
rect 13495 16980 13507 16983
rect 13722 16980 13728 16992
rect 13495 16952 13728 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 13722 16940 13728 16952
rect 13780 16980 13786 16992
rect 13832 16980 13860 17011
rect 14918 16980 14924 16992
rect 13780 16952 13860 16980
rect 14879 16952 14924 16980
rect 13780 16940 13786 16952
rect 14918 16940 14924 16952
rect 14976 16940 14982 16992
rect 15194 16980 15200 16992
rect 15155 16952 15200 16980
rect 15194 16940 15200 16952
rect 15252 16940 15258 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 2041 16779 2099 16785
rect 2041 16776 2053 16779
rect 1452 16748 2053 16776
rect 1452 16736 1458 16748
rect 2041 16745 2053 16748
rect 2087 16776 2099 16779
rect 2406 16776 2412 16788
rect 2087 16748 2412 16776
rect 2087 16745 2099 16748
rect 2041 16739 2099 16745
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 2832 16748 2877 16776
rect 2832 16736 2838 16748
rect 3234 16736 3240 16788
rect 3292 16736 3298 16788
rect 3513 16779 3571 16785
rect 3513 16745 3525 16779
rect 3559 16776 3571 16779
rect 3878 16776 3884 16788
rect 3559 16748 3884 16776
rect 3559 16745 3571 16748
rect 3513 16739 3571 16745
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 4062 16776 4068 16788
rect 4023 16748 4068 16776
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 5166 16736 5172 16788
rect 5224 16776 5230 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 5224 16748 6285 16776
rect 5224 16736 5230 16748
rect 6273 16745 6285 16748
rect 6319 16776 6331 16779
rect 6546 16776 6552 16788
rect 6319 16748 6552 16776
rect 6319 16745 6331 16748
rect 6273 16739 6331 16745
rect 6546 16736 6552 16748
rect 6604 16736 6610 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 9766 16776 9772 16788
rect 9539 16748 9772 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 11609 16779 11667 16785
rect 11609 16745 11621 16779
rect 11655 16745 11667 16779
rect 11974 16776 11980 16788
rect 11935 16748 11980 16776
rect 11609 16739 11667 16745
rect 2682 16668 2688 16720
rect 2740 16668 2746 16720
rect 3252 16708 3280 16736
rect 4246 16708 4252 16720
rect 3252 16680 4252 16708
rect 4246 16668 4252 16680
rect 4304 16708 4310 16720
rect 4525 16711 4583 16717
rect 4525 16708 4537 16711
rect 4304 16680 4537 16708
rect 4304 16668 4310 16680
rect 4525 16677 4537 16680
rect 4571 16708 4583 16711
rect 4798 16708 4804 16720
rect 4571 16680 4804 16708
rect 4571 16677 4583 16680
rect 4525 16671 4583 16677
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 5074 16668 5080 16720
rect 5132 16708 5138 16720
rect 5261 16711 5319 16717
rect 5261 16708 5273 16711
rect 5132 16680 5273 16708
rect 5132 16668 5138 16680
rect 5261 16677 5273 16680
rect 5307 16677 5319 16711
rect 5261 16671 5319 16677
rect 5350 16668 5356 16720
rect 5408 16708 5414 16720
rect 6365 16711 6423 16717
rect 6365 16708 6377 16711
rect 5408 16680 6377 16708
rect 5408 16668 5414 16680
rect 6365 16677 6377 16680
rect 6411 16708 6423 16711
rect 6917 16711 6975 16717
rect 6917 16708 6929 16711
rect 6411 16680 6929 16708
rect 6411 16677 6423 16680
rect 6365 16671 6423 16677
rect 6917 16677 6929 16680
rect 6963 16677 6975 16711
rect 8294 16708 8300 16720
rect 6917 16671 6975 16677
rect 7116 16680 8300 16708
rect 1762 16640 1768 16652
rect 1688 16612 1768 16640
rect 1688 16513 1716 16612
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2700 16640 2728 16668
rect 2700 16612 3188 16640
rect 1854 16532 1860 16584
rect 1912 16572 1918 16584
rect 2133 16575 2191 16581
rect 2133 16572 2145 16575
rect 1912 16544 2145 16572
rect 1912 16532 1918 16544
rect 2133 16541 2145 16544
rect 2179 16541 2191 16575
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2133 16535 2191 16541
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 3160 16572 3188 16612
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3292 16612 3801 16640
rect 3292 16600 3298 16612
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 5626 16640 5632 16652
rect 5587 16612 5632 16640
rect 3789 16603 3847 16609
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 5902 16600 5908 16652
rect 5960 16600 5966 16652
rect 7116 16649 7144 16680
rect 8294 16668 8300 16680
rect 8352 16668 8358 16720
rect 9784 16708 9812 16736
rect 11624 16708 11652 16739
rect 11974 16736 11980 16748
rect 12032 16736 12038 16788
rect 12066 16736 12072 16788
rect 12124 16776 12130 16788
rect 13173 16779 13231 16785
rect 13173 16776 13185 16779
rect 12124 16748 13185 16776
rect 12124 16736 12130 16748
rect 13173 16745 13185 16748
rect 13219 16745 13231 16779
rect 13173 16739 13231 16745
rect 13538 16736 13544 16788
rect 13596 16776 13602 16788
rect 13633 16779 13691 16785
rect 13633 16776 13645 16779
rect 13596 16748 13645 16776
rect 13596 16736 13602 16748
rect 13633 16745 13645 16748
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 14550 16736 14556 16788
rect 14608 16776 14614 16788
rect 14645 16779 14703 16785
rect 14645 16776 14657 16779
rect 14608 16748 14657 16776
rect 14608 16736 14614 16748
rect 14645 16745 14657 16748
rect 14691 16776 14703 16779
rect 15194 16776 15200 16788
rect 14691 16748 15200 16776
rect 14691 16745 14703 16748
rect 14645 16739 14703 16745
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 9784 16680 11652 16708
rect 12710 16668 12716 16720
rect 12768 16708 12774 16720
rect 14185 16711 14243 16717
rect 14185 16708 14197 16711
rect 12768 16680 14197 16708
rect 12768 16668 12774 16680
rect 14185 16677 14197 16680
rect 14231 16677 14243 16711
rect 14185 16671 14243 16677
rect 15565 16711 15623 16717
rect 15565 16677 15577 16711
rect 15611 16708 15623 16711
rect 16114 16708 16120 16720
rect 15611 16680 16120 16708
rect 15611 16677 15623 16680
rect 15565 16671 15623 16677
rect 16114 16668 16120 16680
rect 16172 16668 16178 16720
rect 7101 16643 7159 16649
rect 7101 16609 7113 16643
rect 7147 16609 7159 16643
rect 7650 16640 7656 16652
rect 7611 16612 7656 16640
rect 7101 16603 7159 16609
rect 7650 16600 7656 16612
rect 7708 16600 7714 16652
rect 7742 16600 7748 16652
rect 7800 16640 7806 16652
rect 7909 16643 7967 16649
rect 7909 16640 7921 16643
rect 7800 16612 7921 16640
rect 7800 16600 7806 16612
rect 7909 16609 7921 16612
rect 7955 16609 7967 16643
rect 10318 16640 10324 16652
rect 10279 16612 10324 16640
rect 7909 16603 7967 16609
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 12618 16640 12624 16652
rect 12579 16612 12624 16640
rect 12618 16600 12624 16612
rect 12676 16600 12682 16652
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16640 13599 16643
rect 13630 16640 13636 16652
rect 13587 16612 13636 16640
rect 13587 16609 13599 16612
rect 13541 16603 13599 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 15286 16640 15292 16652
rect 15247 16612 15292 16640
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 4522 16572 4528 16584
rect 3160 16544 4528 16572
rect 4522 16532 4528 16544
rect 4580 16532 4586 16584
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 5166 16572 5172 16584
rect 4755 16544 5172 16572
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 1673 16507 1731 16513
rect 1673 16473 1685 16507
rect 1719 16473 1731 16507
rect 1673 16467 1731 16473
rect 3142 16436 3148 16448
rect 3055 16408 3148 16436
rect 3142 16396 3148 16408
rect 3200 16436 3206 16448
rect 4724 16436 4752 16535
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5920 16513 5948 16600
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6457 16575 6515 16581
rect 6457 16572 6469 16575
rect 6328 16544 6469 16572
rect 6328 16532 6334 16544
rect 6457 16541 6469 16544
rect 6503 16572 6515 16575
rect 6822 16572 6828 16584
rect 6503 16544 6828 16572
rect 6503 16541 6515 16544
rect 6457 16535 6515 16541
rect 6822 16532 6828 16544
rect 6880 16532 6886 16584
rect 7282 16572 7288 16584
rect 7243 16544 7288 16572
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 9858 16532 9864 16584
rect 9916 16572 9922 16584
rect 10413 16575 10471 16581
rect 10413 16572 10425 16575
rect 9916 16544 10425 16572
rect 9916 16532 9922 16544
rect 10413 16541 10425 16544
rect 10459 16541 10471 16575
rect 10413 16535 10471 16541
rect 10505 16575 10563 16581
rect 10505 16541 10517 16575
rect 10551 16541 10563 16575
rect 12066 16572 12072 16584
rect 12027 16544 12072 16572
rect 10505 16535 10563 16541
rect 5905 16507 5963 16513
rect 5905 16473 5917 16507
rect 5951 16473 5963 16507
rect 5905 16467 5963 16473
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 10520 16504 10548 16535
rect 12066 16532 12072 16544
rect 12124 16532 12130 16584
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 13722 16572 13728 16584
rect 12216 16544 12309 16572
rect 13683 16544 13728 16572
rect 12216 16532 12222 16544
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 12176 16504 12204 16532
rect 10192 16476 12204 16504
rect 10192 16464 10198 16476
rect 9030 16436 9036 16448
rect 3200 16408 4752 16436
rect 8991 16408 9036 16436
rect 3200 16396 3206 16408
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 11054 16436 11060 16448
rect 11015 16408 11060 16436
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11333 16439 11391 16445
rect 11333 16436 11345 16439
rect 11296 16408 11345 16436
rect 11296 16396 11302 16408
rect 11333 16405 11345 16408
rect 11379 16405 11391 16439
rect 13078 16436 13084 16448
rect 13039 16408 13084 16436
rect 11333 16399 11391 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2406 16192 2412 16244
rect 2464 16232 2470 16244
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2464 16204 2605 16232
rect 2464 16192 2470 16204
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 4525 16235 4583 16241
rect 4525 16232 4537 16235
rect 2593 16195 2651 16201
rect 2976 16204 4537 16232
rect 2038 16096 2044 16108
rect 1999 16068 2044 16096
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 2976 16105 3004 16204
rect 4525 16201 4537 16204
rect 4571 16232 4583 16235
rect 5074 16232 5080 16244
rect 4571 16204 5080 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 5166 16192 5172 16244
rect 5224 16232 5230 16244
rect 5629 16235 5687 16241
rect 5629 16232 5641 16235
rect 5224 16204 5641 16232
rect 5224 16192 5230 16204
rect 5629 16201 5641 16204
rect 5675 16232 5687 16235
rect 5994 16232 6000 16244
rect 5675 16204 6000 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6270 16232 6276 16244
rect 6231 16204 6276 16232
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 8573 16235 8631 16241
rect 8573 16232 8585 16235
rect 8352 16204 8585 16232
rect 8352 16192 8358 16204
rect 8573 16201 8585 16204
rect 8619 16201 8631 16235
rect 8573 16195 8631 16201
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 10318 16232 10324 16244
rect 9916 16204 10324 16232
rect 9916 16192 9922 16204
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 11974 16232 11980 16244
rect 11931 16204 11980 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 13722 16232 13728 16244
rect 12299 16204 13728 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 13722 16192 13728 16204
rect 13780 16232 13786 16244
rect 14369 16235 14427 16241
rect 14369 16232 14381 16235
rect 13780 16204 14381 16232
rect 13780 16192 13786 16204
rect 14369 16201 14381 16204
rect 14415 16201 14427 16235
rect 14369 16195 14427 16201
rect 4798 16164 4804 16176
rect 4759 16136 4804 16164
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 9950 16164 9956 16176
rect 9911 16136 9956 16164
rect 9950 16124 9956 16136
rect 10008 16124 10014 16176
rect 2225 16099 2283 16105
rect 2225 16065 2237 16099
rect 2271 16096 2283 16099
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2271 16068 2973 16096
rect 2271 16065 2283 16068
rect 2225 16059 2283 16065
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 2961 16059 3019 16065
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4706 16096 4712 16108
rect 4580 16068 4712 16096
rect 4580 16056 4586 16068
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4764 16068 5181 16096
rect 4764 16056 4770 16068
rect 5169 16065 5181 16068
rect 5215 16065 5227 16099
rect 5169 16059 5227 16065
rect 5721 16099 5779 16105
rect 5721 16065 5733 16099
rect 5767 16096 5779 16099
rect 6454 16096 6460 16108
rect 5767 16068 6460 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 9306 16096 9312 16108
rect 9267 16068 9312 16096
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11333 16099 11391 16105
rect 11333 16096 11345 16099
rect 11112 16068 11345 16096
rect 11112 16056 11118 16068
rect 11333 16065 11345 16068
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16096 15807 16099
rect 16482 16096 16488 16108
rect 15795 16068 16488 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 2056 16028 2084 16056
rect 2682 16028 2688 16040
rect 2056 16000 2688 16028
rect 2682 15988 2688 16000
rect 2740 15988 2746 16040
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 3418 16037 3424 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 2832 16000 3157 16028
rect 2832 15988 2838 16000
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3412 16028 3424 16037
rect 3331 16000 3424 16028
rect 3145 15991 3203 15997
rect 3412 15991 3424 16000
rect 3476 16028 3482 16040
rect 3878 16028 3884 16040
rect 3476 16000 3884 16028
rect 3160 15960 3188 15991
rect 3418 15988 3424 15991
rect 3476 15988 3482 16000
rect 3878 15988 3884 16000
rect 3936 15988 3942 16040
rect 5810 15988 5816 16040
rect 5868 16028 5874 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 5868 16000 6929 16028
rect 5868 15988 5874 16000
rect 6917 15997 6929 16000
rect 6963 16028 6975 16031
rect 7006 16028 7012 16040
rect 6963 16000 7012 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 9125 16031 9183 16037
rect 9125 15997 9137 16031
rect 9171 16028 9183 16031
rect 9582 16028 9588 16040
rect 9171 16000 9588 16028
rect 9171 15997 9183 16000
rect 9125 15991 9183 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10686 16028 10692 16040
rect 9824 16000 10692 16028
rect 9824 15988 9830 16000
rect 10686 15988 10692 16000
rect 10744 15988 10750 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11238 16028 11244 16040
rect 11020 16000 11244 16028
rect 11020 15988 11026 16000
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 3786 15960 3792 15972
rect 3160 15932 3792 15960
rect 3786 15920 3792 15932
rect 3844 15920 3850 15972
rect 7162 15963 7220 15969
rect 7162 15960 7174 15963
rect 7024 15932 7174 15960
rect 7024 15904 7052 15932
rect 7162 15929 7174 15932
rect 7208 15929 7220 15963
rect 10870 15960 10876 15972
rect 7162 15923 7220 15929
rect 9876 15932 10876 15960
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 1949 15895 2007 15901
rect 1949 15861 1961 15895
rect 1995 15892 2007 15895
rect 3510 15892 3516 15904
rect 1995 15864 3516 15892
rect 1995 15861 2007 15864
rect 1949 15855 2007 15861
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 6641 15895 6699 15901
rect 6641 15861 6653 15895
rect 6687 15892 6699 15895
rect 7006 15892 7012 15904
rect 6687 15864 7012 15892
rect 6687 15861 6699 15864
rect 6641 15855 6699 15861
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 8297 15895 8355 15901
rect 8297 15861 8309 15895
rect 8343 15892 8355 15895
rect 8386 15892 8392 15904
rect 8343 15864 8392 15892
rect 8343 15861 8355 15864
rect 8297 15855 8355 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 9033 15895 9091 15901
rect 9033 15861 9045 15895
rect 9079 15892 9091 15895
rect 9876 15892 9904 15932
rect 10870 15920 10876 15932
rect 10928 15960 10934 15972
rect 11149 15963 11207 15969
rect 11149 15960 11161 15963
rect 10928 15932 11161 15960
rect 10928 15920 10934 15932
rect 11149 15929 11161 15932
rect 11195 15929 11207 15963
rect 11348 15960 11376 16059
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12989 16031 13047 16037
rect 12989 16028 13001 16031
rect 12492 16000 13001 16028
rect 12492 15988 12498 16000
rect 12989 15997 13001 16000
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13630 15988 13636 16040
rect 13688 16028 13694 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 13688 16000 14657 16028
rect 13688 15988 13694 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 15286 16028 15292 16040
rect 15247 16000 15292 16028
rect 14645 15991 14703 15997
rect 15286 15988 15292 16000
rect 15344 15988 15350 16040
rect 15470 16028 15476 16040
rect 15431 16000 15476 16028
rect 15470 15988 15476 16000
rect 15528 16028 15534 16040
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15528 16000 16221 16028
rect 15528 15988 15534 16000
rect 16209 15997 16221 16000
rect 16255 15997 16267 16031
rect 16209 15991 16267 15997
rect 13078 15960 13084 15972
rect 11348 15932 13084 15960
rect 11149 15923 11207 15929
rect 13078 15920 13084 15932
rect 13136 15960 13142 15972
rect 13256 15963 13314 15969
rect 13256 15960 13268 15963
rect 13136 15932 13268 15960
rect 13136 15920 13142 15932
rect 13256 15929 13268 15932
rect 13302 15960 13314 15963
rect 13814 15960 13820 15972
rect 13302 15932 13820 15960
rect 13302 15929 13314 15932
rect 13256 15923 13314 15929
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 9079 15864 9904 15892
rect 9079 15861 9091 15864
rect 9033 15855 9091 15861
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10505 15895 10563 15901
rect 10505 15892 10517 15895
rect 10100 15864 10517 15892
rect 10100 15852 10106 15864
rect 10505 15861 10517 15864
rect 10551 15861 10563 15895
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10505 15855 10563 15861
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13538 15892 13544 15904
rect 12943 15864 13544 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13538 15852 13544 15864
rect 13596 15852 13602 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2314 15688 2320 15700
rect 2275 15660 2320 15688
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3384 15660 3801 15688
rect 3384 15648 3390 15660
rect 3789 15657 3801 15660
rect 3835 15688 3847 15691
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 3835 15660 4445 15688
rect 3835 15657 3847 15660
rect 3789 15651 3847 15657
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 5074 15688 5080 15700
rect 5035 15660 5080 15688
rect 4433 15651 4491 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 7742 15688 7748 15700
rect 7703 15660 7748 15688
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 8113 15691 8171 15697
rect 8113 15657 8125 15691
rect 8159 15688 8171 15691
rect 8202 15688 8208 15700
rect 8159 15660 8208 15688
rect 8159 15657 8171 15660
rect 8113 15651 8171 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 9493 15691 9551 15697
rect 9493 15657 9505 15691
rect 9539 15688 9551 15691
rect 9582 15688 9588 15700
rect 9539 15660 9588 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 9858 15688 9864 15700
rect 9819 15660 9864 15688
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10192 15660 10333 15688
rect 10192 15648 10198 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10870 15688 10876 15700
rect 10831 15660 10876 15688
rect 10321 15651 10379 15657
rect 3418 15620 3424 15632
rect 3379 15592 3424 15620
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 10336 15620 10364 15651
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12253 15691 12311 15697
rect 12253 15688 12265 15691
rect 12124 15660 12265 15688
rect 12124 15648 12130 15660
rect 12253 15657 12265 15660
rect 12299 15657 12311 15691
rect 13814 15688 13820 15700
rect 13775 15660 13820 15688
rect 12253 15651 12311 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 11977 15623 12035 15629
rect 11977 15620 11989 15623
rect 10336 15592 11989 15620
rect 11977 15589 11989 15592
rect 12023 15589 12035 15623
rect 11977 15583 12035 15589
rect 16298 15580 16304 15632
rect 16356 15620 16362 15632
rect 16393 15623 16451 15629
rect 16393 15620 16405 15623
rect 16356 15592 16405 15620
rect 16356 15580 16362 15592
rect 16393 15589 16405 15592
rect 16439 15589 16451 15623
rect 16393 15583 16451 15589
rect 2774 15512 2780 15564
rect 2832 15552 2838 15564
rect 3436 15552 3464 15580
rect 2832 15524 2877 15552
rect 3436 15524 4660 15552
rect 2832 15512 2838 15524
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 1854 15484 1860 15496
rect 1815 15456 1860 15484
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 2590 15444 2596 15496
rect 2648 15484 2654 15496
rect 2869 15487 2927 15493
rect 2869 15484 2881 15487
rect 2648 15456 2881 15484
rect 2648 15444 2654 15456
rect 2869 15453 2881 15456
rect 2915 15453 2927 15487
rect 2869 15447 2927 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3142 15484 3148 15496
rect 3007 15456 3148 15484
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 2884 15416 2912 15447
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4632 15493 4660 15524
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5721 15555 5779 15561
rect 5721 15552 5733 15555
rect 5592 15524 5733 15552
rect 5592 15512 5598 15524
rect 5721 15521 5733 15524
rect 5767 15552 5779 15555
rect 5810 15552 5816 15564
rect 5767 15524 5816 15552
rect 5767 15521 5779 15524
rect 5721 15515 5779 15521
rect 5810 15512 5816 15524
rect 5868 15512 5874 15564
rect 5994 15561 6000 15564
rect 5988 15552 6000 15561
rect 5955 15524 6000 15552
rect 5988 15515 6000 15524
rect 5994 15512 6000 15515
rect 6052 15512 6058 15564
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15552 8355 15555
rect 8570 15552 8576 15564
rect 8343 15524 8576 15552
rect 8343 15521 8355 15524
rect 8297 15515 8355 15521
rect 8570 15512 8576 15524
rect 8628 15552 8634 15564
rect 10778 15552 10784 15564
rect 8628 15524 10784 15552
rect 8628 15512 8634 15524
rect 10778 15512 10784 15524
rect 10836 15512 10842 15564
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15552 11299 15555
rect 11882 15552 11888 15564
rect 11287 15524 11888 15552
rect 11287 15521 11299 15524
rect 11241 15515 11299 15521
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 12693 15555 12751 15561
rect 12693 15552 12705 15555
rect 11992 15524 12705 15552
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4212 15456 4537 15484
rect 4212 15444 4218 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 8478 15484 8484 15496
rect 8439 15456 8484 15484
rect 4617 15447 4675 15453
rect 8478 15444 8484 15456
rect 8536 15444 8542 15496
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11330 15484 11336 15496
rect 10744 15456 11336 15484
rect 10744 15444 10750 15456
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11422 15444 11428 15496
rect 11480 15484 11486 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11480 15456 11529 15484
rect 11480 15444 11486 15456
rect 11517 15453 11529 15456
rect 11563 15484 11575 15487
rect 11992 15484 12020 15524
rect 12693 15521 12705 15524
rect 12739 15552 12751 15555
rect 13814 15552 13820 15564
rect 12739 15524 13820 15552
rect 12739 15521 12751 15524
rect 12693 15515 12751 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 16114 15552 16120 15564
rect 16075 15524 16120 15552
rect 16114 15512 16120 15524
rect 16172 15512 16178 15564
rect 11563 15456 12020 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12492 15456 12537 15484
rect 12492 15444 12498 15456
rect 3050 15416 3056 15428
rect 2884 15388 3056 15416
rect 3050 15376 3056 15388
rect 3108 15376 3114 15428
rect 3510 15376 3516 15428
rect 3568 15416 3574 15428
rect 4065 15419 4123 15425
rect 4065 15416 4077 15419
rect 3568 15388 4077 15416
rect 3568 15376 3574 15388
rect 4065 15385 4077 15388
rect 4111 15385 4123 15419
rect 4065 15379 4123 15385
rect 10781 15419 10839 15425
rect 10781 15385 10793 15419
rect 10827 15416 10839 15419
rect 11440 15416 11468 15444
rect 10827 15388 11468 15416
rect 10827 15385 10839 15388
rect 10781 15379 10839 15385
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15348 2467 15351
rect 3234 15348 3240 15360
rect 2455 15320 3240 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 5537 15351 5595 15357
rect 5537 15348 5549 15351
rect 5500 15320 5549 15348
rect 5500 15308 5506 15320
rect 5537 15317 5549 15320
rect 5583 15317 5595 15351
rect 5537 15311 5595 15317
rect 7101 15351 7159 15357
rect 7101 15317 7113 15351
rect 7147 15348 7159 15351
rect 7374 15348 7380 15360
rect 7147 15320 7380 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 9122 15348 9128 15360
rect 9083 15320 9128 15348
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 14182 15348 14188 15360
rect 14143 15320 14188 15348
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 1581 15147 1639 15153
rect 1581 15144 1593 15147
rect 1544 15116 1593 15144
rect 1544 15104 1550 15116
rect 1581 15113 1593 15116
rect 1627 15113 1639 15147
rect 1581 15107 1639 15113
rect 2682 15104 2688 15156
rect 2740 15144 2746 15156
rect 2777 15147 2835 15153
rect 2777 15144 2789 15147
rect 2740 15116 2789 15144
rect 2740 15104 2746 15116
rect 2777 15113 2789 15116
rect 2823 15113 2835 15147
rect 5534 15144 5540 15156
rect 2777 15107 2835 15113
rect 4448 15116 5540 15144
rect 3234 15008 3240 15020
rect 3195 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 14968 3298 15020
rect 3418 15008 3424 15020
rect 3379 14980 3424 15008
rect 3418 14968 3424 14980
rect 3476 14968 3482 15020
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 4448 15017 4476 15116
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9033 15147 9091 15153
rect 9033 15144 9045 15147
rect 8352 15116 9045 15144
rect 8352 15104 8358 15116
rect 9033 15113 9045 15116
rect 9079 15113 9091 15147
rect 10686 15144 10692 15156
rect 10647 15116 10692 15144
rect 9033 15107 9091 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 10962 15144 10968 15156
rect 10827 15116 10968 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 13814 15144 13820 15156
rect 13775 15116 13820 15144
rect 13814 15104 13820 15116
rect 13872 15144 13878 15156
rect 14093 15147 14151 15153
rect 14093 15144 14105 15147
rect 13872 15116 14105 15144
rect 13872 15104 13878 15116
rect 14093 15113 14105 15116
rect 14139 15113 14151 15147
rect 14093 15107 14151 15113
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 14240 15116 14473 15144
rect 14240 15104 14246 15116
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 14461 15107 14519 15113
rect 8570 15076 8576 15088
rect 8531 15048 8576 15076
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 16114 15076 16120 15088
rect 16075 15048 16120 15076
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 3844 14980 4445 15008
rect 3844 14968 3850 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 8941 15011 8999 15017
rect 8941 14977 8953 15011
rect 8987 15008 8999 15011
rect 9582 15008 9588 15020
rect 8987 14980 9588 15008
rect 8987 14977 8999 14980
rect 8941 14971 8999 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 11422 15008 11428 15020
rect 11383 14980 11428 15008
rect 11422 14968 11428 14980
rect 11480 14968 11486 15020
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 3145 14943 3203 14949
rect 1443 14912 3096 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2133 14875 2191 14881
rect 2133 14841 2145 14875
rect 2179 14872 2191 14875
rect 2682 14872 2688 14884
rect 2179 14844 2688 14872
rect 2179 14841 2191 14844
rect 2133 14835 2191 14841
rect 2682 14832 2688 14844
rect 2740 14832 2746 14884
rect 3068 14872 3096 14912
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 4062 14940 4068 14952
rect 3191 14912 4068 14940
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 4700 14943 4758 14949
rect 4700 14909 4712 14943
rect 4746 14940 4758 14943
rect 5074 14940 5080 14952
rect 4746 14912 5080 14940
rect 4746 14909 4758 14912
rect 4700 14903 4758 14909
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 6822 14940 6828 14952
rect 6783 14912 6828 14940
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 9180 14912 9413 14940
rect 9180 14900 9186 14912
rect 9401 14909 9413 14912
rect 9447 14940 9459 14943
rect 9674 14940 9680 14952
rect 9447 14912 9680 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9674 14900 9680 14912
rect 9732 14900 9738 14952
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 12434 14940 12440 14952
rect 12032 14912 12440 14940
rect 12032 14900 12038 14912
rect 12434 14900 12440 14912
rect 12492 14940 12498 14952
rect 12492 14912 12537 14940
rect 12492 14900 12498 14912
rect 3694 14872 3700 14884
rect 3068 14844 3700 14872
rect 3694 14832 3700 14844
rect 3752 14832 3758 14884
rect 4798 14832 4804 14884
rect 4856 14872 4862 14884
rect 6641 14875 6699 14881
rect 4856 14844 6500 14872
rect 4856 14832 4862 14844
rect 1854 14764 1860 14816
rect 1912 14804 1918 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 1912 14776 2421 14804
rect 1912 14764 1918 14776
rect 2409 14773 2421 14776
rect 2455 14804 2467 14807
rect 2590 14804 2596 14816
rect 2455 14776 2596 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 4154 14804 4160 14816
rect 4115 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 5810 14804 5816 14816
rect 5771 14776 5816 14804
rect 5810 14764 5816 14776
rect 5868 14804 5874 14816
rect 5994 14804 6000 14816
rect 5868 14776 6000 14804
rect 5868 14764 5874 14776
rect 5994 14764 6000 14776
rect 6052 14804 6058 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 6052 14776 6193 14804
rect 6052 14764 6058 14776
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6472 14804 6500 14844
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7092 14875 7150 14881
rect 7092 14872 7104 14875
rect 6687 14844 7104 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7092 14841 7104 14844
rect 7138 14872 7150 14875
rect 7374 14872 7380 14884
rect 7138 14844 7380 14872
rect 7138 14841 7150 14844
rect 7092 14835 7150 14841
rect 7374 14832 7380 14844
rect 7432 14832 7438 14884
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 12682 14875 12740 14881
rect 12682 14872 12694 14875
rect 12299 14844 12694 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12682 14841 12694 14844
rect 12728 14872 12740 14875
rect 13262 14872 13268 14884
rect 12728 14844 13268 14872
rect 12728 14841 12740 14844
rect 12682 14835 12740 14841
rect 13262 14832 13268 14844
rect 13320 14832 13326 14884
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 6472 14776 8217 14804
rect 6181 14767 6239 14773
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 9548 14776 9593 14804
rect 9548 14764 9554 14776
rect 10134 14764 10140 14816
rect 10192 14804 10198 14816
rect 10229 14807 10287 14813
rect 10229 14804 10241 14807
rect 10192 14776 10241 14804
rect 10192 14764 10198 14776
rect 10229 14773 10241 14776
rect 10275 14804 10287 14807
rect 11146 14804 11152 14816
rect 10275 14776 11152 14804
rect 10275 14773 10287 14776
rect 10229 14767 10287 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 11882 14804 11888 14816
rect 11296 14776 11341 14804
rect 11843 14776 11888 14804
rect 11296 14764 11302 14776
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 3142 14600 3148 14612
rect 3103 14572 3148 14600
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 3418 14560 3424 14612
rect 3476 14600 3482 14612
rect 3513 14603 3571 14609
rect 3513 14600 3525 14603
rect 3476 14572 3525 14600
rect 3476 14560 3482 14572
rect 3513 14569 3525 14572
rect 3559 14569 3571 14603
rect 3513 14563 3571 14569
rect 3697 14603 3755 14609
rect 3697 14569 3709 14603
rect 3743 14600 3755 14603
rect 3786 14600 3792 14612
rect 3743 14572 3792 14600
rect 3743 14569 3755 14572
rect 3697 14563 3755 14569
rect 3712 14532 3740 14563
rect 3786 14560 3792 14572
rect 3844 14560 3850 14612
rect 3970 14560 3976 14612
rect 4028 14600 4034 14612
rect 4065 14603 4123 14609
rect 4065 14600 4077 14603
rect 4028 14572 4077 14600
rect 4028 14560 4034 14572
rect 4065 14569 4077 14572
rect 4111 14569 4123 14603
rect 4430 14600 4436 14612
rect 4391 14572 4436 14600
rect 4065 14563 4123 14569
rect 4430 14560 4436 14572
rect 4488 14560 4494 14612
rect 5718 14600 5724 14612
rect 5679 14572 5724 14600
rect 5718 14560 5724 14572
rect 5776 14560 5782 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 7098 14600 7104 14612
rect 6135 14572 7104 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 7098 14560 7104 14572
rect 7156 14600 7162 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7156 14572 7757 14600
rect 7156 14560 7162 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 7745 14563 7803 14569
rect 8021 14603 8079 14609
rect 8021 14569 8033 14603
rect 8067 14600 8079 14603
rect 9125 14603 9183 14609
rect 9125 14600 9137 14603
rect 8067 14572 9137 14600
rect 8067 14569 8079 14572
rect 8021 14563 8079 14569
rect 9125 14569 9137 14572
rect 9171 14600 9183 14603
rect 9490 14600 9496 14612
rect 9171 14572 9496 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 1504 14504 3740 14532
rect 6549 14535 6607 14541
rect 1504 14476 1532 14504
rect 6549 14501 6561 14535
rect 6595 14501 6607 14535
rect 7760 14532 7788 14563
rect 9490 14560 9496 14572
rect 9548 14560 9554 14612
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11422 14600 11428 14612
rect 11383 14572 11428 14600
rect 11422 14560 11428 14572
rect 11480 14560 11486 14612
rect 13262 14600 13268 14612
rect 13223 14572 13268 14600
rect 13262 14560 13268 14572
rect 13320 14560 13326 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 8938 14532 8944 14544
rect 7760 14504 8944 14532
rect 6549 14495 6607 14501
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1486 14464 1492 14476
rect 1443 14436 1492 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 1664 14467 1722 14473
rect 1664 14433 1676 14467
rect 1710 14464 1722 14467
rect 2866 14464 2872 14476
rect 1710 14436 2872 14464
rect 1710 14433 1722 14436
rect 1664 14427 1722 14433
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3878 14464 3884 14476
rect 3839 14436 3884 14464
rect 3878 14424 3884 14436
rect 3936 14424 3942 14476
rect 3970 14424 3976 14476
rect 4028 14464 4034 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 4028 14436 4537 14464
rect 4028 14424 4034 14436
rect 4525 14433 4537 14436
rect 4571 14464 4583 14467
rect 5905 14467 5963 14473
rect 4571 14436 4743 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4614 14396 4620 14408
rect 4575 14368 4620 14396
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 2498 14288 2504 14340
rect 2556 14328 2562 14340
rect 2777 14331 2835 14337
rect 2777 14328 2789 14331
rect 2556 14300 2789 14328
rect 2556 14288 2562 14300
rect 2777 14297 2789 14300
rect 2823 14328 2835 14331
rect 4632 14328 4660 14356
rect 2823 14300 4660 14328
rect 4715 14328 4743 14436
rect 5905 14433 5917 14467
rect 5951 14464 5963 14467
rect 6089 14467 6147 14473
rect 6089 14464 6101 14467
rect 5951 14436 6101 14464
rect 5951 14433 5963 14436
rect 5905 14427 5963 14433
rect 6089 14433 6101 14436
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6564 14464 6592 14495
rect 8938 14492 8944 14504
rect 8996 14492 9002 14544
rect 11072 14532 11100 14560
rect 11790 14532 11796 14544
rect 11072 14504 11796 14532
rect 11790 14492 11796 14504
rect 11848 14532 11854 14544
rect 12130 14535 12188 14541
rect 12130 14532 12142 14535
rect 11848 14504 12142 14532
rect 11848 14492 11854 14504
rect 12130 14501 12142 14504
rect 12176 14501 12188 14535
rect 12130 14495 12188 14501
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 13633 14535 13691 14541
rect 13633 14532 13645 14535
rect 13596 14504 13645 14532
rect 13596 14492 13602 14504
rect 13633 14501 13645 14504
rect 13679 14532 13691 14535
rect 14001 14535 14059 14541
rect 14001 14532 14013 14535
rect 13679 14504 14013 14532
rect 13679 14501 13691 14504
rect 13633 14495 13691 14501
rect 14001 14501 14013 14504
rect 14047 14532 14059 14535
rect 14182 14532 14188 14544
rect 14047 14504 14188 14532
rect 14047 14501 14059 14504
rect 14001 14495 14059 14501
rect 14182 14492 14188 14504
rect 14240 14492 14246 14544
rect 6512 14436 6592 14464
rect 7929 14467 7987 14473
rect 6512 14424 6518 14436
rect 7929 14433 7941 14467
rect 7975 14464 7987 14467
rect 8202 14464 8208 14476
rect 7975 14436 8208 14464
rect 7975 14433 7987 14436
rect 7929 14427 7987 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 8386 14464 8392 14476
rect 8347 14436 8392 14464
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 9933 14467 9991 14473
rect 9933 14464 9945 14467
rect 8588 14436 9945 14464
rect 8588 14408 8616 14436
rect 9933 14433 9945 14436
rect 9979 14433 9991 14467
rect 9933 14427 9991 14433
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14396 5687 14399
rect 5810 14396 5816 14408
rect 5675 14368 5816 14396
rect 5675 14365 5687 14368
rect 5629 14359 5687 14365
rect 5810 14356 5816 14368
rect 5868 14396 5874 14408
rect 6362 14396 6368 14408
rect 5868 14368 6368 14396
rect 5868 14356 5874 14368
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 6638 14396 6644 14408
rect 6599 14368 6644 14396
rect 6638 14356 6644 14368
rect 6696 14356 6702 14408
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 8478 14396 8484 14408
rect 6788 14368 6833 14396
rect 8439 14368 8484 14396
rect 6788 14356 6794 14368
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8570 14356 8576 14408
rect 8628 14396 8634 14408
rect 8628 14368 8673 14396
rect 8628 14356 8634 14368
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 9088 14368 9689 14396
rect 9088 14356 9094 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 11882 14396 11888 14408
rect 9677 14359 9735 14365
rect 10704 14368 11888 14396
rect 7561 14331 7619 14337
rect 7561 14328 7573 14331
rect 4715 14300 7573 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 7561 14297 7573 14300
rect 7607 14297 7619 14331
rect 7561 14291 7619 14297
rect 5258 14260 5264 14272
rect 5219 14232 5264 14260
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 6178 14260 6184 14272
rect 6139 14232 6184 14260
rect 6178 14220 6184 14232
rect 6236 14220 6242 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6730 14260 6736 14272
rect 6420 14232 6736 14260
rect 6420 14220 6426 14232
rect 6730 14220 6736 14232
rect 6788 14220 6794 14272
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 7374 14260 7380 14272
rect 7331 14232 7380 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 8444 14232 9413 14260
rect 8444 14220 8450 14232
rect 9401 14229 9413 14232
rect 9447 14229 9459 14263
rect 9692 14260 9720 14359
rect 10042 14260 10048 14272
rect 9692 14232 10048 14260
rect 9401 14223 9459 14229
rect 10042 14220 10048 14232
rect 10100 14260 10106 14272
rect 10704 14260 10732 14368
rect 11882 14356 11888 14368
rect 11940 14356 11946 14408
rect 11698 14260 11704 14272
rect 10100 14232 10732 14260
rect 11659 14232 11704 14260
rect 10100 14220 10106 14232
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 13538 14260 13544 14272
rect 11940 14232 13544 14260
rect 11940 14220 11946 14232
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 3694 14056 3700 14068
rect 3655 14028 3700 14056
rect 3694 14016 3700 14028
rect 3752 14016 3758 14068
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 4430 14056 4436 14068
rect 4387 14028 4436 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 4614 14056 4620 14068
rect 4575 14028 4620 14056
rect 4614 14016 4620 14028
rect 4672 14016 4678 14068
rect 5534 14016 5540 14068
rect 5592 14056 5598 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 5592 14028 6285 14056
rect 5592 14016 5598 14028
rect 6273 14025 6285 14028
rect 6319 14056 6331 14059
rect 6638 14056 6644 14068
rect 6319 14028 6644 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 7926 14016 7932 14068
rect 7984 14056 7990 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 7984 14028 8125 14056
rect 7984 14016 7990 14028
rect 8113 14025 8125 14028
rect 8159 14056 8171 14059
rect 8294 14056 8300 14068
rect 8159 14028 8300 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8757 14059 8815 14065
rect 8757 14025 8769 14059
rect 8803 14056 8815 14059
rect 9766 14056 9772 14068
rect 8803 14028 9772 14056
rect 8803 14025 8815 14028
rect 8757 14019 8815 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11238 14056 11244 14068
rect 11195 14028 11244 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11238 14016 11244 14028
rect 11296 14056 11302 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11296 14028 12449 14056
rect 11296 14016 11302 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 13538 14056 13544 14068
rect 13499 14028 13544 14056
rect 12437 14019 12495 14025
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 3329 13991 3387 13997
rect 3329 13988 3341 13991
rect 2924 13960 3341 13988
rect 2924 13948 2930 13960
rect 3329 13957 3341 13960
rect 3375 13988 3387 13991
rect 4798 13988 4804 14000
rect 3375 13960 4804 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 5316 13960 5764 13988
rect 5316 13948 5322 13960
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5736 13929 5764 13960
rect 6454 13948 6460 14000
rect 6512 13988 6518 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6512 13960 6561 13988
rect 6512 13948 6518 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6822 13988 6828 14000
rect 6783 13960 6828 13988
rect 6549 13951 6607 13957
rect 6822 13948 6828 13960
rect 6880 13948 6886 14000
rect 11790 13988 11796 14000
rect 11751 13960 11796 13988
rect 11790 13948 11796 13960
rect 11848 13948 11854 14000
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 5500 13892 5641 13920
rect 5500 13880 5506 13892
rect 5629 13889 5641 13892
rect 5675 13889 5687 13923
rect 5629 13883 5687 13889
rect 5721 13923 5779 13929
rect 5721 13889 5733 13923
rect 5767 13920 5779 13923
rect 6914 13920 6920 13932
rect 5767 13892 6920 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7374 13920 7380 13932
rect 7335 13892 7380 13920
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 9030 13920 9036 13932
rect 8991 13892 9036 13920
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12894 13920 12900 13932
rect 12299 13892 12900 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13081 13923 13139 13929
rect 13081 13889 13093 13923
rect 13127 13920 13139 13923
rect 13262 13920 13268 13932
rect 13127 13892 13268 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13920 14335 13923
rect 14366 13920 14372 13932
rect 14323 13892 14372 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 17862 13920 17868 13932
rect 16991 13892 17868 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 1578 13852 1584 13864
rect 1539 13824 1584 13852
rect 1578 13812 1584 13824
rect 1636 13812 1642 13864
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5123 13824 5580 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 1848 13787 1906 13793
rect 1848 13753 1860 13787
rect 1894 13784 1906 13787
rect 2498 13784 2504 13796
rect 1894 13756 2504 13784
rect 1894 13753 1906 13756
rect 1848 13747 1906 13753
rect 2498 13744 2504 13756
rect 2556 13744 2562 13796
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 2961 13719 3019 13725
rect 2961 13716 2973 13719
rect 2832 13688 2973 13716
rect 2832 13676 2838 13688
rect 2961 13685 2973 13688
rect 3007 13685 3019 13719
rect 3786 13716 3792 13728
rect 3747 13688 3792 13716
rect 2961 13679 3019 13685
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 5166 13716 5172 13728
rect 5127 13688 5172 13716
rect 5166 13676 5172 13688
rect 5224 13676 5230 13728
rect 5552 13725 5580 13824
rect 6178 13812 6184 13864
rect 6236 13852 6242 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6236 13824 7297 13852
rect 6236 13812 6242 13824
rect 7285 13821 7297 13824
rect 7331 13852 7343 13855
rect 8202 13852 8208 13864
rect 7331 13824 8208 13852
rect 7331 13821 7343 13824
rect 7285 13815 7343 13821
rect 8202 13812 8208 13824
rect 8260 13812 8266 13864
rect 8386 13852 8392 13864
rect 8312 13824 8392 13852
rect 5718 13744 5724 13796
rect 5776 13784 5782 13796
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 5776 13756 7205 13784
rect 5776 13744 5782 13756
rect 7193 13753 7205 13756
rect 7239 13784 7251 13787
rect 8312 13784 8340 13824
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8938 13852 8944 13864
rect 8899 13824 8944 13852
rect 8938 13812 8944 13824
rect 8996 13812 9002 13864
rect 13998 13852 14004 13864
rect 13959 13824 14004 13852
rect 13998 13812 14004 13824
rect 14056 13852 14062 13864
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14056 13824 14749 13852
rect 14056 13812 14062 13824
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 16666 13852 16672 13864
rect 16627 13824 16672 13852
rect 14737 13815 14795 13821
rect 16666 13812 16672 13824
rect 16724 13852 16730 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 16724 13824 17417 13852
rect 16724 13812 16730 13824
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 17405 13815 17463 13821
rect 7239 13756 8340 13784
rect 8665 13787 8723 13793
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 8665 13753 8677 13787
rect 8711 13784 8723 13787
rect 9300 13787 9358 13793
rect 9300 13784 9312 13787
rect 8711 13756 9312 13784
rect 8711 13753 8723 13756
rect 8665 13747 8723 13753
rect 9300 13753 9312 13756
rect 9346 13784 9358 13787
rect 9582 13784 9588 13796
rect 9346 13756 9588 13784
rect 9346 13753 9358 13756
rect 9300 13747 9358 13753
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 12584 13756 12817 13784
rect 12584 13744 12590 13756
rect 12805 13753 12817 13756
rect 12851 13753 12863 13787
rect 12805 13747 12863 13753
rect 5537 13719 5595 13725
rect 5537 13685 5549 13719
rect 5583 13716 5595 13719
rect 5994 13716 6000 13728
rect 5583 13688 6000 13716
rect 5583 13685 5595 13688
rect 5537 13679 5595 13685
rect 5994 13676 6000 13688
rect 6052 13676 6058 13728
rect 10042 13676 10048 13728
rect 10100 13716 10106 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 10100 13688 10425 13716
rect 10100 13676 10106 13688
rect 10413 13685 10425 13688
rect 10459 13716 10471 13719
rect 10689 13719 10747 13725
rect 10689 13716 10701 13719
rect 10459 13688 10701 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10689 13685 10701 13688
rect 10735 13685 10747 13719
rect 11238 13716 11244 13728
rect 11199 13688 11244 13716
rect 10689 13679 10747 13685
rect 11238 13676 11244 13688
rect 11296 13676 11302 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 2498 13512 2504 13524
rect 2459 13484 2504 13512
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 3881 13515 3939 13521
rect 2648 13484 3556 13512
rect 2648 13472 2654 13484
rect 2866 13444 2872 13456
rect 2792 13416 2872 13444
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2792 13308 2820 13416
rect 2866 13404 2872 13416
rect 2924 13404 2930 13456
rect 3528 13453 3556 13484
rect 3881 13481 3893 13515
rect 3927 13512 3939 13515
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 3927 13484 4537 13512
rect 3927 13481 3939 13484
rect 3881 13475 3939 13481
rect 4525 13481 4537 13484
rect 4571 13512 4583 13515
rect 5166 13512 5172 13524
rect 4571 13484 5172 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5258 13472 5264 13524
rect 5316 13512 5322 13524
rect 5534 13512 5540 13524
rect 5316 13484 5540 13512
rect 5316 13472 5322 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6178 13512 6184 13524
rect 6139 13484 6184 13512
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 6914 13512 6920 13524
rect 6875 13484 6920 13512
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8665 13515 8723 13521
rect 8665 13512 8677 13515
rect 8536 13484 8677 13512
rect 8536 13472 8542 13484
rect 8665 13481 8677 13484
rect 8711 13481 8723 13515
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 8665 13475 8723 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10045 13515 10103 13521
rect 10045 13512 10057 13515
rect 10008 13484 10057 13512
rect 10008 13472 10014 13484
rect 10045 13481 10057 13484
rect 10091 13512 10103 13515
rect 11238 13512 11244 13524
rect 10091 13484 11244 13512
rect 10091 13481 10103 13484
rect 10045 13475 10103 13481
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 11977 13515 12035 13521
rect 11977 13512 11989 13515
rect 11940 13484 11989 13512
rect 11940 13472 11946 13484
rect 11977 13481 11989 13484
rect 12023 13481 12035 13515
rect 12526 13512 12532 13524
rect 12487 13484 12532 13512
rect 11977 13475 12035 13481
rect 12526 13472 12532 13484
rect 12584 13472 12590 13524
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13262 13512 13268 13524
rect 12943 13484 13268 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13262 13472 13268 13484
rect 13320 13472 13326 13524
rect 3513 13447 3571 13453
rect 3513 13413 3525 13447
rect 3559 13444 3571 13447
rect 7282 13444 7288 13456
rect 3559 13416 7288 13444
rect 3559 13413 3571 13416
rect 3513 13407 3571 13413
rect 7282 13404 7288 13416
rect 7340 13404 7346 13456
rect 8294 13404 8300 13456
rect 8352 13444 8358 13456
rect 9401 13447 9459 13453
rect 9401 13444 9413 13447
rect 8352 13416 9413 13444
rect 8352 13404 8358 13416
rect 9401 13413 9413 13416
rect 9447 13413 9459 13447
rect 9401 13407 9459 13413
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 10137 13447 10195 13453
rect 10137 13444 10149 13447
rect 9916 13416 10149 13444
rect 9916 13404 9922 13416
rect 10137 13413 10149 13416
rect 10183 13413 10195 13447
rect 10137 13407 10195 13413
rect 17586 13404 17592 13456
rect 17644 13444 17650 13456
rect 17681 13447 17739 13453
rect 17681 13444 17693 13447
rect 17644 13416 17693 13444
rect 17644 13404 17650 13416
rect 17681 13413 17693 13416
rect 17727 13413 17739 13447
rect 17681 13407 17739 13413
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13376 6147 13379
rect 6546 13376 6552 13388
rect 6135 13348 6552 13376
rect 6135 13345 6147 13348
rect 6089 13339 6147 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 7653 13379 7711 13385
rect 7653 13345 7665 13379
rect 7699 13376 7711 13379
rect 8110 13376 8116 13388
rect 7699 13348 8116 13376
rect 7699 13345 7711 13348
rect 7653 13339 7711 13345
rect 8110 13336 8116 13348
rect 8168 13336 8174 13388
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8570 13376 8576 13388
rect 8435 13348 8576 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8570 13336 8576 13348
rect 8628 13376 8634 13388
rect 10042 13376 10048 13388
rect 8628 13348 10048 13376
rect 8628 13336 8634 13348
rect 10042 13336 10048 13348
rect 10100 13376 10106 13388
rect 17402 13376 17408 13388
rect 10100 13348 10272 13376
rect 17363 13348 17408 13376
rect 10100 13336 10106 13348
rect 1995 13280 2820 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2866 13268 2872 13320
rect 2924 13308 2930 13320
rect 2961 13311 3019 13317
rect 2961 13308 2973 13311
rect 2924 13280 2973 13308
rect 2924 13268 2930 13280
rect 2961 13277 2973 13280
rect 3007 13277 3019 13311
rect 2961 13271 3019 13277
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4120 13280 4629 13308
rect 4120 13268 4126 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4798 13308 4804 13320
rect 4759 13280 4804 13308
rect 4617 13271 4675 13277
rect 1397 13243 1455 13249
rect 1397 13209 1409 13243
rect 1443 13240 1455 13243
rect 3970 13240 3976 13252
rect 1443 13212 3976 13240
rect 1443 13209 1455 13212
rect 1397 13203 1455 13209
rect 3970 13200 3976 13212
rect 4028 13200 4034 13252
rect 4154 13240 4160 13252
rect 4115 13212 4160 13240
rect 4154 13200 4160 13212
rect 4212 13200 4218 13252
rect 4632 13240 4660 13271
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7742 13308 7748 13320
rect 7703 13280 7748 13308
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 10244 13317 10272 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 12434 13308 12440 13320
rect 11563 13280 12440 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 7285 13243 7343 13249
rect 7285 13240 7297 13243
rect 4632 13212 7297 13240
rect 7285 13209 7297 13212
rect 7331 13209 7343 13243
rect 7852 13240 7880 13271
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 7285 13203 7343 13209
rect 7760 13212 7880 13240
rect 9125 13243 9183 13249
rect 5534 13172 5540 13184
rect 5495 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7760 13172 7788 13212
rect 9125 13209 9137 13243
rect 9171 13240 9183 13243
rect 9582 13240 9588 13252
rect 9171 13212 9588 13240
rect 9171 13209 9183 13212
rect 9125 13203 9183 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 10686 13172 10692 13184
rect 6972 13144 7788 13172
rect 10647 13144 10692 13172
rect 6972 13132 6978 13144
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 11146 13172 11152 13184
rect 11107 13144 11152 13172
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1670 12968 1676 12980
rect 1627 12940 1676 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 1949 12971 2007 12977
rect 1949 12968 1961 12971
rect 1820 12940 1961 12968
rect 1820 12928 1826 12940
rect 1949 12937 1961 12940
rect 1995 12937 2007 12971
rect 1949 12931 2007 12937
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 4890 12968 4896 12980
rect 4755 12940 4896 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6546 12968 6552 12980
rect 6507 12940 6552 12968
rect 6546 12928 6552 12940
rect 6604 12928 6610 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 9033 12971 9091 12977
rect 9033 12968 9045 12971
rect 8536 12940 9045 12968
rect 8536 12928 8542 12940
rect 9033 12937 9045 12940
rect 9079 12937 9091 12971
rect 9033 12931 9091 12937
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10045 12971 10103 12977
rect 10045 12968 10057 12971
rect 9916 12940 10057 12968
rect 9916 12928 9922 12940
rect 10045 12937 10057 12940
rect 10091 12968 10103 12971
rect 10962 12968 10968 12980
rect 10091 12940 10968 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12968 11759 12971
rect 11882 12968 11888 12980
rect 11747 12940 11888 12968
rect 11747 12937 11759 12940
rect 11701 12931 11759 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 14550 12968 14556 12980
rect 14511 12940 14556 12968
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 17402 12968 17408 12980
rect 17363 12940 17408 12968
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 4154 12860 4160 12912
rect 4212 12900 4218 12912
rect 4801 12903 4859 12909
rect 4801 12900 4813 12903
rect 4212 12872 4813 12900
rect 4212 12860 4218 12872
rect 4801 12869 4813 12872
rect 4847 12900 4859 12903
rect 6270 12900 6276 12912
rect 4847 12872 5856 12900
rect 6231 12872 6276 12900
rect 4847 12869 4859 12872
rect 4801 12863 4859 12869
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 1636 12804 2513 12832
rect 1636 12792 1642 12804
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 5718 12832 5724 12844
rect 5679 12804 5724 12832
rect 2501 12795 2559 12801
rect 5718 12792 5724 12804
rect 5776 12792 5782 12844
rect 5828 12832 5856 12872
rect 6270 12860 6276 12872
rect 6328 12860 6334 12912
rect 8202 12900 8208 12912
rect 8163 12872 8208 12900
rect 8202 12860 8208 12872
rect 8260 12860 8266 12912
rect 13814 12900 13820 12912
rect 13775 12872 13820 12900
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 9582 12832 9588 12844
rect 5828 12804 6224 12832
rect 9543 12804 9588 12832
rect 6196 12776 6224 12804
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 11146 12832 11152 12844
rect 11107 12804 11152 12832
rect 11146 12792 11152 12804
rect 11204 12792 11210 12844
rect 14568 12832 14596 12928
rect 14568 12804 14780 12832
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 2590 12764 2596 12776
rect 1443 12736 2596 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 2774 12773 2780 12776
rect 2768 12727 2780 12773
rect 2832 12764 2838 12776
rect 4249 12767 4307 12773
rect 2832 12736 2868 12764
rect 2774 12724 2780 12727
rect 2832 12724 2838 12736
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4798 12764 4804 12776
rect 4295 12736 4804 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 4982 12764 4988 12776
rect 4943 12736 4988 12764
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5316 12736 5641 12764
rect 5316 12724 5322 12736
rect 5629 12733 5641 12736
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 6825 12767 6883 12773
rect 6825 12764 6837 12767
rect 6236 12736 6837 12764
rect 6236 12724 6242 12736
rect 6825 12733 6837 12736
rect 6871 12733 6883 12767
rect 6825 12727 6883 12733
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7081 12767 7139 12773
rect 7081 12764 7093 12767
rect 6972 12736 7093 12764
rect 6972 12724 6978 12736
rect 7081 12733 7093 12736
rect 7127 12733 7139 12767
rect 8846 12764 8852 12776
rect 8807 12736 8852 12764
rect 7081 12727 7139 12733
rect 8846 12724 8852 12736
rect 8904 12764 8910 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 8904 12736 9505 12764
rect 8904 12724 8910 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 10134 12724 10140 12776
rect 10192 12764 10198 12776
rect 10686 12764 10692 12776
rect 10192 12736 10692 12764
rect 10192 12724 10198 12736
rect 10686 12724 10692 12736
rect 10744 12764 10750 12776
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10744 12736 11069 12764
rect 10744 12724 10750 12736
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12526 12764 12532 12776
rect 12483 12736 12532 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 14642 12764 14648 12776
rect 14603 12736 14648 12764
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 14752 12764 14780 12804
rect 14901 12767 14959 12773
rect 14901 12764 14913 12767
rect 14752 12736 14913 12764
rect 14901 12733 14913 12736
rect 14947 12733 14959 12767
rect 14901 12727 14959 12733
rect 3142 12656 3148 12708
rect 3200 12696 3206 12708
rect 4890 12696 4896 12708
rect 3200 12668 4896 12696
rect 3200 12656 3206 12668
rect 4890 12656 4896 12668
rect 4948 12696 4954 12708
rect 5537 12699 5595 12705
rect 5537 12696 5549 12699
rect 4948 12668 5549 12696
rect 4948 12656 4954 12668
rect 5537 12665 5549 12668
rect 5583 12665 5595 12699
rect 5537 12659 5595 12665
rect 7742 12656 7748 12708
rect 7800 12696 7806 12708
rect 8481 12699 8539 12705
rect 8481 12696 8493 12699
rect 7800 12668 8493 12696
rect 7800 12656 7806 12668
rect 8481 12665 8493 12668
rect 8527 12665 8539 12699
rect 9398 12696 9404 12708
rect 9359 12668 9404 12696
rect 8481 12659 8539 12665
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 10505 12699 10563 12705
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 10778 12696 10784 12708
rect 10551 12668 10784 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 10778 12656 10784 12668
rect 10836 12696 10842 12708
rect 10965 12699 11023 12705
rect 10965 12696 10977 12699
rect 10836 12668 10977 12696
rect 10836 12656 10842 12668
rect 10965 12665 10977 12668
rect 11011 12665 11023 12699
rect 12250 12696 12256 12708
rect 12163 12668 12256 12696
rect 10965 12659 11023 12665
rect 12250 12656 12256 12668
rect 12308 12696 12314 12708
rect 12682 12699 12740 12705
rect 12682 12696 12694 12699
rect 12308 12668 12694 12696
rect 12308 12656 12314 12668
rect 12682 12665 12694 12668
rect 12728 12665 12740 12699
rect 12682 12659 12740 12665
rect 1854 12588 1860 12640
rect 1912 12628 1918 12640
rect 2409 12631 2467 12637
rect 2409 12628 2421 12631
rect 1912 12600 2421 12628
rect 1912 12588 1918 12600
rect 2409 12597 2421 12600
rect 2455 12628 2467 12631
rect 2682 12628 2688 12640
rect 2455 12600 2688 12628
rect 2455 12597 2467 12600
rect 2409 12591 2467 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3234 12588 3240 12640
rect 3292 12628 3298 12640
rect 3881 12631 3939 12637
rect 3881 12628 3893 12631
rect 3292 12600 3893 12628
rect 3292 12588 3298 12600
rect 3881 12597 3893 12600
rect 3927 12597 3939 12631
rect 3881 12591 3939 12597
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 10870 12628 10876 12640
rect 10643 12600 10876 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 12400 12600 16037 12628
rect 12400 12588 12406 12600
rect 16025 12597 16037 12600
rect 16071 12597 16083 12631
rect 16025 12591 16083 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4062 12424 4068 12436
rect 3927 12396 4068 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 5442 12424 5448 12436
rect 4571 12396 5448 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 5997 12427 6055 12433
rect 5997 12393 6009 12427
rect 6043 12424 6055 12427
rect 6362 12424 6368 12436
rect 6043 12396 6368 12424
rect 6043 12393 6055 12396
rect 5997 12387 6055 12393
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7469 12427 7527 12433
rect 7469 12424 7481 12427
rect 6972 12396 7481 12424
rect 6972 12384 6978 12396
rect 7469 12393 7481 12396
rect 7515 12424 7527 12427
rect 7745 12427 7803 12433
rect 7745 12424 7757 12427
rect 7515 12396 7757 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7745 12393 7757 12396
rect 7791 12393 7803 12427
rect 7745 12387 7803 12393
rect 8938 12384 8944 12436
rect 8996 12424 9002 12436
rect 9401 12427 9459 12433
rect 9401 12424 9413 12427
rect 8996 12396 9413 12424
rect 8996 12384 9002 12396
rect 9401 12393 9413 12396
rect 9447 12393 9459 12427
rect 9950 12424 9956 12436
rect 9911 12396 9956 12424
rect 9401 12387 9459 12393
rect 9950 12384 9956 12396
rect 10008 12384 10014 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10100 12396 10241 12424
rect 10100 12384 10106 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 12250 12424 12256 12436
rect 12163 12396 12256 12424
rect 10229 12387 10287 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 13078 12424 13084 12436
rect 12492 12396 13084 12424
rect 12492 12384 12498 12396
rect 13078 12384 13084 12396
rect 13136 12424 13142 12436
rect 13449 12427 13507 12433
rect 13449 12424 13461 12427
rect 13136 12396 13461 12424
rect 13136 12384 13142 12396
rect 13449 12393 13461 12396
rect 13495 12393 13507 12427
rect 14642 12424 14648 12436
rect 14603 12396 14648 12424
rect 13449 12387 13507 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 20990 12384 20996 12436
rect 21048 12384 21054 12436
rect 4985 12359 5043 12365
rect 4985 12325 4997 12359
rect 5031 12356 5043 12359
rect 6454 12356 6460 12368
rect 5031 12328 6460 12356
rect 5031 12325 5043 12328
rect 4985 12319 5043 12325
rect 6454 12316 6460 12328
rect 6512 12316 6518 12368
rect 8294 12356 8300 12368
rect 8255 12328 8300 12356
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 11146 12365 11152 12368
rect 11140 12356 11152 12365
rect 11107 12328 11152 12356
rect 11140 12319 11152 12328
rect 11146 12316 11152 12319
rect 11204 12316 11210 12368
rect 12268 12356 12296 12384
rect 13538 12356 13544 12368
rect 12268 12328 13216 12356
rect 13499 12328 13544 12356
rect 2032 12291 2090 12297
rect 2032 12257 2044 12291
rect 2078 12288 2090 12291
rect 2590 12288 2596 12300
rect 2078 12260 2596 12288
rect 2078 12257 2090 12260
rect 2032 12251 2090 12257
rect 2590 12248 2596 12260
rect 2648 12248 2654 12300
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4488 12260 4905 12288
rect 4488 12248 4494 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 5629 12291 5687 12297
rect 5629 12288 5641 12291
rect 4893 12251 4951 12257
rect 5184 12260 5641 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 5184 12229 5212 12260
rect 5629 12257 5641 12260
rect 5675 12288 5687 12291
rect 5718 12288 5724 12300
rect 5675 12260 5724 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 5718 12248 5724 12260
rect 5776 12288 5782 12300
rect 6356 12291 6414 12297
rect 6356 12288 6368 12291
rect 5776 12260 6368 12288
rect 5776 12248 5782 12260
rect 6356 12257 6368 12260
rect 6402 12288 6414 12291
rect 6638 12288 6644 12300
rect 6402 12260 6644 12288
rect 6402 12257 6414 12260
rect 6356 12251 6414 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 9766 12248 9772 12300
rect 9824 12288 9830 12300
rect 10597 12291 10655 12297
rect 10597 12288 10609 12291
rect 9824 12260 10609 12288
rect 9824 12248 9830 12260
rect 10597 12257 10609 12260
rect 10643 12288 10655 12291
rect 11882 12288 11888 12300
rect 10643 12260 11888 12288
rect 10643 12257 10655 12260
rect 10597 12251 10655 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 1765 12223 1823 12229
rect 1765 12220 1777 12223
rect 1452 12192 1777 12220
rect 1452 12180 1458 12192
rect 1765 12189 1777 12192
rect 1811 12189 1823 12223
rect 1765 12183 1823 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 4387 12192 5181 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 5169 12189 5181 12192
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5960 12192 6101 12220
rect 5960 12180 5966 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 12526 12220 12532 12232
rect 10873 12183 10931 12189
rect 12452 12192 12532 12220
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 3421 12155 3479 12161
rect 3421 12152 3433 12155
rect 2832 12124 3433 12152
rect 2832 12112 2838 12124
rect 3421 12121 3433 12124
rect 3467 12121 3479 12155
rect 8110 12152 8116 12164
rect 8071 12124 8116 12152
rect 3421 12115 3479 12121
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 1673 12087 1731 12093
rect 1673 12053 1685 12087
rect 1719 12084 1731 12087
rect 1762 12084 1768 12096
rect 1719 12056 1768 12084
rect 1719 12053 1731 12056
rect 1673 12047 1731 12053
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 2866 12084 2872 12096
rect 2740 12056 2872 12084
rect 2740 12044 2746 12056
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3145 12087 3203 12093
rect 3145 12053 3157 12087
rect 3191 12084 3203 12087
rect 3694 12084 3700 12096
rect 3191 12056 3700 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 3694 12044 3700 12056
rect 3752 12044 3758 12096
rect 9030 12084 9036 12096
rect 8991 12056 9036 12084
rect 9030 12044 9036 12056
rect 9088 12084 9094 12096
rect 9398 12084 9404 12096
rect 9088 12056 9404 12084
rect 9088 12044 9094 12056
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 9858 12044 9864 12096
rect 9916 12084 9922 12096
rect 10413 12087 10471 12093
rect 10413 12084 10425 12087
rect 9916 12056 10425 12084
rect 9916 12044 9922 12056
rect 10413 12053 10425 12056
rect 10459 12084 10471 12087
rect 10888 12084 10916 12183
rect 11238 12084 11244 12096
rect 10459 12056 11244 12084
rect 10459 12053 10471 12056
rect 10413 12047 10471 12053
rect 11238 12044 11244 12056
rect 11296 12084 11302 12096
rect 12452 12084 12480 12192
rect 12526 12180 12532 12192
rect 12584 12220 12590 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12584 12192 12633 12220
rect 12584 12180 12590 12192
rect 12621 12189 12633 12192
rect 12667 12220 12679 12223
rect 13188 12220 13216 12328
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 20806 12316 20812 12368
rect 20864 12356 20870 12368
rect 21008 12356 21036 12384
rect 21177 12359 21235 12365
rect 21177 12356 21189 12359
rect 20864 12328 20944 12356
rect 21008 12328 21189 12356
rect 20864 12316 20870 12328
rect 20916 12297 20944 12328
rect 21177 12325 21189 12328
rect 21223 12325 21235 12359
rect 21177 12319 21235 12325
rect 20901 12291 20959 12297
rect 20901 12257 20913 12291
rect 20947 12257 20959 12291
rect 20901 12251 20959 12257
rect 13446 12220 13452 12232
rect 12667 12192 13124 12220
rect 13188 12192 13452 12220
rect 12667 12189 12679 12192
rect 12621 12183 12679 12189
rect 13096 12152 13124 12192
rect 13446 12180 13452 12192
rect 13504 12220 13510 12232
rect 13633 12223 13691 12229
rect 13633 12220 13645 12223
rect 13504 12192 13645 12220
rect 13504 12180 13510 12192
rect 13633 12189 13645 12192
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 14642 12152 14648 12164
rect 13096 12124 14648 12152
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 11296 12056 12480 12084
rect 13081 12087 13139 12093
rect 11296 12044 11302 12056
rect 13081 12053 13093 12087
rect 13127 12084 13139 12087
rect 13722 12084 13728 12096
rect 13127 12056 13728 12084
rect 13127 12053 13139 12056
rect 13081 12047 13139 12053
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 4062 11880 4068 11892
rect 1452 11852 4068 11880
rect 1452 11840 1458 11852
rect 1670 11704 1676 11756
rect 1728 11744 1734 11756
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1728 11716 1961 11744
rect 1728 11704 1734 11716
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 2498 11744 2504 11756
rect 2459 11716 2504 11744
rect 1949 11707 2007 11713
rect 2498 11704 2504 11716
rect 2556 11704 2562 11756
rect 2976 11753 3004 11852
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 5166 11880 5172 11892
rect 5127 11852 5172 11880
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6454 11880 6460 11892
rect 6319 11852 6460 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6454 11840 6460 11852
rect 6512 11840 6518 11892
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 8113 11883 8171 11889
rect 8113 11880 8125 11883
rect 6788 11852 8125 11880
rect 6788 11840 6794 11852
rect 8113 11849 8125 11852
rect 8159 11880 8171 11883
rect 8159 11852 8984 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 4890 11772 4896 11824
rect 4948 11812 4954 11824
rect 4985 11815 5043 11821
rect 4985 11812 4997 11815
rect 4948 11784 4997 11812
rect 4948 11772 4954 11784
rect 4985 11781 4997 11784
rect 5031 11812 5043 11815
rect 5074 11812 5080 11824
rect 5031 11784 5080 11812
rect 5031 11781 5043 11784
rect 4985 11775 5043 11781
rect 5074 11772 5080 11784
rect 5132 11812 5138 11824
rect 6365 11815 6423 11821
rect 6365 11812 6377 11815
rect 5132 11784 5672 11812
rect 5132 11772 5138 11784
rect 5644 11753 5672 11784
rect 5828 11784 6377 11812
rect 5828 11753 5856 11784
rect 6365 11781 6377 11784
rect 6411 11781 6423 11815
rect 6472 11812 6500 11840
rect 7745 11815 7803 11821
rect 7745 11812 7757 11815
rect 6472 11784 7757 11812
rect 6365 11775 6423 11781
rect 7745 11781 7757 11784
rect 7791 11812 7803 11815
rect 7791 11784 8708 11812
rect 7791 11781 7803 11784
rect 7745 11775 7803 11781
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11713 5871 11747
rect 5813 11707 5871 11713
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6052 11716 6837 11744
rect 6052 11704 6058 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 8570 11744 8576 11756
rect 7515 11716 8576 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 8570 11704 8576 11716
rect 8628 11704 8634 11756
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11676 1915 11679
rect 2516 11676 2544 11704
rect 1903 11648 2544 11676
rect 1903 11645 1915 11648
rect 1857 11639 1915 11645
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 3050 11676 3056 11688
rect 2832 11648 3056 11676
rect 2832 11636 2838 11648
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 5258 11636 5264 11688
rect 5316 11676 5322 11688
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 5316 11648 5549 11676
rect 5316 11636 5322 11648
rect 5537 11645 5549 11648
rect 5583 11676 5595 11679
rect 6086 11676 6092 11688
rect 5583 11648 6092 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6365 11679 6423 11685
rect 6365 11645 6377 11679
rect 6411 11676 6423 11679
rect 6638 11676 6644 11688
rect 6411 11648 6644 11676
rect 6411 11645 6423 11648
rect 6365 11639 6423 11645
rect 6638 11636 6644 11648
rect 6696 11676 6702 11688
rect 8294 11676 8300 11688
rect 6696 11648 8300 11676
rect 6696 11636 6702 11648
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8680 11685 8708 11784
rect 8846 11744 8852 11756
rect 8807 11716 8852 11744
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8956 11676 8984 11852
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9272 11852 9321 11880
rect 9272 11840 9278 11852
rect 9309 11849 9321 11852
rect 9355 11849 9367 11883
rect 9309 11843 9367 11849
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11241 11883 11299 11889
rect 11241 11880 11253 11883
rect 11204 11852 11253 11880
rect 11204 11840 11210 11852
rect 11241 11849 11253 11852
rect 11287 11880 11299 11883
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11287 11852 11529 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11517 11843 11575 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 13078 11880 13084 11892
rect 13039 11852 13084 11880
rect 13078 11840 13084 11852
rect 13136 11840 13142 11892
rect 13446 11880 13452 11892
rect 13407 11852 13452 11880
rect 13446 11840 13452 11852
rect 13504 11840 13510 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13817 11883 13875 11889
rect 13817 11880 13829 11883
rect 13596 11852 13829 11880
rect 13596 11840 13602 11852
rect 13817 11849 13829 11852
rect 13863 11849 13875 11883
rect 13817 11843 13875 11849
rect 9858 11744 9864 11756
rect 9819 11716 9864 11744
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 18322 11744 18328 11756
rect 18283 11716 18328 11744
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 18046 11676 18052 11688
rect 8803 11648 8984 11676
rect 18007 11648 18052 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 18046 11636 18052 11648
rect 18104 11676 18110 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18104 11648 18797 11676
rect 18104 11636 18110 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 18785 11639 18843 11645
rect 3234 11617 3240 11620
rect 2869 11611 2927 11617
rect 2869 11577 2881 11611
rect 2915 11608 2927 11611
rect 3228 11608 3240 11617
rect 2915 11580 3240 11608
rect 2915 11577 2927 11580
rect 2869 11571 2927 11577
rect 3228 11571 3240 11580
rect 3292 11608 3298 11620
rect 3602 11608 3608 11620
rect 3292 11580 3608 11608
rect 3234 11568 3240 11571
rect 3292 11568 3298 11580
rect 3602 11568 3608 11580
rect 3660 11568 3666 11620
rect 9674 11608 9680 11620
rect 8312 11580 9680 11608
rect 1397 11543 1455 11549
rect 1397 11509 1409 11543
rect 1443 11540 1455 11543
rect 1578 11540 1584 11552
rect 1443 11512 1584 11540
rect 1443 11509 1455 11512
rect 1397 11503 1455 11509
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 3326 11540 3332 11552
rect 2648 11512 3332 11540
rect 2648 11500 2654 11512
rect 3326 11500 3332 11512
rect 3384 11540 3390 11552
rect 4341 11543 4399 11549
rect 4341 11540 4353 11543
rect 3384 11512 4353 11540
rect 3384 11500 3390 11512
rect 4341 11509 4353 11512
rect 4387 11509 4399 11543
rect 4341 11503 4399 11509
rect 4430 11500 4436 11552
rect 4488 11540 4494 11552
rect 8312 11549 8340 11580
rect 9674 11568 9680 11580
rect 9732 11568 9738 11620
rect 9769 11611 9827 11617
rect 9769 11577 9781 11611
rect 9815 11608 9827 11611
rect 10042 11608 10048 11620
rect 9815 11580 10048 11608
rect 9815 11577 9827 11580
rect 9769 11571 9827 11577
rect 10042 11568 10048 11580
rect 10100 11617 10106 11620
rect 10100 11611 10164 11617
rect 10100 11577 10118 11611
rect 10152 11577 10164 11611
rect 10100 11571 10164 11577
rect 10100 11568 10106 11571
rect 4617 11543 4675 11549
rect 4617 11540 4629 11543
rect 4488 11512 4629 11540
rect 4488 11500 4494 11512
rect 4617 11509 4629 11512
rect 4663 11509 4675 11543
rect 4617 11503 4675 11509
rect 8297 11543 8355 11549
rect 8297 11509 8309 11543
rect 8343 11509 8355 11543
rect 20898 11540 20904 11552
rect 20859 11512 20904 11540
rect 8297 11503 8355 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 1728 11308 2881 11336
rect 1728 11296 1734 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 4028 11308 4077 11336
rect 4028 11296 4034 11308
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 5258 11336 5264 11348
rect 5219 11308 5264 11336
rect 4065 11299 4123 11305
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5629 11339 5687 11345
rect 5629 11305 5641 11339
rect 5675 11336 5687 11339
rect 6638 11336 6644 11348
rect 5675 11308 6644 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6733 11339 6791 11345
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 6822 11336 6828 11348
rect 6779 11308 6828 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 11057 11339 11115 11345
rect 11057 11336 11069 11339
rect 10100 11308 11069 11336
rect 10100 11296 10106 11308
rect 11057 11305 11069 11308
rect 11103 11305 11115 11339
rect 11057 11299 11115 11305
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 11296 11308 11345 11336
rect 11296 11296 11302 11308
rect 11333 11305 11345 11308
rect 11379 11305 11391 11339
rect 11333 11299 11391 11305
rect 2590 11228 2596 11280
rect 2648 11268 2654 11280
rect 3053 11271 3111 11277
rect 3053 11268 3065 11271
rect 2648 11240 3065 11268
rect 2648 11228 2654 11240
rect 3053 11237 3065 11240
rect 3099 11237 3111 11271
rect 3053 11231 3111 11237
rect 8846 11228 8852 11280
rect 8904 11268 8910 11280
rect 9582 11268 9588 11280
rect 8904 11240 9588 11268
rect 8904 11228 8910 11240
rect 9582 11228 9588 11240
rect 9640 11268 9646 11280
rect 9922 11271 9980 11277
rect 9922 11268 9934 11271
rect 9640 11240 9934 11268
rect 9640 11228 9646 11240
rect 9922 11237 9934 11240
rect 9968 11237 9980 11271
rect 9922 11231 9980 11237
rect 19797 11271 19855 11277
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 21174 11268 21180 11280
rect 19843 11240 21180 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 21174 11228 21180 11240
rect 21232 11228 21238 11280
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 1664 11203 1722 11209
rect 1664 11169 1676 11203
rect 1710 11200 1722 11203
rect 3234 11200 3240 11212
rect 1710 11172 3240 11200
rect 1710 11169 1722 11172
rect 1664 11163 1722 11169
rect 3234 11160 3240 11172
rect 3292 11200 3298 11212
rect 3694 11200 3700 11212
rect 3292 11172 3700 11200
rect 3292 11160 3298 11172
rect 3694 11160 3700 11172
rect 3752 11160 3758 11212
rect 4154 11160 4160 11212
rect 4212 11200 4218 11212
rect 4433 11203 4491 11209
rect 4433 11200 4445 11203
rect 4212 11172 4445 11200
rect 4212 11160 4218 11172
rect 4433 11169 4445 11172
rect 4479 11169 4491 11203
rect 4433 11163 4491 11169
rect 5534 11160 5540 11212
rect 5592 11200 5598 11212
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5592 11172 6009 11200
rect 5592 11160 5598 11172
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 8202 11200 8208 11212
rect 8163 11172 8208 11200
rect 5997 11163 6055 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 9490 11200 9496 11212
rect 8987 11172 9496 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 9490 11160 9496 11172
rect 9548 11200 9554 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9548 11172 9689 11200
rect 9548 11160 9554 11172
rect 9677 11169 9689 11172
rect 9723 11200 9735 11203
rect 9766 11200 9772 11212
rect 9723 11172 9772 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 19518 11200 19524 11212
rect 19479 11172 19524 11200
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 4062 11092 4068 11144
rect 4120 11132 4126 11144
rect 4525 11135 4583 11141
rect 4525 11132 4537 11135
rect 4120 11104 4537 11132
rect 4120 11092 4126 11104
rect 4525 11101 4537 11104
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 2777 11067 2835 11073
rect 2777 11033 2789 11067
rect 2823 11064 2835 11067
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2823 11036 2881 11064
rect 2823 11033 2835 11036
rect 2777 11027 2835 11033
rect 2869 11033 2881 11036
rect 2915 11064 2927 11067
rect 3421 11067 3479 11073
rect 3421 11064 3433 11067
rect 2915 11036 3433 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 3421 11033 3433 11036
rect 3467 11033 3479 11067
rect 4632 11064 4660 11095
rect 3421 11027 3479 11033
rect 3896 11036 4660 11064
rect 3896 11008 3924 11036
rect 5994 11024 6000 11076
rect 6052 11064 6058 11076
rect 6104 11064 6132 11095
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6236 11104 6281 11132
rect 6236 11092 6242 11104
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 7156 11104 8309 11132
rect 7156 11092 7162 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8297 11095 8355 11101
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11101 8539 11135
rect 8481 11095 8539 11101
rect 6052 11036 6132 11064
rect 6052 11024 6058 11036
rect 6362 11024 6368 11076
rect 6420 11064 6426 11076
rect 7009 11067 7067 11073
rect 7009 11064 7021 11067
rect 6420 11036 7021 11064
rect 6420 11024 6426 11036
rect 7009 11033 7021 11036
rect 7055 11064 7067 11067
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 7055 11036 7389 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 7377 11033 7389 11036
rect 7423 11033 7435 11067
rect 7834 11064 7840 11076
rect 7795 11036 7840 11064
rect 7377 11027 7435 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8496 11008 8524 11095
rect 3878 10996 3884 11008
rect 3839 10968 3884 10996
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3881 10795 3939 10801
rect 3881 10761 3893 10795
rect 3927 10792 3939 10795
rect 4154 10792 4160 10804
rect 3927 10764 4160 10792
rect 3927 10761 3939 10764
rect 3881 10755 3939 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7208 10764 7941 10792
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1946 10656 1952 10668
rect 1636 10628 1952 10656
rect 1636 10616 1642 10628
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 7208 10665 7236 10764
rect 7929 10761 7941 10764
rect 7975 10792 7987 10795
rect 8202 10792 8208 10804
rect 7975 10764 8208 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9582 10792 9588 10804
rect 9543 10764 9588 10792
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10625 7251 10659
rect 9600 10656 9628 10752
rect 10042 10684 10048 10736
rect 10100 10724 10106 10736
rect 10413 10727 10471 10733
rect 10413 10724 10425 10727
rect 10100 10696 10425 10724
rect 10100 10684 10106 10696
rect 10413 10693 10425 10696
rect 10459 10693 10471 10727
rect 10413 10687 10471 10693
rect 10686 10656 10692 10668
rect 9600 10628 10692 10656
rect 7193 10619 7251 10625
rect 1762 10548 1768 10600
rect 1820 10588 1826 10600
rect 2148 10588 2176 10619
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10744 10628 10977 10656
rect 10744 10616 10750 10628
rect 10965 10625 10977 10628
rect 11011 10656 11023 10659
rect 11425 10659 11483 10665
rect 11425 10656 11437 10659
rect 11011 10628 11437 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11425 10625 11437 10628
rect 11471 10625 11483 10659
rect 11425 10619 11483 10625
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 19242 10656 19248 10668
rect 18647 10628 19248 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 19889 10659 19947 10665
rect 19889 10625 19901 10659
rect 19935 10656 19947 10659
rect 19978 10656 19984 10668
rect 19935 10628 19984 10656
rect 19935 10625 19947 10628
rect 19889 10619 19947 10625
rect 19978 10616 19984 10628
rect 20036 10616 20042 10668
rect 2774 10588 2780 10600
rect 1820 10560 2780 10588
rect 1820 10548 1826 10560
rect 2774 10548 2780 10560
rect 2832 10588 2838 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2832 10560 3249 10588
rect 2832 10548 2838 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3970 10588 3976 10600
rect 3931 10560 3976 10588
rect 3237 10551 3295 10557
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 8478 10597 8484 10600
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8472 10588 8484 10597
rect 8439 10560 8484 10588
rect 8205 10551 8263 10557
rect 8472 10551 8484 10560
rect 2501 10523 2559 10529
rect 2501 10520 2513 10523
rect 1872 10492 2513 10520
rect 1486 10452 1492 10464
rect 1447 10424 1492 10452
rect 1486 10412 1492 10424
rect 1544 10412 1550 10464
rect 1578 10412 1584 10464
rect 1636 10452 1642 10464
rect 1872 10461 1900 10492
rect 2501 10489 2513 10492
rect 2547 10489 2559 10523
rect 2501 10483 2559 10489
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 4218 10523 4276 10529
rect 4218 10520 4230 10523
rect 3936 10492 4230 10520
rect 3936 10480 3942 10492
rect 4218 10489 4230 10492
rect 4264 10489 4276 10523
rect 4218 10483 4276 10489
rect 5994 10480 6000 10532
rect 6052 10520 6058 10532
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 6052 10492 6377 10520
rect 6052 10480 6058 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 8220 10520 8248 10551
rect 8478 10548 8484 10551
rect 8536 10548 8542 10600
rect 9766 10548 9772 10600
rect 9824 10588 9830 10600
rect 10229 10591 10287 10597
rect 10229 10588 10241 10591
rect 9824 10560 10241 10588
rect 9824 10548 9830 10560
rect 10229 10557 10241 10560
rect 10275 10588 10287 10591
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10275 10560 10885 10588
rect 10275 10557 10287 10560
rect 10229 10551 10287 10557
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 18322 10588 18328 10600
rect 18283 10560 18328 10588
rect 10873 10551 10931 10557
rect 18322 10548 18328 10560
rect 18380 10588 18386 10600
rect 19061 10591 19119 10597
rect 19061 10588 19073 10591
rect 18380 10560 19073 10588
rect 18380 10548 18386 10560
rect 19061 10557 19073 10560
rect 19107 10557 19119 10591
rect 19061 10551 19119 10557
rect 19518 10548 19524 10600
rect 19576 10588 19582 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19576 10560 19625 10588
rect 19576 10548 19582 10560
rect 19613 10557 19625 10560
rect 19659 10588 19671 10591
rect 20349 10591 20407 10597
rect 20349 10588 20361 10591
rect 19659 10560 20361 10588
rect 19659 10557 19671 10560
rect 19613 10551 19671 10557
rect 20349 10557 20361 10560
rect 20395 10557 20407 10591
rect 20349 10551 20407 10557
rect 9490 10520 9496 10532
rect 8220 10492 9496 10520
rect 6365 10483 6423 10489
rect 9490 10480 9496 10492
rect 9548 10480 9554 10532
rect 10781 10523 10839 10529
rect 10781 10520 10793 10523
rect 9876 10492 10793 10520
rect 9876 10464 9904 10492
rect 10781 10489 10793 10492
rect 10827 10489 10839 10523
rect 10781 10483 10839 10489
rect 1857 10455 1915 10461
rect 1857 10452 1869 10455
rect 1636 10424 1869 10452
rect 1636 10412 1642 10424
rect 1857 10421 1869 10424
rect 1903 10421 1915 10455
rect 1857 10415 1915 10421
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3234 10452 3240 10464
rect 3007 10424 3240 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5629 10455 5687 10461
rect 5629 10452 5641 10455
rect 5592 10424 5641 10452
rect 5592 10412 5598 10424
rect 5629 10421 5641 10424
rect 5675 10421 5687 10455
rect 5629 10415 5687 10421
rect 6089 10455 6147 10461
rect 6089 10421 6101 10455
rect 6135 10452 6147 10455
rect 6178 10452 6184 10464
rect 6135 10424 6184 10452
rect 6135 10421 6147 10424
rect 6089 10415 6147 10421
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 9858 10452 9864 10464
rect 9819 10424 9864 10452
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2774 10248 2780 10260
rect 2735 10220 2780 10248
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 4062 10248 4068 10260
rect 3559 10220 4068 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 4525 10251 4583 10257
rect 4525 10248 4537 10251
rect 4304 10220 4537 10248
rect 4304 10208 4310 10220
rect 4525 10217 4537 10220
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 4982 10208 4988 10260
rect 5040 10248 5046 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 5040 10220 5089 10248
rect 5040 10208 5046 10220
rect 5077 10217 5089 10220
rect 5123 10248 5135 10251
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5123 10220 5457 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 7929 10251 7987 10257
rect 7929 10217 7941 10251
rect 7975 10248 7987 10251
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 7975 10220 8309 10248
rect 7975 10217 7987 10220
rect 7929 10211 7987 10217
rect 8297 10217 8309 10220
rect 8343 10248 8355 10251
rect 8478 10248 8484 10260
rect 8343 10220 8484 10248
rect 8343 10217 8355 10220
rect 8297 10211 8355 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 8573 10251 8631 10257
rect 8573 10217 8585 10251
rect 8619 10248 8631 10251
rect 9858 10248 9864 10260
rect 8619 10220 9864 10248
rect 8619 10217 8631 10220
rect 8573 10211 8631 10217
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10042 10248 10048 10260
rect 10003 10220 10048 10248
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 1946 10140 1952 10192
rect 2004 10180 2010 10192
rect 3053 10183 3111 10189
rect 3053 10180 3065 10183
rect 2004 10152 3065 10180
rect 2004 10140 2010 10152
rect 3053 10149 3065 10152
rect 3099 10149 3111 10183
rect 3053 10143 3111 10149
rect 3970 10140 3976 10192
rect 4028 10180 4034 10192
rect 4264 10180 4292 10208
rect 4028 10152 4292 10180
rect 4028 10140 4034 10152
rect 6178 10140 6184 10192
rect 6236 10189 6242 10192
rect 6236 10183 6300 10189
rect 6236 10149 6254 10183
rect 6288 10149 6300 10183
rect 9490 10180 9496 10192
rect 9451 10152 9496 10180
rect 6236 10143 6300 10149
rect 6236 10140 6242 10143
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 9950 10180 9956 10192
rect 9732 10152 9956 10180
rect 9732 10140 9738 10152
rect 9950 10140 9956 10152
rect 10008 10180 10014 10192
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 10008 10152 10149 10180
rect 10008 10140 10014 10152
rect 10137 10149 10149 10152
rect 10183 10149 10195 10183
rect 10137 10143 10195 10149
rect 1670 10121 1676 10124
rect 1664 10112 1676 10121
rect 1631 10084 1676 10112
rect 1664 10075 1676 10084
rect 1670 10072 1676 10075
rect 1728 10072 1734 10124
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4433 10115 4491 10121
rect 4433 10112 4445 10115
rect 3752 10084 4445 10112
rect 3752 10072 3758 10084
rect 4433 10081 4445 10084
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10044 4767 10047
rect 5074 10044 5080 10056
rect 4755 10016 5080 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5828 10016 6009 10044
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5828 9917 5856 10016
rect 5997 10013 6009 10016
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10134 10044 10140 10056
rect 9916 10016 10140 10044
rect 9916 10004 9922 10016
rect 10134 10004 10140 10016
rect 10192 10044 10198 10056
rect 10229 10047 10287 10053
rect 10229 10044 10241 10047
rect 10192 10016 10241 10044
rect 10192 10004 10198 10016
rect 10229 10013 10241 10016
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 9674 9976 9680 9988
rect 9635 9948 9680 9976
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 5813 9911 5871 9917
rect 5813 9908 5825 9911
rect 5224 9880 5825 9908
rect 5224 9868 5230 9880
rect 5813 9877 5825 9880
rect 5859 9908 5871 9911
rect 6362 9908 6368 9920
rect 5859 9880 6368 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 7374 9908 7380 9920
rect 7335 9880 7380 9908
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 1762 9704 1768 9716
rect 1723 9676 1768 9704
rect 1762 9664 1768 9676
rect 1820 9664 1826 9716
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 2556 9676 3188 9704
rect 2556 9664 2562 9676
rect 1780 9568 1808 9664
rect 3160 9568 3188 9676
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 3936 9676 5457 9704
rect 3936 9664 3942 9676
rect 5445 9673 5457 9676
rect 5491 9673 5503 9707
rect 5445 9667 5503 9673
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 6457 9707 6515 9713
rect 6457 9704 6469 9707
rect 6420 9676 6469 9704
rect 6420 9664 6426 9676
rect 6457 9673 6469 9676
rect 6503 9673 6515 9707
rect 8478 9704 8484 9716
rect 8439 9676 8484 9704
rect 6457 9667 6515 9673
rect 3605 9639 3663 9645
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 3970 9636 3976 9648
rect 3651 9608 3976 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 5132 9608 5733 9636
rect 5132 9596 5138 9608
rect 5721 9605 5733 9608
rect 5767 9605 5779 9639
rect 5721 9599 5779 9605
rect 1780 9540 1992 9568
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1854 9500 1860 9512
rect 1452 9472 1860 9500
rect 1452 9460 1458 9472
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 1964 9500 1992 9540
rect 2884 9540 3188 9568
rect 2113 9503 2171 9509
rect 2113 9500 2125 9503
rect 1964 9472 2125 9500
rect 2113 9469 2125 9472
rect 2159 9469 2171 9503
rect 2113 9463 2171 9469
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 2884 9500 2912 9540
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3292 9540 3464 9568
rect 3292 9528 3298 9540
rect 2740 9472 2912 9500
rect 2740 9460 2746 9472
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3326 9500 3332 9512
rect 3108 9472 3332 9500
rect 3108 9460 3114 9472
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 3436 9500 3464 9540
rect 3694 9528 3700 9580
rect 3752 9568 3758 9580
rect 3881 9571 3939 9577
rect 3881 9568 3893 9571
rect 3752 9540 3893 9568
rect 3752 9528 3758 9540
rect 3881 9537 3893 9540
rect 3927 9537 3939 9571
rect 3881 9531 3939 9537
rect 3970 9500 3976 9512
rect 3436 9472 3976 9500
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4338 9509 4344 9512
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9469 4123 9503
rect 4332 9500 4344 9509
rect 4251 9472 4344 9500
rect 4065 9463 4123 9469
rect 4332 9463 4344 9472
rect 4396 9500 4402 9512
rect 5092 9500 5120 9596
rect 6472 9568 6500 9667
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9858 9704 9864 9716
rect 9815 9676 9864 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10042 9664 10048 9716
rect 10100 9704 10106 9716
rect 10413 9707 10471 9713
rect 10413 9704 10425 9707
rect 10100 9676 10425 9704
rect 10100 9664 10106 9676
rect 10413 9673 10425 9676
rect 10459 9673 10471 9707
rect 10413 9667 10471 9673
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6472 9540 7113 9568
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 4396 9472 5120 9500
rect 7116 9500 7144 9531
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10045 9571 10103 9577
rect 10045 9568 10057 9571
rect 10008 9540 10057 9568
rect 10008 9528 10014 9540
rect 10045 9537 10057 9540
rect 10091 9537 10103 9571
rect 10045 9531 10103 9537
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 7116 9472 8769 9500
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 4080 9432 4108 9463
rect 4338 9460 4344 9463
rect 4396 9460 4402 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 7374 9441 7380 9444
rect 7368 9432 7380 9441
rect 2832 9404 4108 9432
rect 7335 9404 7380 9432
rect 2832 9392 2838 9404
rect 7368 9395 7380 9404
rect 7374 9392 7380 9395
rect 7432 9392 7438 9444
rect 3237 9367 3295 9373
rect 3237 9333 3249 9367
rect 3283 9364 3295 9367
rect 3326 9364 3332 9376
rect 3283 9336 3332 9364
rect 3283 9333 3295 9336
rect 3237 9327 3295 9333
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4430 9364 4436 9376
rect 3936 9336 4436 9364
rect 3936 9324 3942 9336
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 1949 9163 2007 9169
rect 1949 9160 1961 9163
rect 1912 9132 1961 9160
rect 1912 9120 1918 9132
rect 1949 9129 1961 9132
rect 1995 9129 2007 9163
rect 2590 9160 2596 9172
rect 2503 9132 2596 9160
rect 1949 9123 2007 9129
rect 1964 9024 1992 9123
rect 2590 9120 2596 9132
rect 2648 9160 2654 9172
rect 3142 9160 3148 9172
rect 2648 9132 3148 9160
rect 2648 9120 2654 9132
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3237 9163 3295 9169
rect 3237 9129 3249 9163
rect 3283 9160 3295 9163
rect 3786 9160 3792 9172
rect 3283 9132 3792 9160
rect 3283 9129 3295 9132
rect 3237 9123 3295 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 4062 9160 4068 9172
rect 4023 9132 4068 9160
rect 4062 9120 4068 9132
rect 4120 9120 4126 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 5258 9160 5264 9172
rect 4847 9132 5264 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 5258 9120 5264 9132
rect 5316 9120 5322 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6236 9132 6469 9160
rect 6236 9120 6242 9132
rect 6457 9129 6469 9132
rect 6503 9129 6515 9163
rect 6457 9123 6515 9129
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 7285 9163 7343 9169
rect 7285 9160 7297 9163
rect 7156 9132 7297 9160
rect 7156 9120 7162 9132
rect 7285 9129 7297 9132
rect 7331 9129 7343 9163
rect 7742 9160 7748 9172
rect 7703 9132 7748 9160
rect 7285 9123 7343 9129
rect 7742 9120 7748 9132
rect 7800 9120 7806 9172
rect 2314 9052 2320 9104
rect 2372 9092 2378 9104
rect 2501 9095 2559 9101
rect 2501 9092 2513 9095
rect 2372 9064 2513 9092
rect 2372 9052 2378 9064
rect 2501 9061 2513 9064
rect 2547 9061 2559 9095
rect 2501 9055 2559 9061
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3384 9064 3893 9092
rect 3384 9052 3390 9064
rect 3881 9061 3893 9064
rect 3927 9092 3939 9095
rect 4338 9092 4344 9104
rect 3927 9064 4344 9092
rect 3927 9061 3939 9064
rect 3881 9055 3939 9061
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 5350 9101 5356 9104
rect 5344 9092 5356 9101
rect 5311 9064 5356 9092
rect 5344 9055 5356 9064
rect 5350 9052 5356 9055
rect 5408 9052 5414 9104
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 6733 9095 6791 9101
rect 6733 9092 6745 9095
rect 6420 9064 6745 9092
rect 6420 9052 6426 9064
rect 6733 9061 6745 9064
rect 6779 9061 6791 9095
rect 7650 9092 7656 9104
rect 7611 9064 7656 9092
rect 6733 9055 6791 9061
rect 7650 9052 7656 9064
rect 7708 9052 7714 9104
rect 2774 9024 2780 9036
rect 1964 8996 2780 9024
rect 2774 8984 2780 8996
rect 2832 9024 2838 9036
rect 5074 9024 5080 9036
rect 2832 8996 5080 9024
rect 2832 8984 2838 8996
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2498 8956 2504 8968
rect 2280 8928 2504 8956
rect 2280 8916 2286 8928
rect 2498 8916 2504 8928
rect 2556 8956 2562 8968
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2556 8928 2697 8956
rect 2556 8916 2562 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8018 8956 8024 8968
rect 7975 8928 8024 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 7193 8891 7251 8897
rect 7193 8857 7205 8891
rect 7239 8888 7251 8891
rect 7374 8888 7380 8900
rect 7239 8860 7380 8888
rect 7239 8857 7251 8860
rect 7193 8851 7251 8857
rect 7374 8848 7380 8860
rect 7432 8888 7438 8900
rect 7944 8888 7972 8919
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 7432 8860 7972 8888
rect 7432 8848 7438 8860
rect 2133 8823 2191 8829
rect 2133 8789 2145 8823
rect 2179 8820 2191 8823
rect 2774 8820 2780 8832
rect 2179 8792 2780 8820
rect 2179 8789 2191 8792
rect 2133 8783 2191 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2314 8616 2320 8628
rect 2271 8588 2320 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3234 8616 3240 8628
rect 3007 8588 3240 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 4522 8616 4528 8628
rect 4483 8588 4528 8616
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 5994 8616 6000 8628
rect 4755 8588 6000 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 7742 8616 7748 8628
rect 7703 8588 7748 8616
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8018 8616 8024 8628
rect 7979 8588 8024 8616
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 7377 8551 7435 8557
rect 7377 8517 7389 8551
rect 7423 8548 7435 8551
rect 7650 8548 7656 8560
rect 7423 8520 7656 8548
rect 7423 8517 7435 8520
rect 7377 8511 7435 8517
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3234 8480 3240 8492
rect 2832 8452 3240 8480
rect 2832 8440 2838 8452
rect 3234 8440 3240 8452
rect 3292 8480 3298 8492
rect 3421 8483 3479 8489
rect 3421 8480 3433 8483
rect 3292 8452 3433 8480
rect 3292 8440 3298 8452
rect 3421 8449 3433 8452
rect 3467 8449 3479 8483
rect 3602 8480 3608 8492
rect 3563 8452 3608 8480
rect 3421 8443 3479 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 5350 8480 5356 8492
rect 4295 8452 5356 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 5350 8440 5356 8452
rect 5408 8480 5414 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5408 8452 5733 8480
rect 5408 8440 5414 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3694 8412 3700 8424
rect 3375 8384 3700 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 5077 8415 5135 8421
rect 5077 8412 5089 8415
rect 4580 8384 5089 8412
rect 4580 8372 4586 8384
rect 5077 8381 5089 8384
rect 5123 8381 5135 8415
rect 5077 8375 5135 8381
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8412 5227 8415
rect 5258 8412 5264 8424
rect 5215 8384 5264 8412
rect 5215 8381 5227 8384
rect 5169 8375 5227 8381
rect 5258 8372 5264 8384
rect 5316 8372 5322 8424
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1673 8075 1731 8081
rect 1673 8041 1685 8075
rect 1719 8072 1731 8075
rect 1854 8072 1860 8084
rect 1719 8044 1860 8072
rect 1719 8041 1731 8044
rect 1673 8035 1731 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2222 8072 2228 8084
rect 2183 8044 2228 8072
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 2958 8072 2964 8084
rect 2915 8044 2964 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3292 8044 3801 8072
rect 3292 8032 3298 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 3789 8035 3847 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4614 8072 4620 8084
rect 4571 8044 4620 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 5074 8072 5080 8084
rect 5035 8044 5080 8072
rect 5074 8032 5080 8044
rect 5132 8072 5138 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5132 8044 5457 8072
rect 5132 8032 5138 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5592 8044 5733 8072
rect 5592 8032 5598 8044
rect 5721 8041 5733 8044
rect 5767 8041 5779 8075
rect 5721 8035 5779 8041
rect 2682 7964 2688 8016
rect 2740 8004 2746 8016
rect 4154 8004 4160 8016
rect 2740 7976 4160 8004
rect 2740 7964 2746 7976
rect 4154 7964 4160 7976
rect 4212 8004 4218 8016
rect 4433 8007 4491 8013
rect 4433 8004 4445 8007
rect 4212 7976 4445 8004
rect 4212 7964 4218 7976
rect 4433 7973 4445 7976
rect 4479 7973 4491 8007
rect 4433 7967 4491 7973
rect 2777 7939 2835 7945
rect 2777 7905 2789 7939
rect 2823 7936 2835 7939
rect 2866 7936 2872 7948
rect 2823 7908 2872 7936
rect 2823 7905 2835 7908
rect 2777 7899 2835 7905
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 3513 7939 3571 7945
rect 3513 7905 3525 7939
rect 3559 7936 3571 7939
rect 3602 7936 3608 7948
rect 3559 7908 3608 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 3050 7868 3056 7880
rect 3011 7840 3056 7868
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4522 7868 4528 7880
rect 4028 7840 4528 7868
rect 4028 7828 4034 7840
rect 4522 7828 4528 7840
rect 4580 7868 4586 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 4580 7840 4629 7868
rect 4580 7828 4586 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 4062 7800 4068 7812
rect 4023 7772 4068 7800
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 4614 7732 4620 7744
rect 2455 7704 4620 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 1854 7528 1860 7540
rect 1719 7500 1860 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 1854 7488 1860 7500
rect 1912 7528 1918 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1912 7500 1961 7528
rect 1912 7488 1918 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2774 7528 2780 7540
rect 2547 7500 2780 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 2958 7528 2964 7540
rect 2915 7500 2964 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 3108 7500 3157 7528
rect 3108 7488 3114 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 3145 7491 3203 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 22373 7531 22431 7537
rect 4580 7500 4625 7528
rect 4580 7488 4586 7500
rect 22373 7497 22385 7531
rect 22419 7528 22431 7531
rect 23566 7528 23572 7540
rect 22419 7500 23572 7528
rect 22419 7497 22431 7500
rect 22373 7491 22431 7497
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 4614 7420 4620 7472
rect 4672 7460 4678 7472
rect 4801 7463 4859 7469
rect 4801 7460 4813 7463
rect 4672 7432 4813 7460
rect 4672 7420 4678 7432
rect 4801 7429 4813 7432
rect 4847 7429 4859 7463
rect 4801 7423 4859 7429
rect 22186 7324 22192 7336
rect 22099 7296 22192 7324
rect 22186 7284 22192 7296
rect 22244 7324 22250 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22244 7296 22753 7324
rect 22244 7284 22250 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 22741 7287 22799 7293
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 22738 6848 22744 6860
rect 22699 6820 22744 6848
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 22925 6715 22983 6721
rect 22925 6681 22937 6715
rect 22971 6712 22983 6715
rect 23382 6712 23388 6724
rect 22971 6684 23388 6712
rect 22971 6681 22983 6684
rect 22925 6675 22983 6681
rect 23382 6672 23388 6684
rect 23440 6672 23446 6724
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 22738 6440 22744 6452
rect 22699 6412 22744 6440
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 23845 6443 23903 6449
rect 23845 6409 23857 6443
rect 23891 6440 23903 6443
rect 25038 6440 25044 6452
rect 23891 6412 25044 6440
rect 23891 6409 23903 6412
rect 23845 6403 23903 6409
rect 25038 6400 25044 6412
rect 25096 6400 25102 6452
rect 23658 6236 23664 6248
rect 23619 6208 23664 6236
rect 23658 6196 23664 6208
rect 23716 6236 23722 6248
rect 24213 6239 24271 6245
rect 24213 6236 24225 6239
rect 23716 6208 24225 6236
rect 23716 6196 23722 6208
rect 24213 6205 24225 6208
rect 24259 6205 24271 6239
rect 24213 6199 24271 6205
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 24762 5896 24768 5908
rect 24167 5868 24768 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 23934 5760 23940 5772
rect 23895 5732 23940 5760
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 23934 5352 23940 5364
rect 23895 5324 23940 5352
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 24486 5148 24492 5160
rect 24447 5120 24492 5148
rect 24486 5108 24492 5120
rect 24544 5148 24550 5160
rect 25041 5151 25099 5157
rect 25041 5148 25053 5151
rect 24544 5120 25053 5148
rect 24544 5108 24550 5120
rect 25041 5117 25053 5120
rect 25087 5117 25099 5151
rect 25041 5111 25099 5117
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24762 4808 24768 4820
rect 24723 4780 24768 4808
rect 24762 4768 24768 4780
rect 24820 4768 24826 4820
rect 24578 4672 24584 4684
rect 24539 4644 24584 4672
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24670 4264 24676 4276
rect 24631 4236 24676 4264
rect 24670 4224 24676 4236
rect 24728 4224 24734 4276
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7466 4128 7472 4140
rect 7064 4100 7472 4128
rect 7064 4088 7070 4100
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 4068 26800 4120 26852
rect 7380 26800 7432 26852
rect 4068 26392 4120 26444
rect 12072 26392 12124 26444
rect 3516 26324 3568 26376
rect 11152 26324 11204 26376
rect 2044 25712 2096 25764
rect 8484 25712 8536 25764
rect 3516 25644 3568 25696
rect 13636 25644 13688 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 6184 25440 6236 25492
rect 6644 25440 6696 25492
rect 8208 25440 8260 25492
rect 4068 25372 4120 25424
rect 11152 25440 11204 25492
rect 13636 25483 13688 25492
rect 13636 25449 13645 25483
rect 13645 25449 13679 25483
rect 13679 25449 13688 25483
rect 13636 25440 13688 25449
rect 2320 25304 2372 25356
rect 2504 25347 2556 25356
rect 2504 25313 2513 25347
rect 2513 25313 2547 25347
rect 2547 25313 2556 25347
rect 2504 25304 2556 25313
rect 4896 25347 4948 25356
rect 4896 25313 4905 25347
rect 4905 25313 4939 25347
rect 4939 25313 4948 25347
rect 4896 25304 4948 25313
rect 4988 25347 5040 25356
rect 4988 25313 4997 25347
rect 4997 25313 5031 25347
rect 5031 25313 5040 25347
rect 4988 25304 5040 25313
rect 4160 25236 4212 25288
rect 6920 25304 6972 25356
rect 7656 25304 7708 25356
rect 8484 25347 8536 25356
rect 8484 25313 8493 25347
rect 8493 25313 8527 25347
rect 8527 25313 8536 25347
rect 8484 25304 8536 25313
rect 9680 25304 9732 25356
rect 10048 25304 10100 25356
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 12348 25236 12400 25288
rect 4712 25168 4764 25220
rect 5632 25168 5684 25220
rect 7288 25168 7340 25220
rect 7380 25168 7432 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 2780 25100 2832 25152
rect 3608 25100 3660 25152
rect 6000 25100 6052 25152
rect 10692 25100 10744 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 4988 24896 5040 24948
rect 9680 24939 9732 24948
rect 9680 24905 9689 24939
rect 9689 24905 9723 24939
rect 9723 24905 9732 24939
rect 9680 24896 9732 24905
rect 10876 24939 10928 24948
rect 10876 24905 10885 24939
rect 10885 24905 10919 24939
rect 10919 24905 10928 24939
rect 10876 24896 10928 24905
rect 4068 24828 4120 24880
rect 3608 24803 3660 24812
rect 3608 24769 3617 24803
rect 3617 24769 3651 24803
rect 3651 24769 3660 24803
rect 3608 24760 3660 24769
rect 4712 24760 4764 24812
rect 5080 24760 5132 24812
rect 5540 24760 5592 24812
rect 6644 24803 6696 24812
rect 6644 24769 6653 24803
rect 6653 24769 6687 24803
rect 6687 24769 6696 24803
rect 6644 24760 6696 24769
rect 7288 24803 7340 24812
rect 7288 24769 7297 24803
rect 7297 24769 7331 24803
rect 7331 24769 7340 24803
rect 7288 24760 7340 24769
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 3516 24735 3568 24744
rect 3516 24701 3525 24735
rect 3525 24701 3559 24735
rect 3559 24701 3568 24735
rect 3516 24692 3568 24701
rect 4620 24692 4672 24744
rect 6000 24692 6052 24744
rect 6920 24692 6972 24744
rect 2412 24624 2464 24676
rect 10140 24828 10192 24880
rect 12348 24760 12400 24812
rect 12624 24760 12676 24812
rect 12992 24803 13044 24812
rect 12992 24769 13001 24803
rect 13001 24769 13035 24803
rect 13035 24769 13044 24803
rect 12992 24760 13044 24769
rect 13360 24760 13412 24812
rect 13820 24760 13872 24812
rect 8668 24692 8720 24744
rect 1400 24556 1452 24608
rect 1860 24556 1912 24608
rect 2320 24599 2372 24608
rect 2320 24565 2329 24599
rect 2329 24565 2363 24599
rect 2363 24565 2372 24599
rect 2320 24556 2372 24565
rect 2688 24556 2740 24608
rect 8208 24624 8260 24676
rect 9588 24624 9640 24676
rect 10232 24667 10284 24676
rect 4160 24599 4212 24608
rect 4160 24565 4169 24599
rect 4169 24565 4203 24599
rect 4203 24565 4212 24599
rect 4160 24556 4212 24565
rect 4896 24599 4948 24608
rect 4896 24565 4905 24599
rect 4905 24565 4939 24599
rect 4939 24565 4948 24599
rect 4896 24556 4948 24565
rect 5172 24599 5224 24608
rect 5172 24565 5181 24599
rect 5181 24565 5215 24599
rect 5215 24565 5224 24599
rect 5172 24556 5224 24565
rect 6000 24556 6052 24608
rect 6828 24599 6880 24608
rect 6828 24565 6837 24599
rect 6837 24565 6871 24599
rect 6871 24565 6880 24599
rect 6828 24556 6880 24565
rect 6920 24556 6972 24608
rect 7564 24556 7616 24608
rect 8392 24556 8444 24608
rect 10232 24633 10241 24667
rect 10241 24633 10275 24667
rect 10275 24633 10284 24667
rect 10232 24624 10284 24633
rect 13084 24624 13136 24676
rect 14004 24667 14056 24676
rect 14004 24633 14013 24667
rect 14013 24633 14047 24667
rect 14047 24633 14056 24667
rect 14004 24624 14056 24633
rect 10692 24556 10744 24608
rect 12164 24556 12216 24608
rect 12624 24556 12676 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 3608 24352 3660 24404
rect 4620 24395 4672 24404
rect 4620 24361 4629 24395
rect 4629 24361 4663 24395
rect 4663 24361 4672 24395
rect 4620 24352 4672 24361
rect 8484 24352 8536 24404
rect 10692 24352 10744 24404
rect 12256 24352 12308 24404
rect 13084 24395 13136 24404
rect 13084 24361 13093 24395
rect 13093 24361 13127 24395
rect 13127 24361 13136 24395
rect 13084 24352 13136 24361
rect 16488 24352 16540 24404
rect 17868 24352 17920 24404
rect 18972 24395 19024 24404
rect 18972 24361 18981 24395
rect 18981 24361 19015 24395
rect 19015 24361 19024 24395
rect 18972 24352 19024 24361
rect 22468 24352 22520 24404
rect 5080 24284 5132 24336
rect 7472 24284 7524 24336
rect 9956 24284 10008 24336
rect 11704 24284 11756 24336
rect 12808 24284 12860 24336
rect 2596 24216 2648 24268
rect 2872 24216 2924 24268
rect 4068 24216 4120 24268
rect 1768 24191 1820 24200
rect 1768 24157 1777 24191
rect 1777 24157 1811 24191
rect 1811 24157 1820 24191
rect 1768 24148 1820 24157
rect 9312 24216 9364 24268
rect 11888 24259 11940 24268
rect 11888 24225 11897 24259
rect 11897 24225 11931 24259
rect 11931 24225 11940 24259
rect 11888 24216 11940 24225
rect 11980 24216 12032 24268
rect 16028 24216 16080 24268
rect 16120 24216 16172 24268
rect 17500 24259 17552 24268
rect 17500 24225 17509 24259
rect 17509 24225 17543 24259
rect 17543 24225 17552 24259
rect 17500 24216 17552 24225
rect 18788 24259 18840 24268
rect 18788 24225 18797 24259
rect 18797 24225 18831 24259
rect 18831 24225 18840 24259
rect 18788 24216 18840 24225
rect 21180 24216 21232 24268
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 10968 24148 11020 24200
rect 12348 24148 12400 24200
rect 14556 24148 14608 24200
rect 10048 24080 10100 24132
rect 12900 24080 12952 24132
rect 17684 24123 17736 24132
rect 17684 24089 17693 24123
rect 17693 24089 17727 24123
rect 17727 24089 17736 24123
rect 17684 24080 17736 24089
rect 1768 24012 1820 24064
rect 2504 24055 2556 24064
rect 2504 24021 2513 24055
rect 2513 24021 2547 24055
rect 2547 24021 2556 24055
rect 2504 24012 2556 24021
rect 2964 24055 3016 24064
rect 2964 24021 2973 24055
rect 2973 24021 3007 24055
rect 3007 24021 3016 24055
rect 2964 24012 3016 24021
rect 4160 24012 4212 24064
rect 6920 24055 6972 24064
rect 6920 24021 6929 24055
rect 6929 24021 6963 24055
rect 6963 24021 6972 24055
rect 6920 24012 6972 24021
rect 8392 24055 8444 24064
rect 8392 24021 8401 24055
rect 8401 24021 8435 24055
rect 8435 24021 8444 24055
rect 8392 24012 8444 24021
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 9864 24012 9916 24064
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 2872 23851 2924 23860
rect 2872 23817 2881 23851
rect 2881 23817 2915 23851
rect 2915 23817 2924 23851
rect 2872 23808 2924 23817
rect 5356 23851 5408 23860
rect 5356 23817 5365 23851
rect 5365 23817 5399 23851
rect 5399 23817 5408 23851
rect 5356 23808 5408 23817
rect 5540 23808 5592 23860
rect 7472 23808 7524 23860
rect 9956 23851 10008 23860
rect 9956 23817 9965 23851
rect 9965 23817 9999 23851
rect 9999 23817 10008 23851
rect 9956 23808 10008 23817
rect 12256 23808 12308 23860
rect 12808 23851 12860 23860
rect 12808 23817 12817 23851
rect 12817 23817 12851 23851
rect 12851 23817 12860 23851
rect 12808 23808 12860 23817
rect 14280 23851 14332 23860
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 16212 23808 16264 23860
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 19248 23808 19300 23860
rect 20260 23808 20312 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 23388 23808 23440 23860
rect 5080 23783 5132 23792
rect 5080 23749 5089 23783
rect 5089 23749 5123 23783
rect 5123 23749 5132 23783
rect 5080 23740 5132 23749
rect 8484 23783 8536 23792
rect 8484 23749 8493 23783
rect 8493 23749 8527 23783
rect 8527 23749 8536 23783
rect 8484 23740 8536 23749
rect 11980 23740 12032 23792
rect 4620 23672 4672 23724
rect 5264 23672 5316 23724
rect 2412 23604 2464 23656
rect 4068 23604 4120 23656
rect 5356 23604 5408 23656
rect 7012 23604 7064 23656
rect 10048 23647 10100 23656
rect 10048 23613 10057 23647
rect 10057 23613 10091 23647
rect 10091 23613 10100 23647
rect 10048 23604 10100 23613
rect 12348 23604 12400 23656
rect 12900 23647 12952 23656
rect 12900 23613 12909 23647
rect 12909 23613 12943 23647
rect 12943 23613 12952 23647
rect 12900 23604 12952 23613
rect 14372 23604 14424 23656
rect 1952 23579 2004 23588
rect 1952 23545 1961 23579
rect 1961 23545 1995 23579
rect 1995 23545 2004 23579
rect 1952 23536 2004 23545
rect 4160 23536 4212 23588
rect 8392 23536 8444 23588
rect 12992 23536 13044 23588
rect 13728 23536 13780 23588
rect 15568 23604 15620 23656
rect 18052 23647 18104 23656
rect 18052 23613 18061 23647
rect 18061 23613 18095 23647
rect 18095 23613 18104 23647
rect 18052 23604 18104 23613
rect 16580 23536 16632 23588
rect 17500 23579 17552 23588
rect 17500 23545 17509 23579
rect 17509 23545 17543 23579
rect 17543 23545 17552 23579
rect 17500 23536 17552 23545
rect 17592 23536 17644 23588
rect 19984 23604 20036 23656
rect 20996 23604 21048 23656
rect 22100 23604 22152 23656
rect 4712 23511 4764 23520
rect 4712 23477 4721 23511
rect 4721 23477 4755 23511
rect 4755 23477 4764 23511
rect 4712 23468 4764 23477
rect 9312 23468 9364 23520
rect 10876 23468 10928 23520
rect 14556 23511 14608 23520
rect 14556 23477 14565 23511
rect 14565 23477 14599 23511
rect 14599 23477 14608 23511
rect 14556 23468 14608 23477
rect 16028 23511 16080 23520
rect 16028 23477 16037 23511
rect 16037 23477 16071 23511
rect 16071 23477 16080 23511
rect 16028 23468 16080 23477
rect 16120 23468 16172 23520
rect 18328 23468 18380 23520
rect 18788 23468 18840 23520
rect 21180 23511 21232 23520
rect 21180 23477 21189 23511
rect 21189 23477 21223 23511
rect 21223 23477 21232 23511
rect 21180 23468 21232 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 2412 23307 2464 23316
rect 2412 23273 2421 23307
rect 2421 23273 2455 23307
rect 2455 23273 2464 23307
rect 2412 23264 2464 23273
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 8300 23264 8352 23316
rect 10968 23264 11020 23316
rect 11428 23264 11480 23316
rect 11888 23264 11940 23316
rect 12348 23264 12400 23316
rect 13728 23264 13780 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 16764 23264 16816 23273
rect 19524 23307 19576 23316
rect 19524 23273 19533 23307
rect 19533 23273 19567 23307
rect 19567 23273 19576 23307
rect 19524 23264 19576 23273
rect 2044 23196 2096 23248
rect 4712 23196 4764 23248
rect 2688 23128 2740 23180
rect 4068 23171 4120 23180
rect 2412 23060 2464 23112
rect 4068 23137 4077 23171
rect 4077 23137 4111 23171
rect 4111 23137 4120 23171
rect 4068 23128 4120 23137
rect 10140 23239 10192 23248
rect 10140 23205 10174 23239
rect 10174 23205 10192 23239
rect 10140 23196 10192 23205
rect 10876 23196 10928 23248
rect 15568 23239 15620 23248
rect 15568 23205 15577 23239
rect 15577 23205 15611 23239
rect 15611 23205 15620 23239
rect 15568 23196 15620 23205
rect 22008 23196 22060 23248
rect 7380 23171 7432 23180
rect 7380 23137 7414 23171
rect 7414 23137 7432 23171
rect 7380 23128 7432 23137
rect 9956 23128 10008 23180
rect 12348 23128 12400 23180
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 16580 23171 16632 23180
rect 16580 23137 16589 23171
rect 16589 23137 16623 23171
rect 16623 23137 16632 23171
rect 16580 23128 16632 23137
rect 19340 23171 19392 23180
rect 19340 23137 19349 23171
rect 19349 23137 19383 23171
rect 19383 23137 19392 23171
rect 19340 23128 19392 23137
rect 20904 23171 20956 23180
rect 20904 23137 20913 23171
rect 20913 23137 20947 23171
rect 20947 23137 20956 23171
rect 20904 23128 20956 23137
rect 2872 22924 2924 22976
rect 5448 22967 5500 22976
rect 5448 22933 5457 22967
rect 5457 22933 5491 22967
rect 5491 22933 5500 22967
rect 5448 22924 5500 22933
rect 6644 22924 6696 22976
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 12900 22924 12952 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 4712 22720 4764 22772
rect 6368 22763 6420 22772
rect 6368 22729 6377 22763
rect 6377 22729 6411 22763
rect 6411 22729 6420 22763
rect 6368 22720 6420 22729
rect 7012 22720 7064 22772
rect 7288 22763 7340 22772
rect 7288 22729 7297 22763
rect 7297 22729 7331 22763
rect 7331 22729 7340 22763
rect 7288 22720 7340 22729
rect 10140 22720 10192 22772
rect 2688 22652 2740 22704
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 3516 22584 3568 22636
rect 5264 22627 5316 22636
rect 2504 22516 2556 22568
rect 5264 22593 5273 22627
rect 5273 22593 5307 22627
rect 5307 22593 5316 22627
rect 5264 22584 5316 22593
rect 5448 22627 5500 22636
rect 5448 22593 5457 22627
rect 5457 22593 5491 22627
rect 5491 22593 5500 22627
rect 5448 22584 5500 22593
rect 7380 22584 7432 22636
rect 8116 22584 8168 22636
rect 9496 22584 9548 22636
rect 9956 22627 10008 22636
rect 9956 22593 9965 22627
rect 9965 22593 9999 22627
rect 9999 22593 10008 22627
rect 9956 22584 10008 22593
rect 4252 22516 4304 22568
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 6644 22516 6696 22568
rect 7748 22559 7800 22568
rect 7748 22525 7757 22559
rect 7757 22525 7791 22559
rect 7791 22525 7800 22559
rect 7748 22516 7800 22525
rect 9864 22559 9916 22568
rect 9864 22525 9873 22559
rect 9873 22525 9907 22559
rect 9907 22525 9916 22559
rect 9864 22516 9916 22525
rect 12164 22720 12216 22772
rect 12348 22652 12400 22704
rect 14556 22720 14608 22772
rect 15292 22720 15344 22772
rect 15752 22763 15804 22772
rect 15752 22729 15761 22763
rect 15761 22729 15795 22763
rect 15795 22729 15804 22763
rect 15752 22720 15804 22729
rect 12992 22584 13044 22636
rect 15384 22584 15436 22636
rect 3700 22448 3752 22500
rect 8300 22491 8352 22500
rect 8300 22457 8309 22491
rect 8309 22457 8343 22491
rect 8343 22457 8352 22491
rect 8300 22448 8352 22457
rect 11336 22491 11388 22500
rect 11336 22457 11345 22491
rect 11345 22457 11379 22491
rect 11379 22457 11388 22491
rect 11336 22448 11388 22457
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 13084 22380 13136 22432
rect 14740 22423 14792 22432
rect 14740 22389 14749 22423
rect 14749 22389 14783 22423
rect 14783 22389 14792 22423
rect 14740 22380 14792 22389
rect 16580 22423 16632 22432
rect 16580 22389 16589 22423
rect 16589 22389 16623 22423
rect 16623 22389 16632 22423
rect 16580 22380 16632 22389
rect 19340 22423 19392 22432
rect 19340 22389 19349 22423
rect 19349 22389 19383 22423
rect 19383 22389 19392 22423
rect 19340 22380 19392 22389
rect 20904 22423 20956 22432
rect 20904 22389 20913 22423
rect 20913 22389 20947 22423
rect 20947 22389 20956 22423
rect 20904 22380 20956 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2504 22176 2556 22228
rect 2688 22219 2740 22228
rect 2688 22185 2697 22219
rect 2697 22185 2731 22219
rect 2731 22185 2740 22219
rect 2688 22176 2740 22185
rect 3516 22219 3568 22228
rect 3516 22185 3525 22219
rect 3525 22185 3559 22219
rect 3559 22185 3568 22219
rect 3516 22176 3568 22185
rect 6368 22176 6420 22228
rect 16304 22219 16356 22228
rect 16304 22185 16313 22219
rect 16313 22185 16347 22219
rect 16347 22185 16356 22219
rect 16304 22176 16356 22185
rect 1584 22083 1636 22092
rect 1584 22049 1593 22083
rect 1593 22049 1627 22083
rect 1627 22049 1636 22083
rect 1584 22040 1636 22049
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 3700 22040 3752 22092
rect 4068 22108 4120 22160
rect 4344 22083 4396 22092
rect 4344 22049 4378 22083
rect 4378 22049 4396 22083
rect 4344 22040 4396 22049
rect 6460 22040 6512 22092
rect 8392 22040 8444 22092
rect 9588 22040 9640 22092
rect 10048 22108 10100 22160
rect 15292 22151 15344 22160
rect 15292 22117 15301 22151
rect 15301 22117 15335 22151
rect 15335 22117 15344 22151
rect 15292 22108 15344 22117
rect 10508 22040 10560 22092
rect 10968 22040 11020 22092
rect 11244 22040 11296 22092
rect 14648 22040 14700 22092
rect 4068 22015 4120 22024
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 8484 22015 8536 22024
rect 7012 21972 7064 21981
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 12992 22015 13044 22024
rect 3056 21947 3108 21956
rect 3056 21913 3065 21947
rect 3065 21913 3099 21947
rect 3099 21913 3108 21947
rect 3056 21904 3108 21913
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 4252 21836 4304 21888
rect 4436 21836 4488 21888
rect 5540 21836 5592 21888
rect 7656 21879 7708 21888
rect 7656 21845 7665 21879
rect 7665 21845 7699 21879
rect 7699 21845 7708 21879
rect 7656 21836 7708 21845
rect 8208 21836 8260 21888
rect 9404 21879 9456 21888
rect 9404 21845 9413 21879
rect 9413 21845 9447 21879
rect 9447 21845 9456 21879
rect 9404 21836 9456 21845
rect 9956 21836 10008 21888
rect 13176 21836 13228 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 2412 21675 2464 21684
rect 2412 21641 2421 21675
rect 2421 21641 2455 21675
rect 2455 21641 2464 21675
rect 2412 21632 2464 21641
rect 3700 21675 3752 21684
rect 3700 21641 3709 21675
rect 3709 21641 3743 21675
rect 3743 21641 3752 21675
rect 3700 21632 3752 21641
rect 4344 21632 4396 21684
rect 5448 21632 5500 21684
rect 1584 21564 1636 21616
rect 2688 21607 2740 21616
rect 2688 21573 2697 21607
rect 2697 21573 2731 21607
rect 2731 21573 2740 21607
rect 2688 21564 2740 21573
rect 2780 21564 2832 21616
rect 4160 21564 4212 21616
rect 6000 21632 6052 21684
rect 10508 21632 10560 21684
rect 13452 21632 13504 21684
rect 13820 21632 13872 21684
rect 2412 21428 2464 21480
rect 3516 21428 3568 21480
rect 4160 21471 4212 21480
rect 4160 21437 4191 21471
rect 4191 21437 4212 21471
rect 4160 21428 4212 21437
rect 8024 21539 8076 21548
rect 8024 21505 8033 21539
rect 8033 21505 8067 21539
rect 8067 21505 8076 21539
rect 8024 21496 8076 21505
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 10784 21496 10836 21548
rect 5724 21428 5776 21480
rect 7656 21428 7708 21480
rect 10968 21428 11020 21480
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 15384 21496 15436 21548
rect 13452 21428 13504 21480
rect 3976 21292 4028 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 6460 21335 6512 21344
rect 6460 21301 6469 21335
rect 6469 21301 6503 21335
rect 6503 21301 6512 21335
rect 6460 21292 6512 21301
rect 7012 21335 7064 21344
rect 7012 21301 7021 21335
rect 7021 21301 7055 21335
rect 7055 21301 7064 21335
rect 7012 21292 7064 21301
rect 7564 21335 7616 21344
rect 7564 21301 7573 21335
rect 7573 21301 7607 21335
rect 7607 21301 7616 21335
rect 7564 21292 7616 21301
rect 8852 21292 8904 21344
rect 9404 21292 9456 21344
rect 10048 21292 10100 21344
rect 11060 21292 11112 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 2964 21131 3016 21140
rect 2964 21097 2973 21131
rect 2973 21097 3007 21131
rect 3007 21097 3016 21131
rect 2964 21088 3016 21097
rect 3516 21131 3568 21140
rect 3516 21097 3525 21131
rect 3525 21097 3559 21131
rect 3559 21097 3568 21131
rect 3516 21088 3568 21097
rect 5724 21131 5776 21140
rect 5724 21097 5733 21131
rect 5733 21097 5767 21131
rect 5767 21097 5776 21131
rect 5724 21088 5776 21097
rect 6920 21088 6972 21140
rect 7564 21088 7616 21140
rect 8116 21131 8168 21140
rect 8116 21097 8125 21131
rect 8125 21097 8159 21131
rect 8159 21097 8168 21131
rect 8116 21088 8168 21097
rect 8392 21131 8444 21140
rect 8392 21097 8401 21131
rect 8401 21097 8435 21131
rect 8435 21097 8444 21131
rect 8392 21088 8444 21097
rect 9312 21131 9364 21140
rect 9312 21097 9321 21131
rect 9321 21097 9355 21131
rect 9355 21097 9364 21131
rect 9312 21088 9364 21097
rect 10784 21088 10836 21140
rect 12072 21131 12124 21140
rect 12072 21097 12081 21131
rect 12081 21097 12115 21131
rect 12115 21097 12124 21131
rect 12072 21088 12124 21097
rect 13084 21088 13136 21140
rect 14648 21088 14700 21140
rect 4436 21020 4488 21072
rect 9680 21020 9732 21072
rect 9956 21063 10008 21072
rect 9956 21029 9968 21063
rect 9968 21029 10008 21063
rect 9956 21020 10008 21029
rect 1952 20995 2004 21004
rect 1952 20961 1961 20995
rect 1961 20961 1995 20995
rect 1995 20961 2004 20995
rect 1952 20952 2004 20961
rect 4068 20995 4120 21004
rect 4068 20961 4077 20995
rect 4077 20961 4111 20995
rect 4111 20961 4120 20995
rect 4068 20952 4120 20961
rect 6368 20952 6420 21004
rect 6828 20952 6880 21004
rect 7012 20995 7064 21004
rect 7012 20961 7046 20995
rect 7046 20961 7064 20995
rect 7012 20952 7064 20961
rect 8576 20952 8628 21004
rect 11888 20995 11940 21004
rect 11888 20961 11897 20995
rect 11897 20961 11931 20995
rect 11931 20961 11940 20995
rect 11888 20952 11940 20961
rect 13084 20952 13136 21004
rect 12992 20927 13044 20936
rect 1952 20816 2004 20868
rect 2320 20748 2372 20800
rect 2780 20791 2832 20800
rect 2780 20757 2789 20791
rect 2789 20757 2823 20791
rect 2823 20757 2832 20791
rect 3884 20791 3936 20800
rect 2780 20748 2832 20757
rect 3884 20757 3893 20791
rect 3893 20757 3927 20791
rect 3927 20757 3936 20791
rect 3884 20748 3936 20757
rect 5448 20791 5500 20800
rect 5448 20757 5457 20791
rect 5457 20757 5491 20791
rect 5491 20757 5500 20791
rect 5448 20748 5500 20757
rect 6092 20791 6144 20800
rect 6092 20757 6101 20791
rect 6101 20757 6135 20791
rect 6135 20757 6144 20791
rect 6092 20748 6144 20757
rect 9588 20748 9640 20800
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 11152 20748 11204 20800
rect 14740 20791 14792 20800
rect 14740 20757 14749 20791
rect 14749 20757 14783 20791
rect 14783 20757 14792 20791
rect 14740 20748 14792 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 4436 20587 4488 20596
rect 4436 20553 4445 20587
rect 4445 20553 4479 20587
rect 4479 20553 4488 20587
rect 4436 20544 4488 20553
rect 7012 20544 7064 20596
rect 8576 20587 8628 20596
rect 8576 20553 8585 20587
rect 8585 20553 8619 20587
rect 8619 20553 8628 20587
rect 8576 20544 8628 20553
rect 9680 20544 9732 20596
rect 10416 20587 10468 20596
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 11152 20587 11204 20596
rect 11152 20553 11161 20587
rect 11161 20553 11195 20587
rect 11195 20553 11204 20587
rect 11152 20544 11204 20553
rect 11888 20587 11940 20596
rect 11888 20553 11897 20587
rect 11897 20553 11931 20587
rect 11931 20553 11940 20587
rect 11888 20544 11940 20553
rect 13084 20544 13136 20596
rect 14556 20544 14608 20596
rect 14740 20587 14792 20596
rect 14740 20553 14749 20587
rect 14749 20553 14783 20587
rect 14783 20553 14792 20587
rect 14740 20544 14792 20553
rect 2412 20519 2464 20528
rect 2412 20485 2421 20519
rect 2421 20485 2455 20519
rect 2455 20485 2464 20519
rect 2412 20476 2464 20485
rect 2136 20408 2188 20460
rect 2228 20408 2280 20460
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 5448 20408 5500 20460
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 5356 20340 5408 20392
rect 2780 20315 2832 20324
rect 2780 20281 2789 20315
rect 2789 20281 2823 20315
rect 2823 20281 2832 20315
rect 6920 20340 6972 20392
rect 8208 20340 8260 20392
rect 9588 20340 9640 20392
rect 13084 20383 13136 20392
rect 13084 20349 13093 20383
rect 13093 20349 13127 20383
rect 13127 20349 13136 20383
rect 13084 20340 13136 20349
rect 2780 20272 2832 20281
rect 9312 20315 9364 20324
rect 9312 20281 9346 20315
rect 9346 20281 9364 20315
rect 9312 20272 9364 20281
rect 10968 20272 11020 20324
rect 13452 20272 13504 20324
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 4068 20204 4120 20256
rect 4988 20247 5040 20256
rect 4988 20213 4997 20247
rect 4997 20213 5031 20247
rect 5031 20213 5040 20247
rect 4988 20204 5040 20213
rect 5080 20204 5132 20256
rect 9680 20204 9732 20256
rect 11336 20204 11388 20256
rect 15292 20247 15344 20256
rect 15292 20213 15301 20247
rect 15301 20213 15335 20247
rect 15335 20213 15344 20247
rect 15292 20204 15344 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 4988 20000 5040 20052
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 8208 20000 8260 20052
rect 8852 20000 8904 20052
rect 9312 20000 9364 20052
rect 11152 20000 11204 20052
rect 12348 20000 12400 20052
rect 13728 20000 13780 20052
rect 5264 19932 5316 19984
rect 5448 19975 5500 19984
rect 5448 19941 5482 19975
rect 5482 19941 5500 19975
rect 5448 19932 5500 19941
rect 8576 19932 8628 19984
rect 9956 19975 10008 19984
rect 9956 19941 9990 19975
rect 9990 19941 10008 19975
rect 9956 19932 10008 19941
rect 10784 19932 10836 19984
rect 11336 19975 11388 19984
rect 11336 19941 11345 19975
rect 11345 19941 11379 19975
rect 11379 19941 11388 19975
rect 11336 19932 11388 19941
rect 16028 19932 16080 19984
rect 2228 19864 2280 19916
rect 4160 19864 4212 19916
rect 7564 19907 7616 19916
rect 7564 19873 7573 19907
rect 7573 19873 7607 19907
rect 7607 19873 7616 19907
rect 7564 19864 7616 19873
rect 8392 19907 8444 19916
rect 8392 19873 8401 19907
rect 8401 19873 8435 19907
rect 8435 19873 8444 19907
rect 8392 19864 8444 19873
rect 13636 19864 13688 19916
rect 15200 19864 15252 19916
rect 15660 19864 15712 19916
rect 2412 19796 2464 19848
rect 3884 19839 3936 19848
rect 2504 19728 2556 19780
rect 3884 19805 3893 19839
rect 3893 19805 3927 19839
rect 3927 19805 3936 19839
rect 5172 19839 5224 19848
rect 3884 19796 3936 19805
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 9312 19796 9364 19848
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 3516 19728 3568 19780
rect 5080 19728 5132 19780
rect 1860 19660 1912 19712
rect 2228 19703 2280 19712
rect 2228 19669 2237 19703
rect 2237 19669 2271 19703
rect 2271 19669 2280 19703
rect 2228 19660 2280 19669
rect 3792 19660 3844 19712
rect 4068 19660 4120 19712
rect 5540 19660 5592 19712
rect 6644 19728 6696 19780
rect 14648 19771 14700 19780
rect 14648 19737 14657 19771
rect 14657 19737 14691 19771
rect 14691 19737 14700 19771
rect 14648 19728 14700 19737
rect 6552 19703 6604 19712
rect 6552 19669 6561 19703
rect 6561 19669 6595 19703
rect 6595 19669 6604 19703
rect 6552 19660 6604 19669
rect 7288 19703 7340 19712
rect 7288 19669 7297 19703
rect 7297 19669 7331 19703
rect 7331 19669 7340 19703
rect 7288 19660 7340 19669
rect 7932 19703 7984 19712
rect 7932 19669 7941 19703
rect 7941 19669 7975 19703
rect 7975 19669 7984 19703
rect 7932 19660 7984 19669
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 11336 19660 11388 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 12440 19660 12492 19669
rect 13084 19660 13136 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 5264 19456 5316 19508
rect 8576 19456 8628 19508
rect 9312 19456 9364 19508
rect 13452 19456 13504 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 15660 19499 15712 19508
rect 15660 19465 15669 19499
rect 15669 19465 15703 19499
rect 15703 19465 15712 19499
rect 15660 19456 15712 19465
rect 6552 19388 6604 19440
rect 7932 19388 7984 19440
rect 4988 19320 5040 19372
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 7288 19363 7340 19372
rect 5264 19320 5316 19329
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 8392 19320 8444 19372
rect 14556 19388 14608 19440
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 9220 19252 9272 19304
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 9772 19252 9824 19304
rect 11152 19252 11204 19304
rect 14648 19320 14700 19372
rect 25044 19320 25096 19372
rect 25320 19320 25372 19372
rect 12348 19252 12400 19304
rect 12440 19295 12492 19304
rect 12440 19261 12449 19295
rect 12449 19261 12483 19295
rect 12483 19261 12492 19295
rect 14464 19295 14516 19304
rect 12440 19252 12492 19261
rect 2504 19184 2556 19236
rect 4988 19227 5040 19236
rect 4988 19193 4997 19227
rect 4997 19193 5031 19227
rect 5031 19193 5040 19227
rect 4988 19184 5040 19193
rect 6920 19184 6972 19236
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 14464 19252 14516 19261
rect 10232 19184 10284 19236
rect 2136 19159 2188 19168
rect 2136 19125 2145 19159
rect 2145 19125 2179 19159
rect 2179 19125 2188 19159
rect 2136 19116 2188 19125
rect 3056 19116 3108 19168
rect 3976 19116 4028 19168
rect 4620 19159 4672 19168
rect 4620 19125 4629 19159
rect 4629 19125 4663 19159
rect 4663 19125 4672 19159
rect 4620 19116 4672 19125
rect 6460 19116 6512 19168
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 9496 19159 9548 19168
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 10048 19116 10100 19168
rect 10692 19184 10744 19236
rect 12532 19184 12584 19236
rect 12900 19184 12952 19236
rect 10968 19159 11020 19168
rect 10968 19125 10977 19159
rect 10977 19125 11011 19159
rect 11011 19125 11020 19159
rect 10968 19116 11020 19125
rect 11336 19116 11388 19168
rect 13636 19116 13688 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2412 18955 2464 18964
rect 2412 18921 2421 18955
rect 2421 18921 2455 18955
rect 2455 18921 2464 18955
rect 2412 18912 2464 18921
rect 4988 18912 5040 18964
rect 6460 18912 6512 18964
rect 7196 18912 7248 18964
rect 7564 18955 7616 18964
rect 7564 18921 7573 18955
rect 7573 18921 7607 18955
rect 7607 18921 7616 18955
rect 7564 18912 7616 18921
rect 8208 18912 8260 18964
rect 9588 18912 9640 18964
rect 12532 18955 12584 18964
rect 12532 18921 12541 18955
rect 12541 18921 12575 18955
rect 12575 18921 12584 18955
rect 12532 18912 12584 18921
rect 12808 18912 12860 18964
rect 13268 18912 13320 18964
rect 13820 18955 13872 18964
rect 13820 18921 13829 18955
rect 13829 18921 13863 18955
rect 13863 18921 13872 18955
rect 13820 18912 13872 18921
rect 14556 18912 14608 18964
rect 2964 18844 3016 18896
rect 6000 18844 6052 18896
rect 9956 18887 10008 18896
rect 9956 18853 9965 18887
rect 9965 18853 9999 18887
rect 9999 18853 10008 18887
rect 9956 18844 10008 18853
rect 10140 18844 10192 18896
rect 2872 18819 2924 18828
rect 2872 18785 2881 18819
rect 2881 18785 2915 18819
rect 2915 18785 2924 18819
rect 2872 18776 2924 18785
rect 3884 18776 3936 18828
rect 5448 18819 5500 18828
rect 5448 18785 5457 18819
rect 5457 18785 5491 18819
rect 5491 18785 5500 18819
rect 5448 18776 5500 18785
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 2780 18708 2832 18760
rect 5172 18640 5224 18692
rect 6092 18776 6144 18828
rect 7932 18776 7984 18828
rect 9036 18776 9088 18828
rect 10048 18776 10100 18828
rect 11336 18844 11388 18896
rect 12348 18844 12400 18896
rect 13360 18844 13412 18896
rect 11152 18776 11204 18828
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9680 18708 9732 18760
rect 10416 18708 10468 18760
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 1676 18572 1728 18624
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 4252 18572 4304 18581
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 7380 18572 7432 18624
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 2872 18368 2924 18420
rect 3056 18368 3108 18420
rect 7288 18368 7340 18420
rect 7932 18411 7984 18420
rect 7932 18377 7941 18411
rect 7941 18377 7975 18411
rect 7975 18377 7984 18411
rect 7932 18368 7984 18377
rect 8392 18411 8444 18420
rect 8392 18377 8401 18411
rect 8401 18377 8435 18411
rect 8435 18377 8444 18411
rect 8392 18368 8444 18377
rect 9496 18368 9548 18420
rect 9772 18300 9824 18352
rect 11060 18300 11112 18352
rect 6000 18232 6052 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 8300 18232 8352 18284
rect 11152 18232 11204 18284
rect 12348 18300 12400 18352
rect 12532 18300 12584 18352
rect 12808 18343 12860 18352
rect 12808 18309 12817 18343
rect 12817 18309 12851 18343
rect 12851 18309 12860 18343
rect 12808 18300 12860 18309
rect 2320 18164 2372 18216
rect 5172 18164 5224 18216
rect 8760 18207 8812 18216
rect 8760 18173 8769 18207
rect 8769 18173 8803 18207
rect 8803 18173 8812 18207
rect 8760 18164 8812 18173
rect 10140 18164 10192 18216
rect 11520 18164 11572 18216
rect 12716 18164 12768 18216
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 13728 18164 13780 18216
rect 1952 18139 2004 18148
rect 1952 18105 1986 18139
rect 1986 18105 2004 18139
rect 1952 18096 2004 18105
rect 2964 18096 3016 18148
rect 3976 18096 4028 18148
rect 4620 18096 4672 18148
rect 6368 18096 6420 18148
rect 8668 18096 8720 18148
rect 10416 18096 10468 18148
rect 13268 18096 13320 18148
rect 2136 18028 2188 18080
rect 2320 18028 2372 18080
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 8300 18071 8352 18080
rect 8300 18037 8309 18071
rect 8309 18037 8343 18071
rect 8343 18037 8352 18071
rect 8300 18028 8352 18037
rect 8576 18028 8628 18080
rect 10048 18028 10100 18080
rect 11060 18028 11112 18080
rect 11428 18028 11480 18080
rect 14556 18071 14608 18080
rect 14556 18037 14565 18071
rect 14565 18037 14599 18071
rect 14599 18037 14608 18071
rect 14556 18028 14608 18037
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2228 17824 2280 17876
rect 2688 17824 2740 17876
rect 3148 17824 3200 17876
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 6276 17824 6328 17876
rect 11152 17867 11204 17876
rect 11152 17833 11161 17867
rect 11161 17833 11195 17867
rect 11195 17833 11204 17867
rect 11152 17824 11204 17833
rect 11520 17867 11572 17876
rect 11520 17833 11529 17867
rect 11529 17833 11563 17867
rect 11563 17833 11572 17867
rect 11520 17824 11572 17833
rect 13268 17867 13320 17876
rect 13268 17833 13277 17867
rect 13277 17833 13311 17867
rect 13311 17833 13320 17867
rect 13268 17824 13320 17833
rect 13728 17867 13780 17876
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 14556 17824 14608 17876
rect 1768 17756 1820 17808
rect 3608 17756 3660 17808
rect 5540 17756 5592 17808
rect 6920 17756 6972 17808
rect 2688 17688 2740 17740
rect 4068 17731 4120 17740
rect 4068 17697 4077 17731
rect 4077 17697 4111 17731
rect 4111 17697 4120 17731
rect 4068 17688 4120 17697
rect 4988 17688 5040 17740
rect 6092 17688 6144 17740
rect 3884 17663 3936 17672
rect 1952 17595 2004 17604
rect 1952 17561 1961 17595
rect 1961 17561 1995 17595
rect 1995 17561 2004 17595
rect 1952 17552 2004 17561
rect 2780 17552 2832 17604
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 6000 17663 6052 17672
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 7656 17688 7708 17740
rect 9956 17688 10008 17740
rect 13084 17688 13136 17740
rect 14648 17688 14700 17740
rect 9772 17620 9824 17672
rect 11428 17620 11480 17672
rect 14004 17663 14056 17672
rect 4068 17552 4120 17604
rect 9680 17552 9732 17604
rect 3332 17484 3384 17536
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 6828 17527 6880 17536
rect 6828 17493 6837 17527
rect 6837 17493 6871 17527
rect 6871 17493 6880 17527
rect 6828 17484 6880 17493
rect 7840 17484 7892 17536
rect 8300 17527 8352 17536
rect 8300 17493 8309 17527
rect 8309 17493 8343 17527
rect 8343 17493 8352 17527
rect 8300 17484 8352 17493
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 9128 17484 9180 17536
rect 10140 17484 10192 17536
rect 14004 17629 14013 17663
rect 14013 17629 14047 17663
rect 14047 17629 14056 17663
rect 14004 17620 14056 17629
rect 12900 17484 12952 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 3148 17280 3200 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 6644 17280 6696 17332
rect 8208 17280 8260 17332
rect 9220 17280 9272 17332
rect 11428 17323 11480 17332
rect 11428 17289 11437 17323
rect 11437 17289 11471 17323
rect 11471 17289 11480 17323
rect 11428 17280 11480 17289
rect 13084 17323 13136 17332
rect 13084 17289 13093 17323
rect 13093 17289 13127 17323
rect 13127 17289 13136 17323
rect 13084 17280 13136 17289
rect 6828 17212 6880 17264
rect 7012 17212 7064 17264
rect 9128 17212 9180 17264
rect 23480 17212 23532 17264
rect 24768 17212 24820 17264
rect 24860 17212 24912 17264
rect 25964 17212 26016 17264
rect 5632 17144 5684 17196
rect 6000 17144 6052 17196
rect 10048 17187 10100 17196
rect 10048 17153 10057 17187
rect 10057 17153 10091 17187
rect 10091 17153 10100 17187
rect 10048 17144 10100 17153
rect 1584 17076 1636 17128
rect 2596 17076 2648 17128
rect 4988 17119 5040 17128
rect 1492 17008 1544 17060
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 5540 17119 5592 17128
rect 5540 17085 5549 17119
rect 5549 17085 5583 17119
rect 5583 17085 5592 17119
rect 5540 17076 5592 17085
rect 6092 17076 6144 17128
rect 10140 17076 10192 17128
rect 14556 17076 14608 17128
rect 3148 17008 3200 17060
rect 5080 17008 5132 17060
rect 2688 16940 2740 16992
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 5172 16983 5224 16992
rect 5172 16949 5181 16983
rect 5181 16949 5215 16983
rect 5215 16949 5224 16983
rect 5172 16940 5224 16949
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 6920 16940 6972 16992
rect 7472 16940 7524 16992
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 13728 16940 13780 16992
rect 14924 16983 14976 16992
rect 14924 16949 14933 16983
rect 14933 16949 14967 16983
rect 14967 16949 14976 16983
rect 14924 16940 14976 16949
rect 15200 16983 15252 16992
rect 15200 16949 15209 16983
rect 15209 16949 15243 16983
rect 15243 16949 15252 16983
rect 15200 16940 15252 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 1400 16736 1452 16788
rect 2412 16736 2464 16788
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 3240 16736 3292 16788
rect 3884 16736 3936 16788
rect 4068 16779 4120 16788
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 4068 16736 4120 16745
rect 4436 16779 4488 16788
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 5172 16736 5224 16788
rect 6552 16736 6604 16788
rect 9772 16736 9824 16788
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 11980 16779 12032 16788
rect 2688 16668 2740 16720
rect 4252 16668 4304 16720
rect 4804 16668 4856 16720
rect 5080 16668 5132 16720
rect 5356 16668 5408 16720
rect 1768 16600 1820 16652
rect 1860 16532 1912 16584
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 3240 16600 3292 16652
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5908 16600 5960 16652
rect 8300 16668 8352 16720
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 12072 16736 12124 16788
rect 13544 16736 13596 16788
rect 14556 16736 14608 16788
rect 15200 16736 15252 16788
rect 12716 16668 12768 16720
rect 16120 16668 16172 16720
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 7748 16600 7800 16652
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 12624 16643 12676 16652
rect 12624 16609 12633 16643
rect 12633 16609 12667 16643
rect 12667 16609 12676 16643
rect 12624 16600 12676 16609
rect 13636 16600 13688 16652
rect 15292 16643 15344 16652
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 4528 16532 4580 16584
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 5172 16532 5224 16584
rect 6276 16532 6328 16584
rect 6828 16532 6880 16584
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 9864 16532 9916 16584
rect 12072 16575 12124 16584
rect 10140 16464 10192 16516
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 13728 16575 13780 16584
rect 12164 16532 12216 16541
rect 13728 16541 13737 16575
rect 13737 16541 13771 16575
rect 13771 16541 13780 16575
rect 13728 16532 13780 16541
rect 9036 16439 9088 16448
rect 3148 16396 3200 16405
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 11060 16439 11112 16448
rect 11060 16405 11069 16439
rect 11069 16405 11103 16439
rect 11103 16405 11112 16439
rect 11060 16396 11112 16405
rect 11244 16396 11296 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2412 16192 2464 16244
rect 2044 16099 2096 16108
rect 2044 16065 2053 16099
rect 2053 16065 2087 16099
rect 2087 16065 2096 16099
rect 2044 16056 2096 16065
rect 5080 16192 5132 16244
rect 5172 16192 5224 16244
rect 6000 16192 6052 16244
rect 6276 16235 6328 16244
rect 6276 16201 6285 16235
rect 6285 16201 6319 16235
rect 6319 16201 6328 16235
rect 6276 16192 6328 16201
rect 8300 16192 8352 16244
rect 9864 16192 9916 16244
rect 10324 16235 10376 16244
rect 10324 16201 10333 16235
rect 10333 16201 10367 16235
rect 10367 16201 10376 16235
rect 10324 16192 10376 16201
rect 11980 16192 12032 16244
rect 13728 16192 13780 16244
rect 4804 16167 4856 16176
rect 4804 16133 4813 16167
rect 4813 16133 4847 16167
rect 4847 16133 4856 16167
rect 4804 16124 4856 16133
rect 9956 16167 10008 16176
rect 9956 16133 9965 16167
rect 9965 16133 9999 16167
rect 9999 16133 10008 16167
rect 9956 16124 10008 16133
rect 4528 16056 4580 16108
rect 4712 16056 4764 16108
rect 6460 16056 6512 16108
rect 9312 16099 9364 16108
rect 9312 16065 9321 16099
rect 9321 16065 9355 16099
rect 9355 16065 9364 16099
rect 9312 16056 9364 16065
rect 11060 16056 11112 16108
rect 2688 15988 2740 16040
rect 2780 15988 2832 16040
rect 3424 16031 3476 16040
rect 3424 15997 3458 16031
rect 3458 15997 3476 16031
rect 3424 15988 3476 15997
rect 3884 15988 3936 16040
rect 5816 15988 5868 16040
rect 7012 15988 7064 16040
rect 9588 15988 9640 16040
rect 9772 15988 9824 16040
rect 10692 16031 10744 16040
rect 10692 15997 10701 16031
rect 10701 15997 10735 16031
rect 10735 15997 10744 16031
rect 10692 15988 10744 15997
rect 10968 15988 11020 16040
rect 11244 16031 11296 16040
rect 11244 15997 11253 16031
rect 11253 15997 11287 16031
rect 11287 15997 11296 16031
rect 11244 15988 11296 15997
rect 3792 15920 3844 15972
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 3516 15852 3568 15904
rect 7012 15852 7064 15904
rect 8392 15852 8444 15904
rect 10876 15920 10928 15972
rect 16488 16056 16540 16108
rect 12440 15988 12492 16040
rect 13636 15988 13688 16040
rect 15292 16031 15344 16040
rect 15292 15997 15301 16031
rect 15301 15997 15335 16031
rect 15335 15997 15344 16031
rect 15292 15988 15344 15997
rect 15476 16031 15528 16040
rect 15476 15997 15485 16031
rect 15485 15997 15519 16031
rect 15519 15997 15528 16031
rect 15476 15988 15528 15997
rect 13084 15920 13136 15972
rect 13820 15920 13872 15972
rect 10048 15852 10100 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 13544 15852 13596 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2320 15691 2372 15700
rect 2320 15657 2329 15691
rect 2329 15657 2363 15691
rect 2363 15657 2372 15691
rect 2320 15648 2372 15657
rect 3332 15648 3384 15700
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 7748 15691 7800 15700
rect 7748 15657 7757 15691
rect 7757 15657 7791 15691
rect 7791 15657 7800 15691
rect 7748 15648 7800 15657
rect 8208 15648 8260 15700
rect 9588 15648 9640 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10140 15648 10192 15700
rect 10876 15691 10928 15700
rect 3424 15623 3476 15632
rect 3424 15589 3433 15623
rect 3433 15589 3467 15623
rect 3467 15589 3476 15623
rect 3424 15580 3476 15589
rect 10876 15657 10885 15691
rect 10885 15657 10919 15691
rect 10919 15657 10928 15691
rect 10876 15648 10928 15657
rect 12072 15648 12124 15700
rect 13820 15691 13872 15700
rect 13820 15657 13829 15691
rect 13829 15657 13863 15691
rect 13863 15657 13872 15691
rect 13820 15648 13872 15657
rect 16304 15580 16356 15632
rect 2780 15555 2832 15564
rect 2780 15521 2789 15555
rect 2789 15521 2823 15555
rect 2823 15521 2832 15555
rect 2780 15512 2832 15521
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 2596 15444 2648 15496
rect 3148 15444 3200 15496
rect 4160 15444 4212 15496
rect 5540 15512 5592 15564
rect 5816 15512 5868 15564
rect 6000 15555 6052 15564
rect 6000 15521 6034 15555
rect 6034 15521 6052 15555
rect 6000 15512 6052 15521
rect 8576 15512 8628 15564
rect 10784 15512 10836 15564
rect 11888 15512 11940 15564
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 10692 15444 10744 15496
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 11428 15444 11480 15496
rect 13820 15512 13872 15564
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16120 15512 16172 15521
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 3056 15376 3108 15428
rect 3516 15376 3568 15428
rect 3240 15308 3292 15360
rect 5448 15308 5500 15360
rect 7380 15308 7432 15360
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1492 15104 1544 15156
rect 2688 15104 2740 15156
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 3424 15011 3476 15020
rect 3424 14977 3433 15011
rect 3433 14977 3467 15011
rect 3467 14977 3476 15011
rect 3424 14968 3476 14977
rect 3792 14968 3844 15020
rect 5540 15104 5592 15156
rect 8300 15104 8352 15156
rect 10692 15147 10744 15156
rect 10692 15113 10701 15147
rect 10701 15113 10735 15147
rect 10735 15113 10744 15147
rect 10692 15104 10744 15113
rect 10968 15104 11020 15156
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 14188 15104 14240 15156
rect 8576 15079 8628 15088
rect 8576 15045 8585 15079
rect 8585 15045 8619 15079
rect 8619 15045 8628 15079
rect 8576 15036 8628 15045
rect 16120 15079 16172 15088
rect 16120 15045 16129 15079
rect 16129 15045 16163 15079
rect 16163 15045 16172 15079
rect 16120 15036 16172 15045
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 11428 15011 11480 15020
rect 11428 14977 11437 15011
rect 11437 14977 11471 15011
rect 11471 14977 11480 15011
rect 11428 14968 11480 14977
rect 2688 14832 2740 14884
rect 4068 14900 4120 14952
rect 5080 14900 5132 14952
rect 6828 14943 6880 14952
rect 6828 14909 6837 14943
rect 6837 14909 6871 14943
rect 6871 14909 6880 14943
rect 6828 14900 6880 14909
rect 9128 14900 9180 14952
rect 9680 14900 9732 14952
rect 11980 14900 12032 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 3700 14832 3752 14884
rect 4804 14832 4856 14884
rect 1860 14764 1912 14816
rect 2596 14764 2648 14816
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 6000 14764 6052 14816
rect 7380 14832 7432 14884
rect 13268 14832 13320 14884
rect 9496 14807 9548 14816
rect 9496 14773 9505 14807
rect 9505 14773 9539 14807
rect 9539 14773 9548 14807
rect 9496 14764 9548 14773
rect 10140 14764 10192 14816
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 11244 14807 11296 14816
rect 11244 14773 11253 14807
rect 11253 14773 11287 14807
rect 11287 14773 11296 14807
rect 11888 14807 11940 14816
rect 11244 14764 11296 14773
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 3424 14560 3476 14612
rect 3792 14560 3844 14612
rect 3976 14560 4028 14612
rect 4436 14603 4488 14612
rect 4436 14569 4445 14603
rect 4445 14569 4479 14603
rect 4479 14569 4488 14603
rect 4436 14560 4488 14569
rect 5724 14603 5776 14612
rect 5724 14569 5733 14603
rect 5733 14569 5767 14603
rect 5767 14569 5776 14603
rect 5724 14560 5776 14569
rect 7104 14560 7156 14612
rect 9496 14560 9548 14612
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11428 14603 11480 14612
rect 11428 14569 11437 14603
rect 11437 14569 11471 14603
rect 11471 14569 11480 14603
rect 11428 14560 11480 14569
rect 13268 14603 13320 14612
rect 13268 14569 13277 14603
rect 13277 14569 13311 14603
rect 13311 14569 13320 14603
rect 13268 14560 13320 14569
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 1492 14424 1544 14476
rect 2872 14424 2924 14476
rect 3884 14467 3936 14476
rect 3884 14433 3893 14467
rect 3893 14433 3927 14467
rect 3927 14433 3936 14467
rect 3884 14424 3936 14433
rect 3976 14424 4028 14476
rect 4620 14399 4672 14408
rect 4620 14365 4629 14399
rect 4629 14365 4663 14399
rect 4663 14365 4672 14399
rect 4620 14356 4672 14365
rect 2504 14288 2556 14340
rect 6460 14424 6512 14476
rect 8944 14492 8996 14544
rect 11796 14492 11848 14544
rect 13544 14492 13596 14544
rect 14188 14492 14240 14544
rect 8208 14424 8260 14476
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 5816 14356 5868 14408
rect 6368 14356 6420 14408
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 8484 14399 8536 14408
rect 6736 14356 6788 14365
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 9036 14356 9088 14408
rect 11888 14399 11940 14408
rect 5264 14263 5316 14272
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 6184 14263 6236 14272
rect 6184 14229 6193 14263
rect 6193 14229 6227 14263
rect 6227 14229 6236 14263
rect 6184 14220 6236 14229
rect 6368 14220 6420 14272
rect 6736 14220 6788 14272
rect 7380 14220 7432 14272
rect 8392 14220 8444 14272
rect 10048 14220 10100 14272
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 11888 14220 11940 14272
rect 13544 14220 13596 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 3700 14059 3752 14068
rect 3700 14025 3709 14059
rect 3709 14025 3743 14059
rect 3743 14025 3752 14059
rect 3700 14016 3752 14025
rect 4436 14016 4488 14068
rect 4620 14059 4672 14068
rect 4620 14025 4629 14059
rect 4629 14025 4663 14059
rect 4663 14025 4672 14059
rect 4620 14016 4672 14025
rect 5540 14016 5592 14068
rect 6644 14016 6696 14068
rect 7932 14016 7984 14068
rect 8300 14016 8352 14068
rect 9772 14016 9824 14068
rect 11244 14016 11296 14068
rect 13544 14059 13596 14068
rect 13544 14025 13553 14059
rect 13553 14025 13587 14059
rect 13587 14025 13596 14059
rect 13544 14016 13596 14025
rect 2872 13948 2924 14000
rect 4804 13948 4856 14000
rect 5264 13948 5316 14000
rect 5448 13880 5500 13932
rect 6460 13948 6512 14000
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 11796 13991 11848 14000
rect 11796 13957 11805 13991
rect 11805 13957 11839 13991
rect 11839 13957 11848 13991
rect 11796 13948 11848 13957
rect 6920 13880 6972 13932
rect 7380 13923 7432 13932
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 9036 13923 9088 13932
rect 9036 13889 9045 13923
rect 9045 13889 9079 13923
rect 9079 13889 9088 13923
rect 9036 13880 9088 13889
rect 12900 13923 12952 13932
rect 12900 13889 12909 13923
rect 12909 13889 12943 13923
rect 12943 13889 12952 13923
rect 12900 13880 12952 13889
rect 13268 13880 13320 13932
rect 14372 13880 14424 13932
rect 17868 13880 17920 13932
rect 1584 13855 1636 13864
rect 1584 13821 1593 13855
rect 1593 13821 1627 13855
rect 1627 13821 1636 13855
rect 1584 13812 1636 13821
rect 2504 13744 2556 13796
rect 2780 13676 2832 13728
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 6184 13812 6236 13864
rect 8208 13812 8260 13864
rect 5724 13744 5776 13796
rect 8392 13812 8444 13864
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 16672 13855 16724 13864
rect 16672 13821 16681 13855
rect 16681 13821 16715 13855
rect 16715 13821 16724 13855
rect 16672 13812 16724 13821
rect 9588 13744 9640 13796
rect 12532 13744 12584 13796
rect 6000 13676 6052 13728
rect 10048 13676 10100 13728
rect 11244 13719 11296 13728
rect 11244 13685 11253 13719
rect 11253 13685 11287 13719
rect 11287 13685 11296 13719
rect 11244 13676 11296 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2504 13515 2556 13524
rect 2504 13481 2513 13515
rect 2513 13481 2547 13515
rect 2547 13481 2556 13515
rect 2504 13472 2556 13481
rect 2596 13472 2648 13524
rect 2872 13447 2924 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2872 13413 2881 13447
rect 2881 13413 2915 13447
rect 2915 13413 2924 13447
rect 2872 13404 2924 13413
rect 5172 13472 5224 13524
rect 5264 13515 5316 13524
rect 5264 13481 5273 13515
rect 5273 13481 5307 13515
rect 5307 13481 5316 13515
rect 5264 13472 5316 13481
rect 5540 13472 5592 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 8484 13472 8536 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 9956 13472 10008 13524
rect 11244 13472 11296 13524
rect 11888 13472 11940 13524
rect 12532 13515 12584 13524
rect 12532 13481 12541 13515
rect 12541 13481 12575 13515
rect 12575 13481 12584 13515
rect 12532 13472 12584 13481
rect 13268 13472 13320 13524
rect 7288 13404 7340 13456
rect 8300 13404 8352 13456
rect 9864 13404 9916 13456
rect 17592 13404 17644 13456
rect 6552 13336 6604 13388
rect 8116 13336 8168 13388
rect 8576 13336 8628 13388
rect 10048 13336 10100 13388
rect 17408 13379 17460 13388
rect 2872 13268 2924 13320
rect 4068 13268 4120 13320
rect 4804 13311 4856 13320
rect 3976 13200 4028 13252
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 17408 13345 17417 13379
rect 17417 13345 17451 13379
rect 17451 13345 17460 13379
rect 17408 13336 17460 13345
rect 12440 13268 12492 13320
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 6920 13132 6972 13184
rect 9588 13200 9640 13252
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 1676 12928 1728 12980
rect 1768 12928 1820 12980
rect 4896 12928 4948 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 6552 12971 6604 12980
rect 6552 12937 6561 12971
rect 6561 12937 6595 12971
rect 6595 12937 6604 12971
rect 6552 12928 6604 12937
rect 8484 12928 8536 12980
rect 9864 12928 9916 12980
rect 10968 12928 11020 12980
rect 11888 12928 11940 12980
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 17408 12971 17460 12980
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 4160 12860 4212 12912
rect 6276 12903 6328 12912
rect 1584 12792 1636 12844
rect 5724 12835 5776 12844
rect 5724 12801 5733 12835
rect 5733 12801 5767 12835
rect 5767 12801 5776 12835
rect 5724 12792 5776 12801
rect 6276 12869 6285 12903
rect 6285 12869 6319 12903
rect 6319 12869 6328 12903
rect 6276 12860 6328 12869
rect 8208 12903 8260 12912
rect 8208 12869 8217 12903
rect 8217 12869 8251 12903
rect 8251 12869 8260 12903
rect 8208 12860 8260 12869
rect 13820 12903 13872 12912
rect 13820 12869 13829 12903
rect 13829 12869 13863 12903
rect 13863 12869 13872 12903
rect 13820 12860 13872 12869
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 2596 12724 2648 12776
rect 2780 12767 2832 12776
rect 2780 12733 2814 12767
rect 2814 12733 2832 12767
rect 2780 12724 2832 12733
rect 4804 12724 4856 12776
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 5264 12724 5316 12776
rect 6184 12724 6236 12776
rect 6920 12724 6972 12776
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 10140 12724 10192 12776
rect 10692 12724 10744 12776
rect 12532 12724 12584 12776
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 3148 12656 3200 12708
rect 4896 12656 4948 12708
rect 7748 12656 7800 12708
rect 9404 12699 9456 12708
rect 9404 12665 9413 12699
rect 9413 12665 9447 12699
rect 9447 12665 9456 12699
rect 9404 12656 9456 12665
rect 10784 12656 10836 12708
rect 12256 12699 12308 12708
rect 12256 12665 12265 12699
rect 12265 12665 12299 12699
rect 12299 12665 12308 12699
rect 12256 12656 12308 12665
rect 1860 12588 1912 12640
rect 2688 12588 2740 12640
rect 3240 12588 3292 12640
rect 10876 12588 10928 12640
rect 12348 12588 12400 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 4068 12384 4120 12436
rect 5448 12384 5500 12436
rect 6368 12384 6420 12436
rect 6920 12384 6972 12436
rect 8944 12384 8996 12436
rect 9956 12427 10008 12436
rect 9956 12393 9965 12427
rect 9965 12393 9999 12427
rect 9999 12393 10008 12427
rect 9956 12384 10008 12393
rect 10048 12384 10100 12436
rect 12256 12427 12308 12436
rect 12256 12393 12265 12427
rect 12265 12393 12299 12427
rect 12299 12393 12308 12427
rect 12256 12384 12308 12393
rect 12440 12384 12492 12436
rect 13084 12384 13136 12436
rect 14648 12427 14700 12436
rect 14648 12393 14657 12427
rect 14657 12393 14691 12427
rect 14691 12393 14700 12427
rect 14648 12384 14700 12393
rect 20996 12384 21048 12436
rect 6460 12316 6512 12368
rect 8300 12359 8352 12368
rect 8300 12325 8309 12359
rect 8309 12325 8343 12359
rect 8343 12325 8352 12359
rect 8300 12316 8352 12325
rect 11152 12359 11204 12368
rect 11152 12325 11186 12359
rect 11186 12325 11204 12359
rect 11152 12316 11204 12325
rect 13544 12359 13596 12368
rect 2596 12248 2648 12300
rect 4436 12248 4488 12300
rect 1400 12180 1452 12232
rect 5724 12248 5776 12300
rect 6644 12248 6696 12300
rect 9772 12248 9824 12300
rect 11888 12248 11940 12300
rect 5908 12180 5960 12232
rect 2780 12112 2832 12164
rect 8116 12155 8168 12164
rect 8116 12121 8125 12155
rect 8125 12121 8159 12155
rect 8159 12121 8168 12155
rect 8116 12112 8168 12121
rect 1768 12044 1820 12096
rect 2688 12044 2740 12096
rect 2872 12044 2924 12096
rect 3700 12044 3752 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 9404 12044 9456 12096
rect 9864 12044 9916 12096
rect 11244 12044 11296 12096
rect 12532 12180 12584 12232
rect 13544 12325 13553 12359
rect 13553 12325 13587 12359
rect 13587 12325 13596 12359
rect 13544 12316 13596 12325
rect 20812 12316 20864 12368
rect 13452 12180 13504 12232
rect 14648 12112 14700 12164
rect 13728 12044 13780 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1400 11840 1452 11892
rect 1676 11704 1728 11756
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 4068 11840 4120 11892
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 6460 11840 6512 11892
rect 6736 11840 6788 11892
rect 4896 11772 4948 11824
rect 5080 11772 5132 11824
rect 6000 11704 6052 11756
rect 8576 11704 8628 11756
rect 2780 11636 2832 11688
rect 3056 11636 3108 11688
rect 5264 11636 5316 11688
rect 6092 11636 6144 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 8300 11636 8352 11688
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 9220 11840 9272 11892
rect 11152 11840 11204 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 13544 11840 13596 11892
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 3240 11611 3292 11620
rect 3240 11577 3274 11611
rect 3274 11577 3292 11611
rect 3240 11568 3292 11577
rect 3608 11568 3660 11620
rect 1584 11500 1636 11552
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 2596 11500 2648 11552
rect 3332 11500 3384 11552
rect 4436 11500 4488 11552
rect 9680 11568 9732 11620
rect 10048 11568 10100 11620
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11296 1728 11348
rect 3976 11296 4028 11348
rect 5264 11339 5316 11348
rect 5264 11305 5273 11339
rect 5273 11305 5307 11339
rect 5307 11305 5316 11339
rect 5264 11296 5316 11305
rect 6644 11296 6696 11348
rect 6828 11296 6880 11348
rect 10048 11296 10100 11348
rect 11244 11296 11296 11348
rect 2596 11228 2648 11280
rect 8852 11228 8904 11280
rect 9588 11228 9640 11280
rect 21180 11228 21232 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 3240 11160 3292 11212
rect 3700 11160 3752 11212
rect 4160 11160 4212 11212
rect 5540 11160 5592 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 9772 11160 9824 11212
rect 19524 11203 19576 11212
rect 19524 11169 19533 11203
rect 19533 11169 19567 11203
rect 19567 11169 19576 11203
rect 19524 11160 19576 11169
rect 4068 11092 4120 11144
rect 6000 11024 6052 11076
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 7104 11092 7156 11144
rect 6368 11024 6420 11076
rect 7840 11067 7892 11076
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 3884 10999 3936 11008
rect 3884 10965 3893 10999
rect 3893 10965 3927 10999
rect 3927 10965 3936 10999
rect 3884 10956 3936 10965
rect 8484 10956 8536 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 4160 10752 4212 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 1584 10616 1636 10668
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 8208 10752 8260 10804
rect 9588 10795 9640 10804
rect 9588 10761 9597 10795
rect 9597 10761 9631 10795
rect 9631 10761 9640 10795
rect 9588 10752 9640 10761
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 10048 10684 10100 10736
rect 1768 10548 1820 10600
rect 10692 10616 10744 10668
rect 19248 10616 19300 10668
rect 19984 10616 20036 10668
rect 2780 10548 2832 10600
rect 3976 10591 4028 10600
rect 3976 10557 3985 10591
rect 3985 10557 4019 10591
rect 4019 10557 4028 10591
rect 3976 10548 4028 10557
rect 8484 10591 8536 10600
rect 8484 10557 8518 10591
rect 8518 10557 8536 10591
rect 1492 10455 1544 10464
rect 1492 10421 1501 10455
rect 1501 10421 1535 10455
rect 1535 10421 1544 10455
rect 1492 10412 1544 10421
rect 1584 10412 1636 10464
rect 3884 10480 3936 10532
rect 6000 10480 6052 10532
rect 8484 10548 8536 10557
rect 9772 10548 9824 10600
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 19524 10548 19576 10600
rect 9496 10480 9548 10532
rect 3240 10412 3292 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 5540 10412 5592 10464
rect 6184 10412 6236 10464
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 4068 10251 4120 10260
rect 4068 10217 4077 10251
rect 4077 10217 4111 10251
rect 4111 10217 4120 10251
rect 4068 10208 4120 10217
rect 4252 10208 4304 10260
rect 4988 10208 5040 10260
rect 8484 10208 8536 10260
rect 9864 10208 9916 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 1952 10140 2004 10192
rect 3976 10140 4028 10192
rect 6184 10140 6236 10192
rect 9496 10183 9548 10192
rect 9496 10149 9505 10183
rect 9505 10149 9539 10183
rect 9539 10149 9548 10183
rect 9496 10140 9548 10149
rect 9680 10140 9732 10192
rect 9956 10140 10008 10192
rect 1676 10115 1728 10124
rect 1676 10081 1710 10115
rect 1710 10081 1728 10115
rect 1676 10072 1728 10081
rect 3700 10072 3752 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 5080 10004 5132 10056
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 5172 9868 5224 9920
rect 9864 10004 9916 10056
rect 10140 10004 10192 10056
rect 9680 9979 9732 9988
rect 9680 9945 9689 9979
rect 9689 9945 9723 9979
rect 9723 9945 9732 9979
rect 9680 9936 9732 9945
rect 6368 9868 6420 9920
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 2504 9664 2556 9716
rect 3884 9664 3936 9716
rect 6368 9664 6420 9716
rect 8484 9707 8536 9716
rect 3976 9596 4028 9648
rect 5080 9596 5132 9648
rect 1400 9460 1452 9512
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 2688 9460 2740 9512
rect 3240 9528 3292 9580
rect 3056 9460 3108 9512
rect 3332 9460 3384 9512
rect 3700 9528 3752 9580
rect 3976 9460 4028 9512
rect 4344 9503 4396 9512
rect 4344 9469 4378 9503
rect 4378 9469 4396 9503
rect 8484 9673 8493 9707
rect 8493 9673 8527 9707
rect 8527 9673 8536 9707
rect 8484 9664 8536 9673
rect 9864 9664 9916 9716
rect 10048 9664 10100 9716
rect 9956 9528 10008 9580
rect 2780 9392 2832 9444
rect 4344 9460 4396 9469
rect 7380 9435 7432 9444
rect 7380 9401 7414 9435
rect 7414 9401 7432 9435
rect 7380 9392 7432 9401
rect 3332 9324 3384 9376
rect 3884 9324 3936 9376
rect 4436 9324 4488 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 1860 9120 1912 9172
rect 2596 9163 2648 9172
rect 2596 9129 2605 9163
rect 2605 9129 2639 9163
rect 2639 9129 2648 9163
rect 2596 9120 2648 9129
rect 3148 9120 3200 9172
rect 3792 9120 3844 9172
rect 4068 9163 4120 9172
rect 4068 9129 4077 9163
rect 4077 9129 4111 9163
rect 4111 9129 4120 9163
rect 4068 9120 4120 9129
rect 5264 9120 5316 9172
rect 6184 9120 6236 9172
rect 7104 9120 7156 9172
rect 7748 9163 7800 9172
rect 7748 9129 7757 9163
rect 7757 9129 7791 9163
rect 7791 9129 7800 9163
rect 7748 9120 7800 9129
rect 2320 9052 2372 9104
rect 3332 9052 3384 9104
rect 4344 9052 4396 9104
rect 5356 9095 5408 9104
rect 5356 9061 5390 9095
rect 5390 9061 5408 9095
rect 5356 9052 5408 9061
rect 6368 9052 6420 9104
rect 7656 9095 7708 9104
rect 7656 9061 7665 9095
rect 7665 9061 7699 9095
rect 7699 9061 7708 9095
rect 7656 9052 7708 9061
rect 2780 8984 2832 9036
rect 5080 9027 5132 9036
rect 5080 8993 5089 9027
rect 5089 8993 5123 9027
rect 5123 8993 5132 9027
rect 5080 8984 5132 8993
rect 2228 8916 2280 8968
rect 2504 8916 2556 8968
rect 7380 8848 7432 8900
rect 8024 8916 8076 8968
rect 2780 8780 2832 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2320 8576 2372 8628
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 3240 8576 3292 8628
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 6000 8576 6052 8628
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 7656 8508 7708 8560
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2780 8440 2832 8492
rect 3240 8440 3292 8492
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 3700 8372 3752 8424
rect 4528 8372 4580 8424
rect 5264 8372 5316 8424
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1860 8032 1912 8084
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 2964 8032 3016 8084
rect 3240 8032 3292 8084
rect 4620 8032 4672 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5540 8032 5592 8084
rect 2688 7964 2740 8016
rect 4160 7964 4212 8016
rect 2872 7896 2924 7948
rect 3608 7896 3660 7948
rect 3056 7871 3108 7880
rect 3056 7837 3065 7871
rect 3065 7837 3099 7871
rect 3099 7837 3108 7871
rect 3056 7828 3108 7837
rect 3976 7828 4028 7880
rect 4528 7828 4580 7880
rect 4068 7803 4120 7812
rect 4068 7769 4077 7803
rect 4077 7769 4111 7803
rect 4111 7769 4120 7803
rect 4068 7760 4120 7769
rect 4620 7692 4672 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1860 7488 1912 7540
rect 2780 7488 2832 7540
rect 2964 7488 3016 7540
rect 3056 7488 3108 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 23572 7488 23624 7540
rect 4620 7420 4672 7472
rect 22192 7327 22244 7336
rect 22192 7293 22201 7327
rect 22201 7293 22235 7327
rect 22235 7293 22244 7327
rect 22192 7284 22244 7293
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 22744 6851 22796 6860
rect 22744 6817 22753 6851
rect 22753 6817 22787 6851
rect 22787 6817 22796 6851
rect 22744 6808 22796 6817
rect 23388 6672 23440 6724
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 22744 6443 22796 6452
rect 22744 6409 22753 6443
rect 22753 6409 22787 6443
rect 22787 6409 22796 6443
rect 22744 6400 22796 6409
rect 25044 6400 25096 6452
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24768 5856 24820 5908
rect 23940 5763 23992 5772
rect 23940 5729 23949 5763
rect 23949 5729 23983 5763
rect 23983 5729 23992 5763
rect 23940 5720 23992 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 23940 5355 23992 5364
rect 23940 5321 23949 5355
rect 23949 5321 23983 5355
rect 23983 5321 23992 5355
rect 23940 5312 23992 5321
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 24492 5151 24544 5160
rect 24492 5117 24501 5151
rect 24501 5117 24535 5151
rect 24535 5117 24544 5151
rect 24492 5108 24544 5117
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24768 4811 24820 4820
rect 24768 4777 24777 4811
rect 24777 4777 24811 4811
rect 24811 4777 24820 4811
rect 24768 4768 24820 4777
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 7012 4088 7064 4140
rect 7472 4088 7524 4140
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3146 27520 3202 28000
rect 3514 27704 3570 27713
rect 3514 27639 3570 27648
rect 308 24449 336 27520
rect 294 24440 350 24449
rect 294 24375 350 24384
rect 860 18873 888 27520
rect 1412 26466 1440 27520
rect 1964 26874 1992 27520
rect 2516 26874 2544 27520
rect 1964 26846 2176 26874
rect 1412 26438 1532 26466
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1412 21593 1440 24550
rect 1398 21584 1454 21593
rect 1398 21519 1454 21528
rect 846 18864 902 18873
rect 846 18799 902 18808
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1412 16794 1440 18702
rect 1504 17066 1532 26438
rect 2044 25764 2096 25770
rect 2044 25706 2096 25712
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1596 23497 1624 25094
rect 1860 24608 1912 24614
rect 1860 24550 1912 24556
rect 1768 24200 1820 24206
rect 1766 24168 1768 24177
rect 1820 24168 1822 24177
rect 1766 24103 1822 24112
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1582 23488 1638 23497
rect 1582 23423 1638 23432
rect 1780 22642 1808 24006
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1872 22098 1900 24550
rect 1950 23624 2006 23633
rect 1950 23559 1952 23568
rect 2004 23559 2006 23568
rect 1952 23530 2004 23536
rect 2056 23254 2084 25706
rect 2044 23248 2096 23254
rect 2044 23190 2096 23196
rect 1584 22092 1636 22098
rect 1584 22034 1636 22040
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1596 21622 1624 22034
rect 1584 21616 1636 21622
rect 1584 21558 1636 21564
rect 1950 21040 2006 21049
rect 1950 20975 1952 20984
rect 2004 20975 2006 20984
rect 1952 20946 2004 20952
rect 1952 20868 2004 20874
rect 1952 20810 2004 20816
rect 1964 20262 1992 20810
rect 2148 20754 2176 26846
rect 2240 26846 2544 26874
rect 2240 23338 2268 26846
rect 2320 25356 2372 25362
rect 2320 25298 2372 25304
rect 2504 25356 2556 25362
rect 2504 25298 2556 25304
rect 2332 24614 2360 25298
rect 2412 24676 2464 24682
rect 2412 24618 2464 24624
rect 2320 24608 2372 24614
rect 2320 24550 2372 24556
rect 2424 23662 2452 24618
rect 2516 24070 2544 25298
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2596 24268 2648 24274
rect 2596 24210 2648 24216
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2502 23896 2558 23905
rect 2608 23882 2636 24210
rect 2558 23854 2636 23882
rect 2502 23831 2504 23840
rect 2556 23831 2558 23840
rect 2504 23802 2556 23808
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2240 23310 2360 23338
rect 2424 23322 2452 23598
rect 2700 23338 2728 24550
rect 2792 24041 2820 25094
rect 2870 24304 2926 24313
rect 2870 24239 2872 24248
rect 2924 24239 2926 24248
rect 2872 24210 2924 24216
rect 2778 24032 2834 24041
rect 2778 23967 2834 23976
rect 2884 23866 2912 24210
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2872 23860 2924 23866
rect 2872 23802 2924 23808
rect 2226 23216 2282 23225
rect 2226 23151 2282 23160
rect 2056 20726 2176 20754
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1582 17368 1638 17377
rect 1582 17303 1584 17312
rect 1636 17303 1638 17312
rect 1584 17274 1636 17280
rect 1688 17218 1716 18566
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1596 17190 1716 17218
rect 1596 17134 1624 17190
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1492 17060 1544 17066
rect 1492 17002 1544 17008
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1490 16688 1546 16697
rect 1490 16623 1546 16632
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 14657 1440 15438
rect 1504 15162 1532 16623
rect 1596 16561 1624 17070
rect 1780 16658 1808 17750
rect 1872 16946 1900 19654
rect 1964 19281 1992 20198
rect 2056 19417 2084 20726
rect 2240 20618 2268 23151
rect 2332 20890 2360 23310
rect 2412 23316 2464 23322
rect 2700 23310 2820 23338
rect 2412 23258 2464 23264
rect 2688 23180 2740 23186
rect 2688 23122 2740 23128
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2502 23080 2558 23089
rect 2424 22438 2452 23054
rect 2502 23015 2558 23024
rect 2516 22574 2544 23015
rect 2700 22710 2728 23122
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2504 22568 2556 22574
rect 2504 22510 2556 22516
rect 2412 22432 2464 22438
rect 2410 22400 2412 22409
rect 2464 22400 2466 22409
rect 2410 22335 2466 22344
rect 2516 22234 2544 22510
rect 2700 22234 2728 22646
rect 2504 22228 2556 22234
rect 2504 22170 2556 22176
rect 2688 22228 2740 22234
rect 2688 22170 2740 22176
rect 2410 22128 2466 22137
rect 2410 22063 2466 22072
rect 2424 21690 2452 22063
rect 2412 21684 2464 21690
rect 2412 21626 2464 21632
rect 2424 21486 2452 21626
rect 2792 21622 2820 23310
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2688 21616 2740 21622
rect 2688 21558 2740 21564
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2412 21480 2464 21486
rect 2412 21422 2464 21428
rect 2700 20913 2728 21558
rect 2686 20904 2742 20913
rect 2332 20862 2636 20890
rect 2320 20800 2372 20806
rect 2320 20742 2372 20748
rect 2148 20590 2268 20618
rect 2148 20466 2176 20590
rect 2332 20482 2360 20742
rect 2412 20528 2464 20534
rect 2240 20466 2360 20482
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2228 20460 2360 20466
rect 2280 20454 2360 20460
rect 2228 20402 2280 20408
rect 2332 20058 2360 20454
rect 2410 20496 2412 20505
rect 2464 20496 2466 20505
rect 2410 20431 2466 20440
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2240 19718 2268 19858
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2042 19408 2098 19417
rect 2042 19343 2098 19352
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1964 17610 1992 18090
rect 2148 18086 2176 19110
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2240 17882 2268 19654
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2332 18222 2360 19246
rect 2424 18970 2452 19790
rect 2504 19780 2556 19786
rect 2504 19722 2556 19728
rect 2516 19242 2544 19722
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1872 16918 2084 16946
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1860 16584 1912 16590
rect 1582 16552 1638 16561
rect 1860 16526 1912 16532
rect 1582 16487 1638 16496
rect 1674 16144 1730 16153
rect 1674 16079 1730 16088
rect 1582 16008 1638 16017
rect 1582 15943 1638 15952
rect 1596 15910 1624 15943
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1398 14648 1454 14657
rect 1398 14583 1454 14592
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 14362 1532 14418
rect 1504 14334 1624 14362
rect 1596 13870 1624 14334
rect 1584 13864 1636 13870
rect 1584 13806 1636 13812
rect 1596 12850 1624 13806
rect 1688 12986 1716 16079
rect 1872 15502 1900 16526
rect 2056 16114 2084 16918
rect 2332 16590 2360 18022
rect 2608 17513 2636 20862
rect 2686 20839 2742 20848
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 2792 20330 2820 20742
rect 2884 20369 2912 22918
rect 2976 22817 3004 24006
rect 2962 22808 3018 22817
rect 2962 22743 3018 22752
rect 3054 22264 3110 22273
rect 3054 22199 3110 22208
rect 3068 21962 3096 22199
rect 3056 21956 3108 21962
rect 3056 21898 3108 21904
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 2976 21146 3004 21247
rect 2964 21140 3016 21146
rect 2964 21082 3016 21088
rect 3056 20460 3108 20466
rect 3056 20402 3108 20408
rect 2870 20360 2926 20369
rect 2780 20324 2832 20330
rect 2870 20295 2926 20304
rect 2780 20266 2832 20272
rect 2792 19700 2820 20266
rect 2700 19672 2820 19700
rect 2700 17882 2728 19672
rect 2962 19408 3018 19417
rect 2962 19343 3018 19352
rect 2976 18902 3004 19343
rect 3068 19174 3096 20402
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 2964 18896 3016 18902
rect 2870 18864 2926 18873
rect 2964 18838 3016 18844
rect 2870 18799 2872 18808
rect 2924 18799 2926 18808
rect 2872 18770 2924 18776
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2792 18193 2820 18702
rect 2884 18426 2912 18770
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2778 18184 2834 18193
rect 2976 18154 3004 18838
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2778 18119 2834 18128
rect 2964 18148 3016 18154
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2594 17504 2650 17513
rect 2594 17439 2650 17448
rect 2594 17368 2650 17377
rect 2594 17303 2650 17312
rect 2608 17134 2636 17303
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2320 16584 2372 16590
rect 2320 16526 2372 16532
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2332 15706 2360 16526
rect 2424 16250 2452 16730
rect 2608 16402 2636 17070
rect 2700 16998 2728 17682
rect 2792 17610 2820 18119
rect 2964 18090 3016 18096
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 2688 16992 2740 16998
rect 2688 16934 2740 16940
rect 2700 16726 2728 16934
rect 2792 16794 2820 17546
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2688 16720 2740 16726
rect 2688 16662 2740 16668
rect 2608 16374 2820 16402
rect 2412 16244 2464 16250
rect 2412 16186 2464 16192
rect 2792 16046 2820 16374
rect 2688 16040 2740 16046
rect 2688 15982 2740 15988
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1860 15496 1912 15502
rect 1858 15464 1860 15473
rect 2596 15496 2648 15502
rect 1912 15464 1914 15473
rect 2596 15438 2648 15444
rect 1858 15399 1914 15408
rect 2608 14822 2636 15438
rect 2700 15162 2728 15982
rect 2976 15586 3004 18090
rect 2792 15570 3004 15586
rect 2780 15564 3004 15570
rect 2832 15558 3004 15564
rect 2780 15506 2832 15512
rect 2688 15156 2740 15162
rect 2688 15098 2740 15104
rect 2688 14884 2740 14890
rect 2688 14826 2740 14832
rect 1860 14816 1912 14822
rect 1860 14758 1912 14764
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1780 13161 1808 13330
rect 1872 13326 1900 14758
rect 2700 14634 2728 14826
rect 2792 14634 2820 15506
rect 3068 15434 3096 18362
rect 3160 17882 3188 27520
rect 3528 26382 3556 27639
rect 3698 27520 3754 28000
rect 4250 27520 4306 28000
rect 4802 27520 4858 28000
rect 5354 27520 5410 28000
rect 5998 27520 6054 28000
rect 6550 27520 6606 28000
rect 7102 27520 7158 28000
rect 7654 27520 7710 28000
rect 8206 27520 8262 28000
rect 8850 27520 8906 28000
rect 9402 27520 9458 28000
rect 9954 27520 10010 28000
rect 10506 27520 10562 28000
rect 11058 27520 11114 28000
rect 11702 27520 11758 28000
rect 12254 27520 12310 28000
rect 12806 27520 12862 28000
rect 13358 27520 13414 28000
rect 13910 27520 13966 28000
rect 14554 27520 14610 28000
rect 15106 27520 15162 28000
rect 15658 27520 15714 28000
rect 16210 27520 16266 28000
rect 16762 27520 16818 28000
rect 17406 27520 17462 28000
rect 17958 27520 18014 28000
rect 18510 27520 18566 28000
rect 19062 27520 19118 28000
rect 19614 27520 19670 28000
rect 20258 27520 20314 28000
rect 20810 27520 20866 28000
rect 21362 27520 21418 28000
rect 21914 27520 21970 28000
rect 22466 27520 22522 28000
rect 23110 27520 23166 28000
rect 23662 27520 23718 28000
rect 24214 27520 24270 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 3516 26376 3568 26382
rect 3516 26318 3568 26324
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3528 24750 3556 25638
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 3620 24818 3648 25094
rect 3608 24812 3660 24818
rect 3608 24754 3660 24760
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3620 24410 3648 24754
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3712 23202 3740 27520
rect 4066 27160 4122 27169
rect 4066 27095 4122 27104
rect 4080 26858 4108 27095
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4066 26480 4122 26489
rect 4066 26415 4068 26424
rect 4120 26415 4122 26424
rect 4068 26386 4120 26392
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4080 25430 4108 25871
rect 4068 25424 4120 25430
rect 4068 25366 4120 25372
rect 4160 25288 4212 25294
rect 4066 25256 4122 25265
rect 4160 25230 4212 25236
rect 4066 25191 4122 25200
rect 4080 24886 4108 25191
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 4172 24614 4200 25230
rect 4264 24834 4292 27520
rect 4816 27418 4844 27520
rect 4816 27390 5304 27418
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 4264 24806 4568 24834
rect 4724 24818 4752 25162
rect 4160 24608 4212 24614
rect 4160 24550 4212 24556
rect 4068 24268 4120 24274
rect 4068 24210 4120 24216
rect 4080 23662 4108 24210
rect 4172 24070 4200 24550
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 3620 23174 3740 23202
rect 4080 23186 4108 23598
rect 4172 23594 4200 24006
rect 4160 23588 4212 23594
rect 4160 23530 4212 23536
rect 4068 23180 4120 23186
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3528 22234 3556 22578
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3528 21486 3556 21517
rect 3516 21480 3568 21486
rect 3514 21448 3516 21457
rect 3568 21448 3570 21457
rect 3514 21383 3570 21392
rect 3528 21146 3556 21383
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3516 19780 3568 19786
rect 3516 19722 3568 19728
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3160 17338 3188 17818
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3160 17218 3188 17274
rect 3160 17190 3280 17218
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16454 3188 17002
rect 3252 16794 3280 17190
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 15502 3188 16390
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 2700 14606 3004 14634
rect 3160 14618 3188 15438
rect 3252 15366 3280 16594
rect 3344 15706 3372 17478
rect 3436 16164 3464 18566
rect 3528 16232 3556 19722
rect 3620 17814 3648 23174
rect 4068 23122 4120 23128
rect 3698 22536 3754 22545
rect 3698 22471 3700 22480
rect 3752 22471 3754 22480
rect 3700 22442 3752 22448
rect 4080 22166 4108 23122
rect 4252 22568 4304 22574
rect 4252 22510 4304 22516
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 3712 22001 3740 22034
rect 4068 22024 4120 22030
rect 3698 21992 3754 22001
rect 4068 21966 4120 21972
rect 3698 21927 3754 21936
rect 3712 21690 3740 21927
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 3896 20262 3924 20742
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 19854 3924 20198
rect 3884 19848 3936 19854
rect 3988 19825 4016 21286
rect 4080 21010 4108 21966
rect 4264 21894 4292 22510
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4356 21690 4384 22034
rect 4436 21888 4488 21894
rect 4436 21830 4488 21836
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4172 21486 4200 21558
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4448 21078 4476 21830
rect 4436 21072 4488 21078
rect 4436 21014 4488 21020
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4448 20602 4476 21014
rect 4436 20596 4488 20602
rect 4436 20538 4488 20544
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 20097 4108 20198
rect 4066 20088 4122 20097
rect 4066 20023 4122 20032
rect 4158 19952 4214 19961
rect 4158 19887 4160 19896
rect 4212 19887 4214 19896
rect 4160 19858 4212 19864
rect 3884 19790 3936 19796
rect 3974 19816 4030 19825
rect 3974 19751 4030 19760
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3804 18630 3832 19654
rect 3976 19168 4028 19174
rect 4080 19145 4108 19654
rect 4172 19310 4200 19858
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3976 19110 4028 19116
rect 4066 19136 4122 19145
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3698 18048 3754 18057
rect 3698 17983 3754 17992
rect 3608 17808 3660 17814
rect 3608 17750 3660 17756
rect 3528 16204 3648 16232
rect 3436 16136 3556 16164
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15638 3464 15982
rect 3528 15910 3556 16136
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15026 3280 15302
rect 3436 15026 3464 15574
rect 3528 15434 3556 15846
rect 3516 15428 3568 15434
rect 3516 15370 3568 15376
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3436 14618 3464 14962
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2516 13802 2544 14282
rect 2884 14006 2912 14418
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2516 13530 2544 13738
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1766 13152 1822 13161
rect 1766 13087 1822 13096
rect 1780 12986 1808 13087
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1872 12646 1900 13262
rect 2608 12782 2636 13466
rect 2792 12782 2820 13670
rect 2884 13462 2912 13942
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12481 2728 12582
rect 2502 12472 2558 12481
rect 2502 12407 2558 12416
rect 2686 12472 2742 12481
rect 2686 12407 2742 12416
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11898 1440 12174
rect 1768 12096 1820 12102
rect 2516 12050 2544 12407
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 1768 12038 1820 12044
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1412 11218 1440 11834
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1596 10674 1624 11494
rect 1688 11354 1716 11698
rect 1780 11558 1808 12038
rect 2332 12022 2544 12050
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1490 10568 1546 10577
rect 1490 10503 1546 10512
rect 1504 10470 1532 10503
rect 1492 10464 1544 10470
rect 1492 10406 1544 10412
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1596 8498 1624 10406
rect 1688 10130 1716 11290
rect 1780 11257 1808 11494
rect 1766 11248 1822 11257
rect 1766 11183 1822 11192
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1688 9178 1716 10066
rect 1780 9722 1808 10542
rect 1964 10198 1992 10610
rect 1952 10192 2004 10198
rect 1952 10134 2004 10140
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1872 9178 1900 9454
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1872 8090 1900 9114
rect 2332 9110 2360 12022
rect 2502 11792 2558 11801
rect 2502 11727 2504 11736
rect 2556 11727 2558 11736
rect 2504 11698 2556 11704
rect 2608 11558 2636 12242
rect 2792 12170 2820 12718
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11286 2636 11494
rect 2596 11280 2648 11286
rect 2596 11222 2648 11228
rect 2700 9874 2728 12038
rect 2792 11694 2820 12106
rect 2884 12102 2912 13262
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2870 11928 2926 11937
rect 2870 11863 2926 11872
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10266 2820 10542
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2516 9846 2728 9874
rect 2516 9722 2544 9846
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2608 9710 2820 9738
rect 2608 9602 2636 9710
rect 2792 9625 2820 9710
rect 2516 9574 2636 9602
rect 2778 9616 2834 9625
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2240 8090 2268 8910
rect 2332 8634 2360 9046
rect 2516 8974 2544 9574
rect 2778 9551 2834 9560
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2608 8634 2636 9114
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2594 8528 2650 8537
rect 2594 8463 2650 8472
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1872 7546 1900 8026
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 2608 2689 2636 8463
rect 2700 8022 2728 9454
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 9042 2820 9386
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8498 2820 8774
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2884 7954 2912 11863
rect 2976 8090 3004 14606
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3424 14612 3476 14618
rect 3424 14554 3476 14560
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3068 9625 3096 11630
rect 3054 9616 3110 9625
rect 3054 9551 3110 9560
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2884 7562 2912 7890
rect 2792 7546 2912 7562
rect 2976 7546 3004 8026
rect 3068 7886 3096 9454
rect 3160 9178 3188 12650
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 3252 11626 3280 12582
rect 3620 12424 3648 16204
rect 3712 15065 3740 17983
rect 3804 17377 3832 18566
rect 3896 17678 3924 18770
rect 3988 18154 4016 19110
rect 4066 19071 4122 19080
rect 4252 18624 4304 18630
rect 4250 18592 4252 18601
rect 4304 18592 4306 18601
rect 4250 18527 4306 18536
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 4250 17912 4306 17921
rect 4250 17847 4252 17856
rect 4304 17847 4306 17856
rect 4252 17818 4304 17824
rect 4066 17776 4122 17785
rect 4122 17720 4200 17728
rect 4066 17711 4068 17720
rect 4120 17700 4200 17720
rect 4068 17682 4120 17688
rect 3884 17672 3936 17678
rect 3882 17640 3884 17649
rect 3936 17640 3938 17649
rect 3882 17575 3938 17584
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 3790 17368 3846 17377
rect 3790 17303 3846 17312
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3896 16794 3924 16934
rect 4080 16794 4108 17546
rect 4172 17338 4200 17700
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4436 16788 4488 16794
rect 4540 16776 4568 24806
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4620 24744 4672 24750
rect 4620 24686 4672 24692
rect 4632 24410 4660 24686
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4620 23724 4672 23730
rect 4620 23666 4672 23672
rect 4632 22658 4660 23666
rect 4724 23526 4752 24754
rect 4908 24614 4936 25298
rect 5000 24954 5028 25298
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 5080 24812 5132 24818
rect 5080 24754 5132 24760
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4724 23254 4752 23462
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 4724 22778 4752 23190
rect 4712 22772 4764 22778
rect 4712 22714 4764 22720
rect 4632 22630 4752 22658
rect 4618 19272 4674 19281
rect 4618 19207 4674 19216
rect 4632 19174 4660 19207
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4632 17882 4660 18090
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4488 16748 4568 16776
rect 4436 16730 4488 16736
rect 3896 16046 3924 16730
rect 3884 16040 3936 16046
rect 3884 15982 3936 15988
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3698 15056 3754 15065
rect 3804 15026 3832 15914
rect 3974 15056 4030 15065
rect 3698 14991 3754 15000
rect 3792 15020 3844 15026
rect 3974 14991 4030 15000
rect 3792 14962 3844 14968
rect 3698 14920 3754 14929
rect 3698 14855 3700 14864
rect 3752 14855 3754 14864
rect 3700 14826 3752 14832
rect 3712 14074 3740 14826
rect 3804 14618 3832 14962
rect 3988 14618 4016 14991
rect 4080 14958 4108 16730
rect 4252 16720 4304 16726
rect 4252 16662 4304 16668
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4172 14822 4200 15438
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3882 14512 3938 14521
rect 3882 14447 3884 14456
rect 3936 14447 3938 14456
rect 3976 14476 4028 14482
rect 3884 14418 3936 14424
rect 3976 14418 4028 14424
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3436 12396 3648 12424
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10470 3280 11154
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3252 9586 3280 10406
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3344 9518 3372 11494
rect 3332 9512 3384 9518
rect 3238 9480 3294 9489
rect 3332 9454 3384 9460
rect 3238 9415 3294 9424
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3252 8634 3280 9415
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 9110 3372 9318
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3252 8090 3280 8434
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 3068 7546 3096 7822
rect 2780 7540 2912 7546
rect 2832 7534 2912 7540
rect 2964 7540 3016 7546
rect 2780 7482 2832 7488
rect 2964 7482 3016 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3436 6882 3464 12396
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3608 11620 3660 11626
rect 3608 11562 3660 11568
rect 3620 8498 3648 11562
rect 3712 11218 3740 12038
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3698 10704 3754 10713
rect 3698 10639 3754 10648
rect 3712 10130 3740 10639
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9586 3740 10066
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3804 9178 3832 13670
rect 3988 13258 4016 14418
rect 4172 14385 4200 14758
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 4158 13424 4214 13433
rect 4158 13359 4214 13368
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4080 12442 4108 13262
rect 4172 13258 4200 13359
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4172 12322 4200 12854
rect 4080 12294 4200 12322
rect 4080 11898 4108 12294
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10538 3924 10950
rect 3988 10713 4016 11290
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3896 9926 3924 10474
rect 3988 10441 4016 10542
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 4080 10266 4108 11086
rect 4172 10810 4200 11154
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3976 10192 4028 10198
rect 4172 10146 4200 10746
rect 4264 10266 4292 16662
rect 4540 16590 4568 16748
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4540 16114 4568 16526
rect 4724 16232 4752 22630
rect 4908 19009 4936 24550
rect 5092 24342 5120 24754
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5080 24336 5132 24342
rect 5080 24278 5132 24284
rect 5092 23798 5120 24278
rect 5184 23905 5212 24550
rect 5170 23896 5226 23905
rect 5170 23831 5226 23840
rect 5080 23792 5132 23798
rect 5078 23760 5080 23769
rect 5132 23760 5134 23769
rect 5276 23730 5304 27390
rect 5368 24585 5396 27520
rect 6012 25242 6040 27520
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 5552 25226 5672 25242
rect 5552 25220 5684 25226
rect 5552 25214 5632 25220
rect 5552 24818 5580 25214
rect 6012 25214 6132 25242
rect 5632 25162 5684 25168
rect 6000 25152 6052 25158
rect 6000 25094 6052 25100
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 6012 24750 6040 25094
rect 6104 24857 6132 25214
rect 6090 24848 6146 24857
rect 6090 24783 6146 24792
rect 6000 24744 6052 24750
rect 5538 24712 5594 24721
rect 6000 24686 6052 24692
rect 5538 24647 5594 24656
rect 5354 24576 5410 24585
rect 5354 24511 5410 24520
rect 5354 24168 5410 24177
rect 5354 24103 5410 24112
rect 5368 23866 5396 24103
rect 5552 23866 5580 24647
rect 6000 24608 6052 24614
rect 6196 24596 6224 25434
rect 6052 24568 6224 24596
rect 6000 24550 6052 24556
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5356 23860 5408 23866
rect 5356 23802 5408 23808
rect 5540 23860 5592 23866
rect 5540 23802 5592 23808
rect 5078 23695 5134 23704
rect 5264 23724 5316 23730
rect 5264 23666 5316 23672
rect 5368 23662 5396 23802
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5170 22672 5226 22681
rect 5276 22642 5304 23423
rect 5354 23352 5410 23361
rect 5354 23287 5410 23296
rect 5170 22607 5226 22616
rect 5264 22636 5316 22642
rect 5184 22574 5212 22607
rect 5264 22578 5316 22584
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 5368 20398 5396 23287
rect 6012 23225 6040 24550
rect 6274 24440 6330 24449
rect 6274 24375 6330 24384
rect 5998 23216 6054 23225
rect 5998 23151 6054 23160
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 22642 5488 22918
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 5460 21690 5488 22578
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5998 21856 6054 21865
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5552 21457 5580 21830
rect 5622 21788 5918 21808
rect 5998 21791 6054 21800
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6012 21690 6040 21791
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5724 21480 5776 21486
rect 5538 21448 5594 21457
rect 5724 21422 5776 21428
rect 5538 21383 5594 21392
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 21185 5488 21286
rect 5446 21176 5502 21185
rect 5736 21146 5764 21422
rect 5446 21111 5502 21120
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5448 20800 5500 20806
rect 5448 20742 5500 20748
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 5460 20466 5488 20742
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5000 20058 5028 20198
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 5000 19378 5028 19994
rect 5092 19825 5120 20198
rect 5460 19990 5488 20402
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5172 19848 5224 19854
rect 5078 19816 5134 19825
rect 5172 19790 5224 19796
rect 5078 19751 5080 19760
rect 5132 19751 5134 19760
rect 5080 19722 5132 19728
rect 5092 19691 5120 19722
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4986 19272 5042 19281
rect 4986 19207 4988 19216
rect 5040 19207 5042 19216
rect 4988 19178 5040 19184
rect 4894 19000 4950 19009
rect 5000 18970 5028 19178
rect 4894 18935 4950 18944
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5184 18698 5212 19790
rect 5276 19514 5304 19926
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5264 19508 5316 19514
rect 5552 19496 5580 19654
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5552 19468 5672 19496
rect 5264 19450 5316 19456
rect 5264 19372 5316 19378
rect 5644 19360 5672 19468
rect 5264 19314 5316 19320
rect 5460 19332 5672 19360
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5184 18222 5212 18634
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5000 17134 5028 17682
rect 5078 17504 5134 17513
rect 5078 17439 5134 17448
rect 4988 17128 5040 17134
rect 4908 17088 4988 17116
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4632 16204 4752 16232
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4632 14770 4660 16204
rect 4816 16182 4844 16662
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4356 14742 4660 14770
rect 4356 12753 4384 14742
rect 4434 14648 4490 14657
rect 4434 14583 4436 14592
rect 4488 14583 4490 14592
rect 4436 14554 4488 14560
rect 4448 14074 4476 14554
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 14074 4660 14350
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4434 13832 4490 13841
rect 4434 13767 4490 13776
rect 4342 12744 4398 12753
rect 4342 12679 4398 12688
rect 4448 12424 4476 13767
rect 4356 12396 4476 12424
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 3976 10134 4028 10140
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9722 3924 9862
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9654 4016 10134
rect 4080 10118 4200 10146
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3792 9172 3844 9178
rect 3712 9132 3792 9160
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3620 7954 3648 8434
rect 3712 8430 3740 9132
rect 3792 9114 3844 9120
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3344 6854 3464 6882
rect 2962 6216 3018 6225
rect 2962 6151 3018 6160
rect 2594 2680 2650 2689
rect 2594 2615 2650 2624
rect 2976 377 3004 6151
rect 3344 3369 3372 6854
rect 3422 6760 3478 6769
rect 3422 6695 3478 6704
rect 3330 3360 3386 3369
rect 3330 3295 3386 3304
rect 3436 1465 3464 6695
rect 3896 3913 3924 9318
rect 3988 7886 4016 9454
rect 4080 9178 4108 10118
rect 4356 9761 4384 12396
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4448 11558 4476 12242
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 4342 9752 4398 9761
rect 4342 9687 4398 9696
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4356 9110 4384 9454
rect 4448 9382 4476 11494
rect 4724 10033 4752 16050
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14006 4844 14826
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12889 4844 13262
rect 4908 12986 4936 17088
rect 4988 17070 5040 17076
rect 5092 17066 5120 17439
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5092 16726 5120 17002
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16794 5212 16934
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5080 16720 5132 16726
rect 5000 16680 5080 16708
rect 5000 14804 5028 16680
rect 5080 16662 5132 16668
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 16250 5212 16526
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5092 15706 5120 16186
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 5092 14958 5120 15642
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5000 14776 5120 14804
rect 4986 14512 5042 14521
rect 4986 14447 5042 14456
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4802 12880 4858 12889
rect 4802 12815 4858 12824
rect 4816 12782 4844 12815
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4908 12714 4936 12922
rect 5000 12782 5028 14447
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4896 11824 4948 11830
rect 4894 11792 4896 11801
rect 4948 11792 4950 11801
rect 4894 11727 4950 11736
rect 5000 10266 5028 12718
rect 5092 11830 5120 14776
rect 5276 14498 5304 19314
rect 5460 18834 5488 19332
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6012 18290 6040 18838
rect 6104 18834 6132 20742
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18284 6052 18290
rect 6000 18226 6052 18232
rect 5540 17808 5592 17814
rect 5540 17750 5592 17756
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 16726 5396 17478
rect 5552 17134 5580 17750
rect 6012 17678 6040 18226
rect 6104 17746 6132 18770
rect 6288 17882 6316 24375
rect 6564 23361 6592 27520
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 6656 24818 6684 25434
rect 6920 25356 6972 25362
rect 6920 25298 6972 25304
rect 6644 24812 6696 24818
rect 6644 24754 6696 24760
rect 6932 24750 6960 25298
rect 6920 24744 6972 24750
rect 6972 24692 7052 24698
rect 6920 24686 7052 24692
rect 6932 24670 7052 24686
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 6550 23352 6606 23361
rect 6550 23287 6606 23296
rect 6840 23089 6868 24550
rect 6932 24070 6960 24550
rect 7024 24449 7052 24670
rect 7010 24440 7066 24449
rect 7010 24375 7066 24384
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23225 6960 24006
rect 7024 23662 7052 24142
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 7024 23322 7052 23598
rect 7116 23497 7144 27520
rect 7380 26852 7432 26858
rect 7380 26794 7432 26800
rect 7392 25226 7420 26794
rect 7668 25362 7696 27520
rect 8220 25498 8248 27520
rect 8484 25764 8536 25770
rect 8484 25706 8536 25712
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 8496 25362 8524 25706
rect 7656 25356 7708 25362
rect 7656 25298 7708 25304
rect 8484 25356 8536 25362
rect 8484 25298 8536 25304
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7300 24818 7328 25162
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7102 23488 7158 23497
rect 7102 23423 7158 23432
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6918 23216 6974 23225
rect 6918 23151 6974 23160
rect 6826 23080 6882 23089
rect 6826 23015 6882 23024
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6380 22234 6408 22714
rect 6656 22574 6684 22918
rect 7024 22778 7052 23258
rect 7300 22778 7328 24754
rect 7484 24342 7512 24754
rect 7576 24614 7604 25230
rect 8208 24676 8260 24682
rect 8260 24636 8340 24664
rect 8208 24618 8260 24624
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7472 24336 7524 24342
rect 7472 24278 7524 24284
rect 7484 23866 7512 24278
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7746 23488 7802 23497
rect 7746 23423 7802 23432
rect 7380 23180 7432 23186
rect 7380 23122 7432 23128
rect 7012 22772 7064 22778
rect 7012 22714 7064 22720
rect 7288 22772 7340 22778
rect 7288 22714 7340 22720
rect 7392 22642 7420 23122
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7760 22574 7788 23423
rect 8022 23352 8078 23361
rect 8312 23322 8340 24636
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8404 24070 8432 24550
rect 8496 24410 8524 25298
rect 8668 24744 8720 24750
rect 8668 24686 8720 24692
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8680 24070 8708 24686
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8404 23594 8432 24006
rect 8484 23792 8536 23798
rect 8482 23760 8484 23769
rect 8536 23760 8538 23769
rect 8482 23695 8538 23704
rect 8680 23633 8708 24006
rect 8666 23624 8722 23633
rect 8392 23588 8444 23594
rect 8666 23559 8722 23568
rect 8392 23530 8444 23536
rect 8864 23497 8892 27520
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9324 23526 9352 24210
rect 9312 23520 9364 23526
rect 8850 23488 8906 23497
rect 9312 23462 9364 23468
rect 8850 23423 8906 23432
rect 8022 23287 8078 23296
rect 8300 23316 8352 23322
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 7748 22568 7800 22574
rect 7748 22510 7800 22516
rect 6368 22228 6420 22234
rect 6368 22170 6420 22176
rect 6380 21010 6408 22170
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6472 21350 6500 22034
rect 6460 21344 6512 21350
rect 6458 21312 6460 21321
rect 6512 21312 6514 21321
rect 6458 21247 6514 21256
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6656 19786 6684 22510
rect 6920 22024 6972 22030
rect 6920 21966 6972 21972
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6932 21146 6960 21966
rect 7024 21350 7052 21966
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7668 21486 7696 21830
rect 8036 21554 8064 23287
rect 8300 23258 8352 23264
rect 9324 22681 9352 23462
rect 9416 23361 9444 27520
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9692 24954 9720 25298
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 9692 24857 9720 24890
rect 9678 24848 9734 24857
rect 9678 24783 9734 24792
rect 9588 24676 9640 24682
rect 9588 24618 9640 24624
rect 9402 23352 9458 23361
rect 9402 23287 9458 23296
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9310 22672 9366 22681
rect 8116 22636 8168 22642
rect 9508 22642 9536 22918
rect 9310 22607 9366 22616
rect 9496 22636 9548 22642
rect 8116 22578 8168 22584
rect 9496 22578 9548 22584
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7656 21480 7708 21486
rect 7656 21422 7708 21428
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 7564 21344 7616 21350
rect 7564 21286 7616 21292
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 7024 21010 7052 21286
rect 7576 21146 7604 21286
rect 7564 21140 7616 21146
rect 7564 21082 7616 21088
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 6840 20466 6868 20946
rect 7024 20602 7052 20946
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6932 20058 6960 20334
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 6564 19446 6592 19654
rect 6552 19440 6604 19446
rect 6552 19382 6604 19388
rect 7300 19378 7328 19654
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 6920 19236 6972 19242
rect 6920 19178 6972 19184
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6472 18970 6500 19110
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6368 18148 6420 18154
rect 6368 18090 6420 18096
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6092 17740 6144 17746
rect 6092 17682 6144 17688
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5906 17232 5962 17241
rect 5632 17196 5684 17202
rect 6012 17202 6040 17614
rect 6288 17338 6316 17818
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 5906 17167 5962 17176
rect 6000 17196 6052 17202
rect 5632 17138 5684 17144
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5644 16658 5672 17138
rect 5920 16658 5948 17167
rect 6000 17138 6052 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5998 16280 6054 16289
rect 5998 16215 6000 16224
rect 6052 16215 6054 16224
rect 6000 16186 6052 16192
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5828 15570 5856 15982
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 6000 15564 6052 15570
rect 6000 15506 6052 15512
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5276 14470 5396 14498
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5276 14006 5304 14214
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5172 13728 5224 13734
rect 5172 13670 5224 13676
rect 5184 13530 5212 13670
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5170 13288 5226 13297
rect 5170 13223 5226 13232
rect 5184 12986 5212 13223
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5276 12782 5304 13466
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5368 12322 5396 14470
rect 5460 13938 5488 15302
rect 5552 15162 5580 15506
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 6012 14822 6040 15506
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 14521 5764 14554
rect 5722 14512 5778 14521
rect 5722 14447 5778 14456
rect 5828 14414 5856 14758
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 12442 5488 13874
rect 5552 13530 5580 14010
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 13530 5764 13738
rect 6000 13728 6052 13734
rect 6000 13670 6052 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12832 5580 13126
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5724 12844 5776 12850
rect 5552 12804 5724 12832
rect 5724 12786 5776 12792
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5368 12294 5488 12322
rect 5736 12306 5764 12786
rect 5906 12336 5962 12345
rect 5170 12200 5226 12209
rect 5170 12135 5226 12144
rect 5184 11898 5212 12135
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 11824 5132 11830
rect 5080 11766 5132 11772
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5276 11354 5304 11630
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5170 10432 5226 10441
rect 5170 10367 5226 10376
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5080 10056 5132 10062
rect 4526 10024 4582 10033
rect 4526 9959 4582 9968
rect 4710 10024 4766 10033
rect 5080 9998 5132 10004
rect 4710 9959 4766 9968
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4540 8634 4568 9959
rect 5092 9654 5120 9998
rect 5184 9926 5212 10367
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 5184 9466 5212 9862
rect 5092 9438 5212 9466
rect 5092 9042 5120 9438
rect 5276 9178 5304 11290
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4540 8430 4568 8570
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 5092 8090 5120 8978
rect 5276 8430 5304 9114
rect 5368 9110 5396 10406
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8498 5396 9046
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5264 8424 5316 8430
rect 5264 8366 5316 8372
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4066 7848 4122 7857
rect 4066 7783 4068 7792
rect 4120 7783 4122 7792
rect 4068 7754 4120 7760
rect 4172 7546 4200 7958
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7546 4568 7822
rect 4632 7750 4660 8026
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4632 7478 4660 7686
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 3882 3904 3938 3913
rect 3882 3839 3938 3848
rect 5460 3505 5488 12294
rect 5724 12300 5776 12306
rect 5906 12271 5962 12280
rect 5724 12242 5776 12248
rect 5920 12238 5948 12271
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 6012 11762 6040 13670
rect 6104 13410 6132 17070
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6288 16250 6316 16526
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6380 15688 6408 18090
rect 6472 16114 6500 18906
rect 6840 18465 6868 19110
rect 6932 18630 6960 19178
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 18970 7236 19110
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6552 18080 6604 18086
rect 6550 18048 6552 18057
rect 6604 18048 6606 18057
rect 6550 17983 6606 17992
rect 6932 17814 6960 18566
rect 7300 18426 7328 19314
rect 7576 18970 7604 19858
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7668 18737 7696 21422
rect 8128 21146 8156 22578
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8220 21554 8248 21830
rect 8312 21729 8340 22442
rect 9404 22432 9456 22438
rect 8482 22400 8538 22409
rect 9404 22374 9456 22380
rect 8482 22335 8538 22344
rect 8392 22092 8444 22098
rect 8392 22034 8444 22040
rect 8298 21720 8354 21729
rect 8298 21655 8354 21664
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8022 20904 8078 20913
rect 8022 20839 8078 20848
rect 8036 20058 8064 20839
rect 8220 20641 8248 21490
rect 8404 21146 8432 22034
rect 8496 22030 8524 22335
rect 9416 22137 9444 22374
rect 9402 22128 9458 22137
rect 9600 22098 9628 24618
rect 9968 24426 9996 27520
rect 10520 25786 10548 27520
rect 11072 27418 11100 27520
rect 11072 27390 11284 27418
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 10520 25758 10824 25786
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10060 24585 10088 25298
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 10046 24576 10102 24585
rect 10046 24511 10102 24520
rect 9876 24398 9996 24426
rect 9876 24313 9904 24398
rect 9956 24336 10008 24342
rect 9862 24304 9918 24313
rect 9956 24278 10008 24284
rect 9862 24239 9918 24248
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9678 22672 9734 22681
rect 9678 22607 9734 22616
rect 9402 22063 9458 22072
rect 9588 22092 9640 22098
rect 9588 22034 9640 22040
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 9310 21448 9366 21457
rect 9310 21383 9366 21392
rect 8852 21344 8904 21350
rect 8852 21286 8904 21292
rect 8392 21140 8444 21146
rect 8392 21082 8444 21088
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8206 20632 8262 20641
rect 8588 20602 8616 20946
rect 8206 20567 8262 20576
rect 8576 20596 8628 20602
rect 8220 20398 8248 20567
rect 8576 20538 8628 20544
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8390 20088 8446 20097
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8208 20052 8260 20058
rect 8390 20023 8446 20032
rect 8208 19994 8260 20000
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 7944 19446 7972 19654
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 8220 18970 8248 19994
rect 8404 19922 8432 20023
rect 8588 19990 8616 20538
rect 8864 20058 8892 21286
rect 9324 21146 9352 21383
rect 9416 21350 9444 21830
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9692 21162 9720 22607
rect 9876 22574 9904 24006
rect 9968 23866 9996 24278
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 10060 23662 10088 24074
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9956 23180 10008 23186
rect 10060 23168 10088 23598
rect 10152 23254 10180 24822
rect 10230 24712 10286 24721
rect 10230 24647 10232 24656
rect 10284 24647 10286 24656
rect 10232 24618 10284 24624
rect 10704 24614 10732 25094
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10704 24410 10732 24550
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10008 23140 10088 23168
rect 9956 23122 10008 23128
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9864 22568 9916 22574
rect 9864 22510 9916 22516
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22137 9812 22374
rect 9770 22128 9826 22137
rect 9770 22063 9826 22072
rect 9968 21894 9996 22578
rect 10060 22166 10088 23140
rect 10152 22778 10180 23190
rect 10140 22772 10192 22778
rect 10140 22714 10192 22720
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9312 21140 9364 21146
rect 9692 21134 9904 21162
rect 9312 21082 9364 21088
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 20398 9628 20742
rect 9692 20602 9720 21014
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 9324 20058 9352 20266
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8404 19378 8432 19858
rect 8588 19514 8616 19926
rect 9324 19854 9352 19994
rect 9692 19854 9720 20198
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9324 19514 9352 19790
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 9416 19310 9444 19654
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8390 18864 8446 18873
rect 7932 18828 7984 18834
rect 9048 18834 9076 19110
rect 8390 18799 8446 18808
rect 9036 18828 9088 18834
rect 7932 18770 7984 18776
rect 7654 18728 7710 18737
rect 7654 18663 7710 18672
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7392 18290 7420 18566
rect 7944 18426 7972 18770
rect 8404 18426 8432 18799
rect 9036 18770 9088 18776
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8312 18086 8340 18226
rect 8390 18184 8446 18193
rect 8390 18119 8446 18128
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6564 16794 6592 16934
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6380 15660 6500 15688
rect 6472 14482 6500 15660
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 14278 6408 14350
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6196 13870 6224 14214
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6182 13696 6238 13705
rect 6182 13631 6238 13640
rect 6196 13530 6224 13631
rect 6184 13524 6236 13530
rect 6236 13484 6316 13512
rect 6184 13466 6236 13472
rect 6104 13382 6224 13410
rect 6196 12866 6224 13382
rect 6288 12918 6316 13484
rect 6380 13326 6408 14214
rect 6472 14006 6500 14418
rect 6656 14414 6684 17274
rect 6840 17270 6868 17478
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6932 16998 6960 17750
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 6920 16992 6972 16998
rect 6840 16952 6920 16980
rect 6840 16590 6868 16952
rect 6920 16934 6972 16940
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 7024 16046 7052 17206
rect 7668 17105 7696 17682
rect 8312 17542 8340 18022
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 7654 17096 7710 17105
rect 7654 17031 7710 17040
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6656 14074 6684 14350
rect 6748 14278 6776 14350
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6840 14113 6868 14894
rect 6826 14104 6882 14113
rect 6644 14068 6696 14074
rect 6696 14028 6776 14056
rect 6826 14039 6882 14048
rect 6644 14010 6696 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6104 12838 6224 12866
rect 6276 12912 6328 12918
rect 6276 12854 6328 12860
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6104 11694 6132 12838
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 12424 6224 12718
rect 6380 12442 6408 13262
rect 6368 12436 6420 12442
rect 6196 12396 6316 12424
rect 6288 12345 6316 12396
rect 6368 12378 6420 12384
rect 6472 12374 6500 13942
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6564 12986 6592 13330
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6460 12368 6512 12374
rect 6274 12336 6330 12345
rect 6564 12345 6592 12922
rect 6460 12310 6512 12316
rect 6550 12336 6606 12345
rect 6274 12271 6330 12280
rect 6288 11914 6316 12271
rect 6288 11886 6408 11914
rect 6472 11898 6500 12310
rect 6550 12271 6606 12280
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10470 5580 11154
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 6012 10538 6040 11018
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 8090 5580 10406
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 6012 8634 6040 10474
rect 6196 10470 6224 11086
rect 6380 11082 6408 11886
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6656 11694 6684 12242
rect 6748 11898 6776 14028
rect 6828 14000 6880 14006
rect 6826 13968 6828 13977
rect 6880 13968 6882 13977
rect 6826 13903 6882 13912
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6932 13530 6960 13874
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6932 13190 6960 13466
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6932 12782 6960 13126
rect 7024 12889 7052 15846
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7010 12880 7066 12889
rect 7010 12815 7066 12824
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6932 12442 6960 12718
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7116 12288 7144 14554
rect 7300 13462 7328 16526
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 14890 7420 15302
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7392 14278 7420 14826
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13938 7420 14214
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 6840 12260 7144 12288
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6840 11354 6868 12260
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10198 6224 10406
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6196 9382 6224 10134
rect 6380 9926 6408 11018
rect 6656 10169 6684 11290
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7116 10810 7144 11086
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6642 10160 6698 10169
rect 6642 10095 6698 10104
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9722 6408 9862
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6380 9110 6408 9658
rect 7116 9178 7144 10746
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9450 7420 9862
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 7392 8906 7420 9386
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 7484 4146 7512 16934
rect 7668 16658 7696 17031
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7748 16652 7800 16658
rect 7852 16640 7880 17478
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7800 16612 7880 16640
rect 7748 16594 7800 16600
rect 7760 15706 7788 16594
rect 8220 15706 8248 17274
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8312 16250 8340 16662
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8220 14482 8248 15642
rect 8312 15162 8340 16186
rect 8404 15910 8432 18119
rect 8496 17785 8524 18702
rect 8758 18456 8814 18465
rect 8758 18391 8814 18400
rect 8772 18222 8800 18391
rect 8760 18216 8812 18222
rect 8666 18184 8722 18193
rect 8760 18158 8812 18164
rect 8666 18119 8668 18128
rect 8720 18119 8722 18128
rect 8668 18090 8720 18096
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8482 17776 8538 17785
rect 8482 17711 8538 17720
rect 8588 17542 8616 18022
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 8588 17241 8616 17478
rect 9140 17270 9168 17478
rect 9232 17338 9260 19246
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9402 18728 9458 18737
rect 9402 18663 9458 18672
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9128 17264 9180 17270
rect 8574 17232 8630 17241
rect 9180 17212 9260 17218
rect 9128 17206 9260 17212
rect 8574 17167 8630 17176
rect 9140 17190 9260 17206
rect 9140 17141 9168 17190
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 16289 9076 16390
rect 9034 16280 9090 16289
rect 9034 16215 9090 16224
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8390 15328 8446 15337
rect 8390 15263 8446 15272
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8404 14482 8432 15263
rect 8496 14929 8524 15438
rect 8588 15094 8616 15506
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 9140 14958 9168 15302
rect 9128 14952 9180 14958
rect 8482 14920 8538 14929
rect 9128 14894 9180 14900
rect 8482 14855 8538 14864
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8404 14362 8432 14418
rect 8312 14334 8432 14362
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8312 14074 8340 14334
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7748 13320 7800 13326
rect 7746 13288 7748 13297
rect 7800 13288 7802 13297
rect 7746 13223 7802 13232
rect 7760 12714 7788 13223
rect 7748 12708 7800 12714
rect 7748 12650 7800 12656
rect 7838 11112 7894 11121
rect 7838 11047 7840 11056
rect 7892 11047 7894 11056
rect 7840 11018 7892 11024
rect 7746 10024 7802 10033
rect 7746 9959 7802 9968
rect 7654 9344 7710 9353
rect 7654 9279 7710 9288
rect 7668 9110 7696 9279
rect 7760 9178 7788 9959
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7656 9104 7708 9110
rect 7656 9046 7708 9052
rect 7668 8566 7696 9046
rect 7760 8634 7788 9114
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7944 6769 7972 14010
rect 8404 13870 8432 14214
rect 8208 13864 8260 13870
rect 8392 13864 8444 13870
rect 8260 13812 8340 13818
rect 8208 13806 8340 13812
rect 8392 13806 8444 13812
rect 8220 13790 8340 13806
rect 8312 13462 8340 13790
rect 8496 13530 8524 14350
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8300 13456 8352 13462
rect 8300 13398 8352 13404
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8128 12209 8156 13330
rect 8496 12986 8524 13466
rect 8588 13394 8616 14350
rect 8956 13870 8984 14486
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9048 14113 9076 14350
rect 9232 14249 9260 17190
rect 9310 16552 9366 16561
rect 9310 16487 9366 16496
rect 9324 16114 9352 16487
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9218 14240 9274 14249
rect 9218 14175 9274 14184
rect 9034 14104 9090 14113
rect 9034 14039 9090 14048
rect 9048 13938 9076 14039
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8208 12912 8260 12918
rect 8206 12880 8208 12889
rect 8260 12880 8262 12889
rect 8206 12815 8262 12824
rect 8852 12776 8904 12782
rect 8850 12744 8852 12753
rect 8904 12744 8906 12753
rect 8850 12679 8906 12688
rect 8956 12442 8984 13806
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8300 12368 8352 12374
rect 8298 12336 8300 12345
rect 8352 12336 8354 12345
rect 8298 12271 8354 12280
rect 8114 12200 8170 12209
rect 8114 12135 8116 12144
rect 8168 12135 8170 12144
rect 8298 12200 8354 12209
rect 8298 12135 8354 12144
rect 8116 12106 8168 12112
rect 8312 11694 8340 12135
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8576 11756 8628 11762
rect 8852 11756 8904 11762
rect 8628 11716 8852 11744
rect 8576 11698 8628 11704
rect 8852 11698 8904 11704
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8864 11286 8892 11698
rect 8852 11280 8904 11286
rect 8852 11222 8904 11228
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8220 10810 8248 11154
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8496 10606 8524 10950
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 10266 8524 10542
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8496 9722 8524 10202
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8634 8064 8910
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7930 6760 7986 6769
rect 7930 6695 7986 6704
rect 9048 6225 9076 12038
rect 9232 11898 9260 14175
rect 9416 12714 9444 18663
rect 9508 18630 9536 19110
rect 9600 18970 9628 19314
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9692 18766 9720 19790
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 19145 9812 19246
rect 9770 19136 9826 19145
rect 9770 19071 9826 19080
rect 9770 19000 9826 19009
rect 9770 18935 9826 18944
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9508 18426 9536 18566
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9784 18358 9812 18935
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9588 16040 9640 16046
rect 9692 16028 9720 17546
rect 9784 16794 9812 17614
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9876 16590 9904 21134
rect 9968 21078 9996 21830
rect 10520 21690 10548 22034
rect 10796 22001 10824 25758
rect 11164 25498 11192 26318
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10888 24954 10916 25298
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 11256 24834 11284 27390
rect 11164 24806 11284 24834
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10888 23254 10916 23462
rect 10980 23322 11008 24142
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10876 23248 10928 23254
rect 10876 23190 10928 23196
rect 10980 22098 11008 23258
rect 10968 22092 11020 22098
rect 10968 22034 11020 22040
rect 10782 21992 10838 22001
rect 10782 21927 10838 21936
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10138 21448 10194 21457
rect 10138 21383 10194 21392
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9968 18902 9996 19926
rect 10060 19825 10088 21286
rect 10046 19816 10102 19825
rect 10046 19751 10102 19760
rect 10060 19174 10088 19751
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 10060 18834 10088 19110
rect 10152 18902 10180 21383
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10796 21146 10824 21490
rect 10968 21480 11020 21486
rect 11164 21468 11192 24806
rect 11716 24342 11744 27520
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 11704 24336 11756 24342
rect 11704 24278 11756 24284
rect 11978 24304 12034 24313
rect 11888 24268 11940 24274
rect 11978 24239 11980 24248
rect 11888 24210 11940 24216
rect 12032 24239 12034 24248
rect 11980 24210 12032 24216
rect 11900 23322 11928 24210
rect 11992 23798 12020 24210
rect 11980 23792 12032 23798
rect 11980 23734 12032 23740
rect 11428 23316 11480 23322
rect 11428 23258 11480 23264
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11020 21440 11192 21468
rect 11256 21457 11284 22034
rect 11348 21865 11376 22442
rect 11334 21856 11390 21865
rect 11334 21791 11390 21800
rect 11242 21448 11298 21457
rect 10968 21422 11020 21428
rect 11242 21383 11298 21392
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10414 20632 10470 20641
rect 10414 20567 10416 20576
rect 10468 20567 10470 20576
rect 10416 20538 10468 20544
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10796 19990 10824 21082
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10244 19242 10548 19258
rect 10232 19236 10548 19242
rect 10284 19230 10548 19236
rect 10520 19224 10548 19230
rect 10692 19236 10744 19242
rect 10520 19196 10692 19224
rect 10232 19178 10284 19184
rect 10692 19178 10744 19184
rect 10980 19174 11008 20266
rect 11072 19961 11100 21286
rect 11152 20800 11204 20806
rect 11152 20742 11204 20748
rect 11164 20602 11192 20742
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11164 20058 11192 20538
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11348 19990 11376 20198
rect 11336 19984 11388 19990
rect 11058 19952 11114 19961
rect 11336 19926 11388 19932
rect 11058 19887 11114 19896
rect 11348 19718 11376 19926
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10152 18222 10180 18838
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10428 18154 10456 18702
rect 10980 18601 11008 19110
rect 11164 18834 11192 19246
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18902 11376 19110
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 10966 18592 11022 18601
rect 10966 18527 11022 18536
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 11072 18086 11100 18294
rect 11164 18290 11192 18770
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 16794 9996 17682
rect 10060 17202 10088 18022
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 11072 17762 11100 18022
rect 11164 17882 11192 18226
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11072 17734 11192 17762
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10152 17134 10180 17478
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9864 16584 9916 16590
rect 9916 16544 9996 16572
rect 9864 16526 9916 16532
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9640 16000 9720 16028
rect 9772 16040 9824 16046
rect 9588 15982 9640 15988
rect 9772 15982 9824 15988
rect 9600 15706 9628 15982
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14929 9628 14962
rect 9680 14952 9732 14958
rect 9586 14920 9642 14929
rect 9680 14894 9732 14900
rect 9586 14855 9642 14864
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9508 14618 9536 14758
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13258 9628 13738
rect 9692 13530 9720 14894
rect 9784 14074 9812 15982
rect 9876 15706 9904 16186
rect 9968 16182 9996 16544
rect 10152 16522 10180 17070
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 9956 16176 10008 16182
rect 9956 16118 10008 16124
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9968 14906 9996 16118
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9876 14878 9996 14906
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9600 12889 9628 13194
rect 9586 12880 9642 12889
rect 9586 12815 9588 12824
rect 9640 12815 9642 12824
rect 9588 12786 9640 12792
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 12102 9444 12650
rect 9784 12306 9812 14010
rect 9876 13462 9904 14878
rect 10060 14278 10088 15846
rect 10152 15706 10180 16458
rect 10336 16250 10364 16594
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10690 16144 10746 16153
rect 11072 16114 11100 16390
rect 10690 16079 10746 16088
rect 11060 16108 11112 16114
rect 10704 16046 10732 16079
rect 11060 16050 11112 16056
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10796 15570 10824 15846
rect 10888 15706 10916 15914
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10704 15162 10732 15438
rect 10980 15162 11008 15982
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11058 14920 11114 14929
rect 11058 14855 11114 14864
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10152 13841 10180 14758
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11072 14618 11100 14855
rect 11164 14822 11192 17734
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11256 16046 11284 16390
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11348 15502 11376 18838
rect 11440 18086 11468 23258
rect 11886 21040 11942 21049
rect 11886 20975 11888 20984
rect 11940 20975 11942 20984
rect 11888 20946 11940 20952
rect 11900 20602 11928 20946
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 19553 11928 19790
rect 11886 19544 11942 19553
rect 11886 19479 11942 19488
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11532 17882 11560 18158
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 17338 11468 17614
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11992 16794 12020 23734
rect 12084 21146 12112 26386
rect 12164 24608 12216 24614
rect 12164 24550 12216 24556
rect 12176 22778 12204 24550
rect 12268 24410 12296 27520
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12360 24818 12388 25230
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12636 24614 12664 24754
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12256 24404 12308 24410
rect 12256 24346 12308 24352
rect 12268 23866 12296 24346
rect 12820 24342 12848 27520
rect 13266 24848 13322 24857
rect 12992 24812 13044 24818
rect 13372 24818 13400 27520
rect 13636 25696 13688 25702
rect 13636 25638 13688 25644
rect 13648 25498 13676 25638
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13266 24783 13322 24792
rect 13360 24812 13412 24818
rect 12992 24754 13044 24760
rect 12808 24336 12860 24342
rect 12808 24278 12860 24284
rect 12348 24200 12400 24206
rect 12346 24168 12348 24177
rect 12400 24168 12402 24177
rect 12346 24103 12402 24112
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12360 23662 12388 24103
rect 12820 23866 12848 24278
rect 12900 24132 12952 24138
rect 12900 24074 12952 24080
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12912 23662 12940 24074
rect 13004 24070 13032 24754
rect 13084 24676 13136 24682
rect 13084 24618 13136 24624
rect 13096 24410 13124 24618
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12360 23322 12388 23598
rect 12348 23316 12400 23322
rect 12348 23258 12400 23264
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12164 22772 12216 22778
rect 12164 22714 12216 22720
rect 12360 22710 12388 23122
rect 12912 22982 12940 23598
rect 13004 23594 13032 24006
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 12900 22976 12952 22982
rect 12952 22924 13032 22930
rect 12900 22918 13032 22924
rect 12912 22902 13032 22918
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 13004 22642 13032 22902
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13004 22030 13032 22578
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12898 21584 12954 21593
rect 12898 21519 12954 21528
rect 12912 21486 12940 21519
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 13004 20942 13032 21966
rect 13096 21842 13124 22374
rect 13176 21888 13228 21894
rect 13096 21836 13176 21842
rect 13096 21830 13228 21836
rect 13096 21814 13216 21830
rect 13096 21554 13124 21814
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 13096 21146 13124 21490
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13084 21004 13136 21010
rect 13084 20946 13136 20952
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13096 20602 13124 20946
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13084 20392 13136 20398
rect 13084 20334 13136 20340
rect 12348 20052 12400 20058
rect 12348 19994 12400 20000
rect 12360 19310 12388 19994
rect 13096 19718 13124 20334
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12452 19310 12480 19654
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12544 18970 12572 19178
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12360 18358 12388 18838
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11992 16250 12020 16730
rect 12084 16590 12112 16730
rect 12162 16688 12218 16697
rect 12162 16623 12218 16632
rect 12176 16590 12204 16623
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11428 15496 11480 15502
rect 11428 15438 11480 15444
rect 11440 15026 11468 15438
rect 11428 15020 11480 15026
rect 11428 14962 11480 14968
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11256 14074 11284 14758
rect 11440 14618 11468 14962
rect 11900 14822 11928 15506
rect 11992 15337 12020 16186
rect 12084 15706 12112 16526
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12452 15502 12480 15982
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 11978 15328 12034 15337
rect 11978 15263 12034 15272
rect 12452 14958 12480 15438
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 11888 14816 11940 14822
rect 11886 14784 11888 14793
rect 11940 14784 11942 14793
rect 11886 14719 11942 14728
rect 11992 14634 12020 14894
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11900 14606 12020 14634
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11704 14272 11756 14278
rect 11702 14240 11704 14249
rect 11756 14240 11758 14249
rect 11702 14175 11758 14184
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11808 14006 11836 14486
rect 11900 14414 11928 14606
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 14278 11928 14350
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 14000 11848 14006
rect 11796 13942 11848 13948
rect 10138 13832 10194 13841
rect 10138 13767 10194 13776
rect 10048 13728 10100 13734
rect 10048 13670 10100 13676
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9876 12986 9904 13398
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9968 12442 9996 13466
rect 10060 13394 10088 13670
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 11256 13530 11284 13670
rect 11900 13530 11928 14214
rect 12544 13802 12572 18294
rect 12728 18222 12756 18566
rect 12820 18358 12848 18906
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12912 18222 12940 19178
rect 13280 18970 13308 24783
rect 13360 24754 13412 24760
rect 13820 24812 13872 24818
rect 13820 24754 13872 24760
rect 13542 24576 13598 24585
rect 13542 24511 13598 24520
rect 13450 21720 13506 21729
rect 13450 21655 13452 21664
rect 13504 21655 13506 21664
rect 13452 21626 13504 21632
rect 13464 21486 13492 21626
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 20482 13492 21422
rect 13372 20454 13492 20482
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13372 18902 13400 20454
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13464 19854 13492 20266
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13464 19514 13492 19790
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13360 18896 13412 18902
rect 13360 18838 13412 18844
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 17542 12940 18158
rect 13280 18154 13308 18702
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13280 17882 13308 18090
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 13096 17338 13124 17682
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12714 17096 12770 17105
rect 12714 17031 12770 17040
rect 12728 16998 12756 17031
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12728 16726 12756 16934
rect 13556 16794 13584 24511
rect 13728 23588 13780 23594
rect 13728 23530 13780 23536
rect 13740 23322 13768 23530
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13832 21690 13860 24754
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13728 20052 13780 20058
rect 13924 20040 13952 27520
rect 14568 24857 14596 27520
rect 15120 25242 15148 27520
rect 15672 27418 15700 27520
rect 14844 25214 15148 25242
rect 15488 27390 15700 27418
rect 14554 24848 14610 24857
rect 14554 24783 14610 24792
rect 14002 24712 14058 24721
rect 14002 24647 14004 24656
rect 14056 24647 14058 24656
rect 14004 24618 14056 24624
rect 14844 24585 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 14830 24576 14886 24585
rect 14830 24511 14886 24520
rect 14556 24200 14608 24206
rect 14278 24168 14334 24177
rect 14556 24142 14608 24148
rect 14278 24103 14334 24112
rect 14292 23866 14320 24103
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 13780 20012 13952 20040
rect 13728 19994 13780 20000
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13648 19174 13676 19858
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13648 18737 13676 19110
rect 13832 18970 13860 19450
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13634 18728 13690 18737
rect 13634 18663 13690 18672
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16153 12664 16594
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 13096 15978 13124 16390
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 13556 15910 13584 16730
rect 13648 16658 13676 18663
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13740 17882 13768 18158
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 14004 17672 14056 17678
rect 14002 17640 14004 17649
rect 14056 17640 14058 17649
rect 14002 17575 14058 17584
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13648 16046 13676 16594
rect 13740 16590 13768 16934
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 16250 13768 16526
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 16040 13688 16046
rect 13636 15982 13688 15988
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13832 15706 13860 15914
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 15162 13860 15506
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14200 15162 14228 15302
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13280 14618 13308 14826
rect 14094 14784 14150 14793
rect 14094 14719 14150 14728
rect 14108 14618 14136 14719
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 12898 14376 12954 14385
rect 12898 14311 12954 14320
rect 12912 13938 12940 14311
rect 13280 13938 13308 14554
rect 14200 14550 14228 15098
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 13556 14278 13584 14486
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 14074 13584 14214
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 14384 13938 14412 23598
rect 14568 23526 14596 24142
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14556 23520 14608 23526
rect 14556 23462 14608 23468
rect 14568 22778 14596 23462
rect 15382 23216 15438 23225
rect 15292 23180 15344 23186
rect 15382 23151 15438 23160
rect 15292 23122 15344 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22778 15332 23122
rect 14556 22772 14608 22778
rect 14556 22714 14608 22720
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15396 22642 15424 23151
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14648 22092 14700 22098
rect 14648 22034 14700 22040
rect 14660 21554 14688 22034
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 21146 14688 21490
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14752 20806 14780 22374
rect 15292 22160 15344 22166
rect 15292 22102 15344 22108
rect 15382 22128 15438 22137
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21593 15332 22102
rect 15382 22063 15438 22072
rect 15290 21584 15346 21593
rect 15396 21554 15424 22063
rect 15290 21519 15346 21528
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14752 20602 14780 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14462 19544 14518 19553
rect 14462 19479 14518 19488
rect 14476 19310 14504 19479
rect 14568 19446 14596 20538
rect 15198 20496 15254 20505
rect 15198 20431 15254 20440
rect 15212 19922 15240 20431
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14568 18970 14596 19382
rect 14660 19378 14688 19722
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 15304 19281 15332 20198
rect 15290 19272 15346 19281
rect 15290 19207 15346 19216
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 14568 17882 14596 18022
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14568 17134 14596 17818
rect 14660 17746 14688 19110
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14648 17740 14700 17746
rect 14648 17682 14700 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14568 16794 14596 17070
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14936 16697 14964 16934
rect 15212 16794 15240 16934
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 14922 16688 14978 16697
rect 14922 16623 14978 16632
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 16046 15332 16594
rect 15488 16130 15516 27390
rect 16028 24268 16080 24274
rect 16028 24210 16080 24216
rect 16120 24268 16172 24274
rect 16120 24210 16172 24216
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15580 23254 15608 23598
rect 16040 23526 16068 24210
rect 16132 23526 16160 24210
rect 16224 23866 16252 27520
rect 16488 24404 16540 24410
rect 16776 24392 16804 27520
rect 16540 24364 16804 24392
rect 16488 24346 16540 24352
rect 17420 23905 17448 27520
rect 17682 24440 17738 24449
rect 17682 24375 17738 24384
rect 17868 24404 17920 24410
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 16394 23896 16450 23905
rect 16212 23860 16264 23866
rect 16394 23831 16396 23840
rect 16212 23802 16264 23808
rect 16448 23831 16450 23840
rect 17406 23896 17462 23905
rect 17406 23831 17462 23840
rect 16396 23802 16448 23808
rect 16408 23594 16620 23610
rect 17512 23594 17540 24210
rect 17696 24138 17724 24375
rect 17972 24392 18000 27520
rect 17920 24364 18000 24392
rect 17868 24346 17920 24352
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 16408 23588 16632 23594
rect 16408 23582 16580 23588
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 16120 23520 16172 23526
rect 16120 23462 16172 23468
rect 15568 23248 15620 23254
rect 15568 23190 15620 23196
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15672 19514 15700 19858
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15764 18873 15792 22714
rect 16040 19990 16068 23462
rect 16028 19984 16080 19990
rect 16028 19926 16080 19932
rect 15750 18864 15806 18873
rect 15750 18799 15806 18808
rect 16132 16726 16160 23462
rect 16302 22536 16358 22545
rect 16302 22471 16358 22480
rect 16316 22234 16344 22471
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16408 22114 16436 23582
rect 16580 23530 16632 23536
rect 17500 23588 17552 23594
rect 17500 23530 17552 23536
rect 17592 23588 17644 23594
rect 17592 23530 17644 23536
rect 16762 23488 16818 23497
rect 16762 23423 16818 23432
rect 16776 23322 16804 23423
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16592 22438 16620 23122
rect 16580 22432 16632 22438
rect 16580 22374 16632 22380
rect 16316 22086 16436 22114
rect 16120 16720 16172 16726
rect 16120 16662 16172 16668
rect 15396 16102 15516 16130
rect 15292 16040 15344 16046
rect 15290 16008 15292 16017
rect 15344 16008 15346 16017
rect 15290 15943 15346 15952
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15396 14385 15424 16102
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15382 14376 15438 14385
rect 15382 14311 15438 14320
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14554 13968 14610 13977
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 14372 13932 14424 13938
rect 14554 13903 14610 13912
rect 14372 13874 14424 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13530 12572 13738
rect 13280 13530 13308 13874
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 12532 13524 12584 13530
rect 12532 13466 12584 13472
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10060 12442 10088 13330
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 10704 12782 10732 13126
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10152 12481 10180 12718
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10138 12472 10194 12481
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 10048 12436 10100 12442
rect 10289 12464 10585 12484
rect 10138 12407 10194 12416
rect 10048 12378 10100 12384
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9876 11762 9904 12038
rect 9864 11756 9916 11762
rect 9784 11716 9864 11744
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9508 10538 9536 11154
rect 9600 10810 9628 11222
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9496 10532 9548 10538
rect 9496 10474 9548 10480
rect 9508 10198 9536 10474
rect 9692 10198 9720 11562
rect 9784 11218 9812 11716
rect 9864 11698 9916 11704
rect 10048 11620 10100 11626
rect 10048 11562 10100 11568
rect 10060 11354 10088 11562
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10048 11348 10100 11354
rect 10100 11308 10180 11336
rect 10048 11290 10100 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 10048 10736 10100 10742
rect 10048 10678 10100 10684
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9680 10192 9732 10198
rect 9680 10134 9732 10140
rect 9678 10024 9734 10033
rect 9678 9959 9680 9968
rect 9732 9959 9734 9968
rect 9680 9930 9732 9936
rect 9784 8945 9812 10542
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10266 9904 10406
rect 10060 10266 10088 10678
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 9722 9904 9998
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9968 9586 9996 10134
rect 10060 9722 10088 10202
rect 10152 10062 10180 11308
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10704 10266 10732 10610
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 9770 8936 9826 8945
rect 9770 8871 9826 8880
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10796 7993 10824 12650
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10888 12345 10916 12582
rect 10874 12336 10930 12345
rect 10874 12271 10930 12280
rect 10980 8537 11008 12922
rect 11164 12850 11192 13126
rect 11900 12986 11928 13466
rect 12544 13410 12572 13466
rect 14016 13433 14044 13806
rect 14002 13424 14058 13433
rect 12544 13382 12664 13410
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11164 12374 11192 12786
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12268 12442 12296 12650
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11164 11898 11192 12310
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11256 11354 11284 12038
rect 11900 11898 11928 12242
rect 12360 12209 12388 12582
rect 12452 12442 12480 13262
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12544 12238 12572 12718
rect 12532 12232 12584 12238
rect 12346 12200 12402 12209
rect 12532 12174 12584 12180
rect 12346 12135 12402 12144
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 10966 8528 11022 8537
rect 10966 8463 11022 8472
rect 10782 7984 10838 7993
rect 10782 7919 10838 7928
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 9034 6216 9090 6225
rect 9034 6151 9090 6160
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 5446 3496 5502 3505
rect 5446 3431 5502 3440
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 3422 1456 3478 1465
rect 3422 1391 3478 1400
rect 7024 480 7052 4082
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 12636 1329 12664 13382
rect 14002 13359 14058 13368
rect 14568 12986 14596 13903
rect 15488 13841 15516 15982
rect 16316 15638 16344 22086
rect 16592 19394 16620 22374
rect 16500 19366 16620 19394
rect 16500 16114 16528 19366
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16132 15094 16160 15506
rect 16120 15088 16172 15094
rect 16118 15056 16120 15065
rect 16172 15056 16174 15065
rect 16118 14991 16174 15000
rect 16672 13864 16724 13870
rect 15474 13832 15530 13841
rect 16672 13806 16724 13812
rect 15474 13767 15530 13776
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 13820 12912 13872 12918
rect 13818 12880 13820 12889
rect 13872 12880 13874 12889
rect 13818 12815 13874 12824
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14660 12442 14688 12718
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 13096 11898 13124 12378
rect 13544 12368 13596 12374
rect 13542 12336 13544 12345
rect 13596 12336 13598 12345
rect 13542 12271 13598 12280
rect 13726 12336 13782 12345
rect 13726 12271 13782 12280
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 11898 13492 12174
rect 13556 11898 13584 12271
rect 13740 12102 13768 12271
rect 14660 12170 14688 12378
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 16684 9489 16712 13806
rect 17604 13462 17632 23530
rect 18064 14090 18092 23598
rect 18328 23520 18380 23526
rect 18524 23497 18552 27520
rect 18970 24712 19026 24721
rect 18970 24647 19026 24656
rect 18984 24410 19012 24647
rect 19076 24449 19104 27520
rect 19628 25786 19656 27520
rect 19444 25758 19656 25786
rect 19062 24440 19118 24449
rect 18972 24404 19024 24410
rect 19062 24375 19118 24384
rect 18972 24346 19024 24352
rect 18788 24268 18840 24274
rect 18788 24210 18840 24216
rect 18800 23526 18828 24210
rect 19248 23860 19300 23866
rect 19444 23848 19472 25758
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20272 23866 20300 27520
rect 20824 24721 20852 27520
rect 20810 24712 20866 24721
rect 20810 24647 20866 24656
rect 21180 24268 21232 24274
rect 21180 24210 21232 24216
rect 20442 24032 20498 24041
rect 20442 23967 20498 23976
rect 20456 23866 20484 23967
rect 19300 23820 19472 23848
rect 20260 23860 20312 23866
rect 19248 23802 19300 23808
rect 20260 23802 20312 23808
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 19984 23656 20036 23662
rect 19522 23624 19578 23633
rect 19984 23598 20036 23604
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 19522 23559 19578 23568
rect 18788 23520 18840 23526
rect 18328 23462 18380 23468
rect 18510 23488 18566 23497
rect 17880 14062 18092 14090
rect 17880 13938 17908 14062
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17420 12986 17448 13330
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 16670 9480 16726 9489
rect 16670 9415 16726 9424
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 17420 7857 17448 12922
rect 18340 11762 18368 23462
rect 18788 23462 18840 23468
rect 18510 23423 18566 23432
rect 19536 23322 19564 23559
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22438 19380 23122
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18064 10577 18092 11630
rect 18326 10704 18382 10713
rect 19352 10690 19380 22374
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 11121 19564 11154
rect 19522 11112 19578 11121
rect 19522 11047 19578 11056
rect 19536 10810 19564 11047
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19260 10674 19380 10690
rect 19996 10674 20024 23598
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20916 22438 20944 23122
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20812 12368 20864 12374
rect 20916 12345 20944 22374
rect 21008 12442 21036 23598
rect 21192 23526 21220 24210
rect 21376 23633 21404 27520
rect 21928 24041 21956 27520
rect 22480 24410 22508 27520
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 21914 24032 21970 24041
rect 21914 23967 21970 23976
rect 23124 23905 23152 27520
rect 21546 23896 21602 23905
rect 21546 23831 21548 23840
rect 21600 23831 21602 23840
rect 23110 23896 23166 23905
rect 23676 23882 23704 27520
rect 24228 24834 24256 27520
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 23400 23866 23704 23882
rect 23110 23831 23166 23840
rect 23388 23860 23704 23866
rect 21548 23802 21600 23808
rect 23440 23854 23704 23860
rect 23768 24806 24256 24834
rect 24674 24848 24730 24857
rect 23388 23802 23440 23808
rect 22100 23656 22152 23662
rect 21362 23624 21418 23633
rect 21362 23559 21418 23568
rect 22020 23604 22100 23610
rect 22020 23598 22152 23604
rect 22020 23582 22140 23598
rect 21180 23520 21232 23526
rect 21180 23462 21232 23468
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20812 12310 20864 12316
rect 20902 12336 20958 12345
rect 20824 11540 20852 12310
rect 20902 12271 20958 12280
rect 20904 11552 20956 11558
rect 20824 11512 20904 11540
rect 20904 11494 20956 11500
rect 18326 10639 18382 10648
rect 19248 10668 19380 10674
rect 18340 10606 18368 10639
rect 19300 10662 19380 10668
rect 19984 10668 20036 10674
rect 19248 10610 19300 10616
rect 19984 10610 20036 10616
rect 18328 10600 18380 10606
rect 18050 10568 18106 10577
rect 18328 10542 18380 10548
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 18050 10503 18106 10512
rect 19536 10169 19564 10542
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19522 10160 19578 10169
rect 19522 10095 19578 10104
rect 20916 10033 20944 11494
rect 21192 11286 21220 23462
rect 22020 23254 22048 23582
rect 22008 23248 22060 23254
rect 22008 23190 22060 23196
rect 23480 17264 23532 17270
rect 23480 17206 23532 17212
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 17406 7848 17462 7857
rect 17406 7783 17462 7792
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 22192 7336 22244 7342
rect 22190 7304 22192 7313
rect 22244 7304 22246 7313
rect 22190 7239 22246 7248
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 22742 6896 22798 6905
rect 22742 6831 22744 6840
rect 22796 6831 22798 6840
rect 22744 6802 22796 6808
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 22756 6458 22784 6802
rect 23492 6746 23520 17206
rect 23768 12594 23796 24806
rect 24674 24783 24730 24792
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 23676 12566 23796 12594
rect 23676 12458 23704 12566
rect 23584 12430 23704 12458
rect 23584 7546 23612 12430
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23400 6730 23520 6746
rect 23388 6724 23520 6730
rect 23440 6718 23520 6724
rect 23388 6666 23440 6672
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 23662 6352 23718 6361
rect 23662 6287 23718 6296
rect 23676 6254 23704 6287
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 23938 5808 23994 5817
rect 23938 5743 23940 5752
rect 23992 5743 23994 5752
rect 23940 5714 23992 5720
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 23952 5370 23980 5714
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 24783
rect 24780 17270 24808 27520
rect 25332 19378 25360 27520
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 25320 19372 25372 19378
rect 25320 19314 25372 19320
rect 24768 17264 24820 17270
rect 24768 17206 24820 17212
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24872 5930 24900 17206
rect 25056 6458 25084 19314
rect 25976 17270 26004 27520
rect 26528 24857 26556 27520
rect 26514 24848 26570 24857
rect 27080 24834 27108 27520
rect 26514 24783 26570 24792
rect 26712 24806 27108 24834
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 26712 17082 26740 24806
rect 27632 18193 27660 27520
rect 27618 18184 27674 18193
rect 27618 18119 27674 18128
rect 26344 17054 26740 17082
rect 25044 6452 25096 6458
rect 25044 6394 25096 6400
rect 24780 5914 24900 5930
rect 24768 5908 24900 5914
rect 24820 5902 24900 5908
rect 24768 5850 24820 5856
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24490 5264 24546 5273
rect 24490 5199 24546 5208
rect 24504 5166 24532 5199
rect 24492 5160 24544 5166
rect 24492 5102 24544 5108
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 26344 4865 26372 17054
rect 24766 4856 24822 4865
rect 24766 4791 24768 4800
rect 24820 4791 24822 4800
rect 26330 4856 26386 4865
rect 26330 4791 26386 4800
rect 24768 4762 24820 4768
rect 24582 4720 24638 4729
rect 24582 4655 24584 4664
rect 24636 4655 24638 4664
rect 24584 4626 24636 4632
rect 24596 4570 24624 4626
rect 24596 4542 24716 4570
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24688 4282 24716 4542
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 20994 3496 21050 3505
rect 20994 3431 21050 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 12622 1320 12678 1329
rect 12622 1255 12678 1264
rect 21008 480 21036 3431
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 2962 368 3018 377
rect 2962 303 3018 312
rect 7010 0 7066 480
rect 20994 0 21050 480
<< via2 >>
rect 3514 27648 3570 27704
rect 294 24384 350 24440
rect 1398 21528 1454 21584
rect 846 18808 902 18864
rect 1766 24148 1768 24168
rect 1768 24148 1820 24168
rect 1820 24148 1822 24168
rect 1766 24112 1822 24148
rect 1582 23432 1638 23488
rect 1950 23588 2006 23624
rect 1950 23568 1952 23588
rect 1952 23568 2004 23588
rect 2004 23568 2006 23588
rect 1950 21004 2006 21040
rect 1950 20984 1952 21004
rect 1952 20984 2004 21004
rect 2004 20984 2006 21004
rect 2502 23860 2558 23896
rect 2502 23840 2504 23860
rect 2504 23840 2556 23860
rect 2556 23840 2558 23860
rect 2870 24268 2926 24304
rect 2870 24248 2872 24268
rect 2872 24248 2924 24268
rect 2924 24248 2926 24268
rect 2778 23976 2834 24032
rect 2226 23160 2282 23216
rect 1582 17332 1638 17368
rect 1582 17312 1584 17332
rect 1584 17312 1636 17332
rect 1636 17312 1638 17332
rect 1490 16632 1546 16688
rect 2502 23024 2558 23080
rect 2410 22380 2412 22400
rect 2412 22380 2464 22400
rect 2464 22380 2466 22400
rect 2410 22344 2466 22380
rect 2410 22072 2466 22128
rect 2410 20476 2412 20496
rect 2412 20476 2464 20496
rect 2464 20476 2466 20496
rect 2410 20440 2466 20476
rect 2042 19352 2098 19408
rect 1950 19216 2006 19272
rect 1582 16496 1638 16552
rect 1674 16088 1730 16144
rect 1582 15952 1638 16008
rect 1398 14592 1454 14648
rect 2686 20848 2742 20904
rect 2962 22752 3018 22808
rect 3054 22208 3110 22264
rect 2962 21256 3018 21312
rect 2870 20304 2926 20360
rect 2962 19352 3018 19408
rect 2870 18828 2926 18864
rect 2870 18808 2872 18828
rect 2872 18808 2924 18828
rect 2924 18808 2926 18828
rect 2778 18128 2834 18184
rect 2594 17448 2650 17504
rect 2594 17312 2650 17368
rect 1858 15444 1860 15464
rect 1860 15444 1912 15464
rect 1912 15444 1914 15464
rect 1858 15408 1914 15444
rect 4066 27104 4122 27160
rect 4066 26444 4122 26480
rect 4066 26424 4068 26444
rect 4068 26424 4120 26444
rect 4120 26424 4122 26444
rect 4066 25880 4122 25936
rect 4066 25200 4122 25256
rect 3514 21428 3516 21448
rect 3516 21428 3568 21448
rect 3568 21428 3570 21448
rect 3514 21392 3570 21428
rect 3698 22500 3754 22536
rect 3698 22480 3700 22500
rect 3700 22480 3752 22500
rect 3752 22480 3754 22500
rect 3698 21936 3754 21992
rect 4066 20032 4122 20088
rect 4158 19916 4214 19952
rect 4158 19896 4160 19916
rect 4160 19896 4212 19916
rect 4212 19896 4214 19916
rect 3974 19760 4030 19816
rect 3698 17992 3754 18048
rect 1766 13096 1822 13152
rect 2502 12416 2558 12472
rect 2686 12416 2742 12472
rect 1490 10512 1546 10568
rect 1766 11192 1822 11248
rect 2502 11756 2558 11792
rect 2502 11736 2504 11756
rect 2504 11736 2556 11756
rect 2556 11736 2558 11756
rect 2870 11872 2926 11928
rect 2778 9560 2834 9616
rect 2594 8472 2650 8528
rect 3054 9560 3110 9616
rect 4066 19080 4122 19136
rect 4250 18572 4252 18592
rect 4252 18572 4304 18592
rect 4304 18572 4306 18592
rect 4250 18536 4306 18572
rect 4250 17876 4306 17912
rect 4250 17856 4252 17876
rect 4252 17856 4304 17876
rect 4304 17856 4306 17876
rect 4066 17740 4122 17776
rect 4066 17720 4068 17740
rect 4068 17720 4120 17740
rect 4120 17720 4122 17740
rect 3882 17620 3884 17640
rect 3884 17620 3936 17640
rect 3936 17620 3938 17640
rect 3882 17584 3938 17620
rect 3790 17312 3846 17368
rect 4618 19216 4674 19272
rect 3698 15000 3754 15056
rect 3974 15000 4030 15056
rect 3698 14884 3754 14920
rect 3698 14864 3700 14884
rect 3700 14864 3752 14884
rect 3752 14864 3754 14884
rect 3882 14476 3938 14512
rect 3882 14456 3884 14476
rect 3884 14456 3936 14476
rect 3936 14456 3938 14476
rect 3238 9424 3294 9480
rect 3698 10648 3754 10704
rect 4158 14320 4214 14376
rect 4158 13368 4214 13424
rect 3974 10648 4030 10704
rect 3974 10376 4030 10432
rect 5170 23840 5226 23896
rect 5078 23740 5080 23760
rect 5080 23740 5132 23760
rect 5132 23740 5134 23760
rect 5078 23704 5134 23740
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 6090 24792 6146 24848
rect 5538 24656 5594 24712
rect 5354 24520 5410 24576
rect 5354 24112 5410 24168
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5262 23432 5318 23488
rect 5170 22616 5226 22672
rect 5354 23296 5410 23352
rect 6274 24384 6330 24440
rect 5998 23160 6054 23216
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5998 21800 6054 21856
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5538 21392 5594 21448
rect 5446 21120 5502 21176
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5078 19780 5134 19816
rect 5078 19760 5080 19780
rect 5080 19760 5132 19780
rect 5132 19760 5134 19780
rect 4986 19236 5042 19272
rect 4986 19216 4988 19236
rect 4988 19216 5040 19236
rect 5040 19216 5042 19236
rect 4894 18944 4950 19000
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5078 17448 5134 17504
rect 4434 14612 4490 14648
rect 4434 14592 4436 14612
rect 4436 14592 4488 14612
rect 4488 14592 4490 14612
rect 4434 13776 4490 13832
rect 4342 12688 4398 12744
rect 2962 6160 3018 6216
rect 2594 2624 2650 2680
rect 3422 6704 3478 6760
rect 3330 3304 3386 3360
rect 4342 9696 4398 9752
rect 4986 14456 5042 14512
rect 4802 12824 4858 12880
rect 4894 11772 4896 11792
rect 4896 11772 4948 11792
rect 4948 11772 4950 11792
rect 4894 11736 4950 11772
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 6550 23296 6606 23352
rect 7010 24384 7066 24440
rect 7102 23432 7158 23488
rect 6918 23160 6974 23216
rect 6826 23024 6882 23080
rect 7746 23432 7802 23488
rect 8022 23296 8078 23352
rect 8482 23740 8484 23760
rect 8484 23740 8536 23760
rect 8536 23740 8538 23760
rect 8482 23704 8538 23740
rect 8666 23568 8722 23624
rect 8850 23432 8906 23488
rect 6458 21292 6460 21312
rect 6460 21292 6512 21312
rect 6512 21292 6514 21312
rect 6458 21256 6514 21292
rect 9678 24792 9734 24848
rect 9402 23296 9458 23352
rect 9310 22616 9366 22672
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5906 17176 5962 17232
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5998 16244 6054 16280
rect 5998 16224 6000 16244
rect 6000 16224 6052 16244
rect 6052 16224 6054 16244
rect 5170 13232 5226 13288
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5722 14456 5778 14512
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5170 12144 5226 12200
rect 5170 10376 5226 10432
rect 4526 9968 4582 10024
rect 4710 9968 4766 10024
rect 4066 7812 4122 7848
rect 4066 7792 4068 7812
rect 4068 7792 4120 7812
rect 4120 7792 4122 7812
rect 3882 3848 3938 3904
rect 5906 12280 5962 12336
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 6826 18400 6882 18456
rect 6550 18028 6552 18048
rect 6552 18028 6604 18048
rect 6604 18028 6606 18048
rect 6550 17992 6606 18028
rect 8482 22344 8538 22400
rect 8298 21664 8354 21720
rect 8022 20848 8078 20904
rect 9402 22072 9458 22128
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10046 24520 10102 24576
rect 9862 24248 9918 24304
rect 9678 22616 9734 22672
rect 9310 21392 9366 21448
rect 8206 20576 8262 20632
rect 8390 20032 8446 20088
rect 10230 24676 10286 24712
rect 10230 24656 10232 24676
rect 10232 24656 10284 24676
rect 10284 24656 10286 24676
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 9770 22072 9826 22128
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 8390 18808 8446 18864
rect 7654 18672 7710 18728
rect 8390 18128 8446 18184
rect 6182 13640 6238 13696
rect 7654 17040 7710 17096
rect 6826 14048 6882 14104
rect 6274 12280 6330 12336
rect 6550 12280 6606 12336
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6826 13948 6828 13968
rect 6828 13948 6880 13968
rect 6880 13948 6882 13968
rect 6826 13912 6882 13948
rect 7010 12824 7066 12880
rect 6642 10104 6698 10160
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 8758 18400 8814 18456
rect 8666 18148 8722 18184
rect 8666 18128 8668 18148
rect 8668 18128 8720 18148
rect 8720 18128 8722 18148
rect 8482 17720 8538 17776
rect 9402 18672 9458 18728
rect 8574 17176 8630 17232
rect 9034 16224 9090 16280
rect 8390 15272 8446 15328
rect 8482 14864 8538 14920
rect 7746 13268 7748 13288
rect 7748 13268 7800 13288
rect 7800 13268 7802 13288
rect 7746 13232 7802 13268
rect 7838 11076 7894 11112
rect 7838 11056 7840 11076
rect 7840 11056 7892 11076
rect 7892 11056 7894 11076
rect 7746 9968 7802 10024
rect 7654 9288 7710 9344
rect 9310 16496 9366 16552
rect 9218 14184 9274 14240
rect 9034 14048 9090 14104
rect 8206 12860 8208 12880
rect 8208 12860 8260 12880
rect 8260 12860 8262 12880
rect 8206 12824 8262 12860
rect 8850 12724 8852 12744
rect 8852 12724 8904 12744
rect 8904 12724 8906 12744
rect 8850 12688 8906 12724
rect 8298 12316 8300 12336
rect 8300 12316 8352 12336
rect 8352 12316 8354 12336
rect 8298 12280 8354 12316
rect 8114 12164 8170 12200
rect 8114 12144 8116 12164
rect 8116 12144 8168 12164
rect 8168 12144 8170 12164
rect 8298 12144 8354 12200
rect 7930 6704 7986 6760
rect 9770 19080 9826 19136
rect 9770 18944 9826 19000
rect 10782 21936 10838 21992
rect 10138 21392 10194 21448
rect 10046 19760 10102 19816
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 11978 24268 12034 24304
rect 11978 24248 11980 24268
rect 11980 24248 12032 24268
rect 12032 24248 12034 24268
rect 11334 21800 11390 21856
rect 11242 21392 11298 21448
rect 10414 20596 10470 20632
rect 10414 20576 10416 20596
rect 10416 20576 10468 20596
rect 10468 20576 10470 20596
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 11058 19896 11114 19952
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10966 18536 11022 18592
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9586 14864 9642 14920
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 9586 12844 9642 12880
rect 9586 12824 9588 12844
rect 9588 12824 9640 12844
rect 9640 12824 9642 12844
rect 10690 16088 10746 16144
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 11058 14864 11114 14920
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 11886 21004 11942 21040
rect 11886 20984 11888 21004
rect 11888 20984 11940 21004
rect 11940 20984 11942 21004
rect 11886 19488 11942 19544
rect 13266 24792 13322 24848
rect 12346 24148 12348 24168
rect 12348 24148 12400 24168
rect 12400 24148 12402 24168
rect 12346 24112 12402 24148
rect 12898 21528 12954 21584
rect 12162 16632 12218 16688
rect 11978 15272 12034 15328
rect 11886 14764 11888 14784
rect 11888 14764 11940 14784
rect 11940 14764 11942 14784
rect 11886 14728 11942 14764
rect 11702 14220 11704 14240
rect 11704 14220 11756 14240
rect 11756 14220 11758 14240
rect 11702 14184 11758 14220
rect 10138 13776 10194 13832
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 13542 24520 13598 24576
rect 13450 21684 13506 21720
rect 13450 21664 13452 21684
rect 13452 21664 13504 21684
rect 13504 21664 13506 21684
rect 12714 17040 12770 17096
rect 14554 24792 14610 24848
rect 14002 24676 14058 24712
rect 14002 24656 14004 24676
rect 14004 24656 14056 24676
rect 14056 24656 14058 24676
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 14830 24520 14886 24576
rect 14278 24112 14334 24168
rect 13634 18672 13690 18728
rect 12622 16088 12678 16144
rect 14002 17620 14004 17640
rect 14004 17620 14056 17640
rect 14056 17620 14058 17640
rect 14002 17584 14058 17620
rect 14094 14728 14150 14784
rect 12898 14320 12954 14376
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15382 23160 15438 23216
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 22072 15438 22128
rect 15290 21528 15346 21584
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14462 19488 14518 19544
rect 15198 20440 15254 20496
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15290 19216 15346 19272
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14922 16632 14978 16688
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 17682 24384 17738 24440
rect 16394 23860 16450 23896
rect 16394 23840 16396 23860
rect 16396 23840 16448 23860
rect 16448 23840 16450 23860
rect 17406 23840 17462 23896
rect 15750 18808 15806 18864
rect 16302 22480 16358 22536
rect 16762 23432 16818 23488
rect 15290 15988 15292 16008
rect 15292 15988 15344 16008
rect 15344 15988 15346 16008
rect 15290 15952 15346 15988
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15382 14320 15438 14376
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14554 13912 14610 13968
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10138 12416 10194 12472
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 9678 9988 9734 10024
rect 9678 9968 9680 9988
rect 9680 9968 9732 9988
rect 9732 9968 9734 9988
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 9770 8880 9826 8936
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10874 12280 10930 12336
rect 12346 12144 12402 12200
rect 10966 8472 11022 8528
rect 10782 7928 10838 7984
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 9034 6160 9090 6216
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 5446 3440 5502 3496
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 3422 1400 3478 1456
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 14002 13368 14058 13424
rect 16118 15036 16120 15056
rect 16120 15036 16172 15056
rect 16172 15036 16174 15056
rect 16118 15000 16174 15036
rect 15474 13776 15530 13832
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 13818 12860 13820 12880
rect 13820 12860 13872 12880
rect 13872 12860 13874 12880
rect 13818 12824 13874 12860
rect 13542 12316 13544 12336
rect 13544 12316 13596 12336
rect 13596 12316 13598 12336
rect 13542 12280 13598 12316
rect 13726 12280 13782 12336
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 18970 24656 19026 24712
rect 19062 24384 19118 24440
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20810 24656 20866 24712
rect 20442 23976 20498 24032
rect 19522 23568 19578 23624
rect 16670 9424 16726 9480
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 18510 23432 18566 23488
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 18326 10648 18382 10704
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19522 11056 19578 11112
rect 21914 23976 21970 24032
rect 21546 23860 21602 23896
rect 21546 23840 21548 23860
rect 21548 23840 21600 23860
rect 21600 23840 21602 23860
rect 23110 23840 23166 23896
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 21362 23568 21418 23624
rect 20902 12280 20958 12336
rect 18050 10512 18106 10568
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19522 10104 19578 10160
rect 20902 9968 20958 10024
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 17406 7792 17462 7848
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 22190 7284 22192 7304
rect 22192 7284 22244 7304
rect 22244 7284 22246 7304
rect 22190 7248 22246 7284
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 22742 6860 22798 6896
rect 22742 6840 22744 6860
rect 22744 6840 22796 6860
rect 22796 6840 22798 6860
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 24674 24792 24730 24848
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 23662 6296 23718 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 23938 5772 23994 5808
rect 23938 5752 23940 5772
rect 23940 5752 23992 5772
rect 23992 5752 23994 5772
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 26514 24792 26570 24848
rect 27618 18128 27674 18184
rect 24490 5208 24546 5264
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24766 4820 24822 4856
rect 24766 4800 24768 4820
rect 24768 4800 24820 4820
rect 24820 4800 24822 4820
rect 26330 4800 26386 4856
rect 24582 4684 24638 4720
rect 24582 4664 24584 4684
rect 24584 4664 24636 4684
rect 24636 4664 24638 4684
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 20994 3440 21050 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 12622 1264 12678 1320
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 2962 312 3018 368
<< metal3 >>
rect 0 27706 480 27736
rect 3509 27706 3575 27709
rect 0 27704 3575 27706
rect 0 27648 3514 27704
rect 3570 27648 3575 27704
rect 0 27646 3575 27648
rect 0 27616 480 27646
rect 3509 27643 3575 27646
rect 0 27162 480 27192
rect 4061 27162 4127 27165
rect 0 27160 4127 27162
rect 0 27104 4066 27160
rect 4122 27104 4127 27160
rect 0 27102 4127 27104
rect 0 27072 480 27102
rect 4061 27099 4127 27102
rect 0 26482 480 26512
rect 4061 26482 4127 26485
rect 0 26480 4127 26482
rect 0 26424 4066 26480
rect 4122 26424 4127 26480
rect 0 26422 4127 26424
rect 0 26392 480 26422
rect 4061 26419 4127 26422
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 0 25258 480 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 480 25198
rect 4061 25195 4127 25198
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 6085 24850 6151 24853
rect 9673 24850 9739 24853
rect 6085 24848 9739 24850
rect 6085 24792 6090 24848
rect 6146 24792 9678 24848
rect 9734 24792 9739 24848
rect 6085 24790 9739 24792
rect 6085 24787 6151 24790
rect 9673 24787 9739 24790
rect 13261 24850 13327 24853
rect 14549 24850 14615 24853
rect 13261 24848 14615 24850
rect 13261 24792 13266 24848
rect 13322 24792 14554 24848
rect 14610 24792 14615 24848
rect 13261 24790 14615 24792
rect 13261 24787 13327 24790
rect 14549 24787 14615 24790
rect 24669 24850 24735 24853
rect 26509 24850 26575 24853
rect 24669 24848 26575 24850
rect 24669 24792 24674 24848
rect 24730 24792 26514 24848
rect 26570 24792 26575 24848
rect 24669 24790 26575 24792
rect 24669 24787 24735 24790
rect 26509 24787 26575 24790
rect 0 24714 480 24744
rect 5533 24714 5599 24717
rect 0 24712 5599 24714
rect 0 24656 5538 24712
rect 5594 24656 5599 24712
rect 0 24654 5599 24656
rect 0 24624 480 24654
rect 5533 24651 5599 24654
rect 10225 24714 10291 24717
rect 13997 24714 14063 24717
rect 10225 24712 14063 24714
rect 10225 24656 10230 24712
rect 10286 24656 14002 24712
rect 14058 24656 14063 24712
rect 10225 24654 14063 24656
rect 10225 24651 10291 24654
rect 13997 24651 14063 24654
rect 18965 24714 19031 24717
rect 20805 24714 20871 24717
rect 18965 24712 20871 24714
rect 18965 24656 18970 24712
rect 19026 24656 20810 24712
rect 20866 24656 20871 24712
rect 18965 24654 20871 24656
rect 18965 24651 19031 24654
rect 20805 24651 20871 24654
rect 5349 24578 5415 24581
rect 10041 24578 10107 24581
rect 5349 24576 10107 24578
rect 5349 24520 5354 24576
rect 5410 24520 10046 24576
rect 10102 24520 10107 24576
rect 5349 24518 10107 24520
rect 5349 24515 5415 24518
rect 10041 24515 10107 24518
rect 13537 24578 13603 24581
rect 14825 24578 14891 24581
rect 13537 24576 14891 24578
rect 13537 24520 13542 24576
rect 13598 24520 14830 24576
rect 14886 24520 14891 24576
rect 13537 24518 14891 24520
rect 13537 24515 13603 24518
rect 14825 24515 14891 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 289 24442 355 24445
rect 6269 24442 6335 24445
rect 289 24440 6335 24442
rect 289 24384 294 24440
rect 350 24384 6274 24440
rect 6330 24384 6335 24440
rect 289 24382 6335 24384
rect 289 24379 355 24382
rect 6269 24379 6335 24382
rect 7005 24442 7071 24445
rect 17677 24442 17743 24445
rect 19057 24442 19123 24445
rect 7005 24440 10058 24442
rect 7005 24384 7010 24440
rect 7066 24384 10058 24440
rect 7005 24382 10058 24384
rect 7005 24379 7071 24382
rect 2865 24306 2931 24309
rect 9857 24306 9923 24309
rect 2865 24304 9923 24306
rect 2865 24248 2870 24304
rect 2926 24248 9862 24304
rect 9918 24248 9923 24304
rect 2865 24246 9923 24248
rect 9998 24306 10058 24382
rect 17677 24440 19123 24442
rect 17677 24384 17682 24440
rect 17738 24384 19062 24440
rect 19118 24384 19123 24440
rect 17677 24382 19123 24384
rect 17677 24379 17743 24382
rect 19057 24379 19123 24382
rect 11973 24306 12039 24309
rect 9998 24304 12039 24306
rect 9998 24248 11978 24304
rect 12034 24248 12039 24304
rect 9998 24246 12039 24248
rect 2865 24243 2931 24246
rect 9857 24243 9923 24246
rect 11973 24243 12039 24246
rect 1761 24170 1827 24173
rect 5349 24170 5415 24173
rect 1761 24168 5415 24170
rect 1761 24112 1766 24168
rect 1822 24112 5354 24168
rect 5410 24112 5415 24168
rect 1761 24110 5415 24112
rect 1761 24107 1827 24110
rect 5349 24107 5415 24110
rect 12341 24170 12407 24173
rect 14273 24170 14339 24173
rect 12341 24168 14339 24170
rect 12341 24112 12346 24168
rect 12402 24112 14278 24168
rect 14334 24112 14339 24168
rect 12341 24110 14339 24112
rect 12341 24107 12407 24110
rect 14273 24107 14339 24110
rect 0 24034 480 24064
rect 2773 24034 2839 24037
rect 0 24032 2839 24034
rect 0 23976 2778 24032
rect 2834 23976 2839 24032
rect 0 23974 2839 23976
rect 0 23944 480 23974
rect 2773 23971 2839 23974
rect 20437 24034 20503 24037
rect 21909 24034 21975 24037
rect 20437 24032 21975 24034
rect 20437 23976 20442 24032
rect 20498 23976 21914 24032
rect 21970 23976 21975 24032
rect 20437 23974 21975 23976
rect 20437 23971 20503 23974
rect 21909 23971 21975 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2497 23898 2563 23901
rect 5165 23898 5231 23901
rect 2497 23896 5231 23898
rect 2497 23840 2502 23896
rect 2558 23840 5170 23896
rect 5226 23840 5231 23896
rect 2497 23838 5231 23840
rect 2497 23835 2563 23838
rect 5165 23835 5231 23838
rect 16389 23898 16455 23901
rect 17401 23898 17467 23901
rect 16389 23896 17467 23898
rect 16389 23840 16394 23896
rect 16450 23840 17406 23896
rect 17462 23840 17467 23896
rect 16389 23838 17467 23840
rect 16389 23835 16455 23838
rect 17401 23835 17467 23838
rect 21541 23898 21607 23901
rect 23105 23898 23171 23901
rect 21541 23896 23171 23898
rect 21541 23840 21546 23896
rect 21602 23840 23110 23896
rect 23166 23840 23171 23896
rect 21541 23838 23171 23840
rect 21541 23835 21607 23838
rect 23105 23835 23171 23838
rect 5073 23762 5139 23765
rect 8477 23762 8543 23765
rect 5073 23760 8543 23762
rect 5073 23704 5078 23760
rect 5134 23704 8482 23760
rect 8538 23704 8543 23760
rect 5073 23702 8543 23704
rect 5073 23699 5139 23702
rect 8477 23699 8543 23702
rect 1945 23626 2011 23629
rect 8661 23626 8727 23629
rect 1945 23624 8727 23626
rect 1945 23568 1950 23624
rect 2006 23568 8666 23624
rect 8722 23568 8727 23624
rect 1945 23566 8727 23568
rect 1945 23563 2011 23566
rect 8661 23563 8727 23566
rect 19517 23626 19583 23629
rect 21357 23626 21423 23629
rect 19517 23624 21423 23626
rect 19517 23568 19522 23624
rect 19578 23568 21362 23624
rect 21418 23568 21423 23624
rect 19517 23566 21423 23568
rect 19517 23563 19583 23566
rect 21357 23563 21423 23566
rect 0 23490 480 23520
rect 1577 23490 1643 23493
rect 0 23488 1643 23490
rect 0 23432 1582 23488
rect 1638 23432 1643 23488
rect 0 23430 1643 23432
rect 0 23400 480 23430
rect 1577 23427 1643 23430
rect 5257 23490 5323 23493
rect 7097 23490 7163 23493
rect 5257 23488 7163 23490
rect 5257 23432 5262 23488
rect 5318 23432 7102 23488
rect 7158 23432 7163 23488
rect 5257 23430 7163 23432
rect 5257 23427 5323 23430
rect 7097 23427 7163 23430
rect 7741 23490 7807 23493
rect 8845 23490 8911 23493
rect 7741 23488 8911 23490
rect 7741 23432 7746 23488
rect 7802 23432 8850 23488
rect 8906 23432 8911 23488
rect 7741 23430 8911 23432
rect 7741 23427 7807 23430
rect 8845 23427 8911 23430
rect 16757 23490 16823 23493
rect 18505 23490 18571 23493
rect 16757 23488 18571 23490
rect 16757 23432 16762 23488
rect 16818 23432 18510 23488
rect 18566 23432 18571 23488
rect 16757 23430 18571 23432
rect 16757 23427 16823 23430
rect 18505 23427 18571 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5349 23354 5415 23357
rect 6545 23354 6611 23357
rect 5349 23352 6611 23354
rect 5349 23296 5354 23352
rect 5410 23296 6550 23352
rect 6606 23296 6611 23352
rect 5349 23294 6611 23296
rect 5349 23291 5415 23294
rect 6545 23291 6611 23294
rect 8017 23354 8083 23357
rect 9397 23354 9463 23357
rect 8017 23352 9463 23354
rect 8017 23296 8022 23352
rect 8078 23296 9402 23352
rect 9458 23296 9463 23352
rect 8017 23294 9463 23296
rect 8017 23291 8083 23294
rect 9397 23291 9463 23294
rect 2221 23218 2287 23221
rect 5993 23218 6059 23221
rect 2221 23216 6059 23218
rect 2221 23160 2226 23216
rect 2282 23160 5998 23216
rect 6054 23160 6059 23216
rect 2221 23158 6059 23160
rect 2221 23155 2287 23158
rect 5993 23155 6059 23158
rect 6913 23218 6979 23221
rect 15377 23218 15443 23221
rect 6913 23216 15443 23218
rect 6913 23160 6918 23216
rect 6974 23160 15382 23216
rect 15438 23160 15443 23216
rect 6913 23158 15443 23160
rect 6913 23155 6979 23158
rect 15377 23155 15443 23158
rect 2497 23082 2563 23085
rect 6821 23082 6887 23085
rect 2497 23080 6887 23082
rect 2497 23024 2502 23080
rect 2558 23024 6826 23080
rect 6882 23024 6887 23080
rect 2497 23022 6887 23024
rect 2497 23019 2563 23022
rect 6821 23019 6887 23022
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2957 22810 3023 22813
rect 0 22808 3023 22810
rect 0 22752 2962 22808
rect 3018 22752 3023 22808
rect 0 22750 3023 22752
rect 0 22720 480 22750
rect 2957 22747 3023 22750
rect 5165 22674 5231 22677
rect 9305 22674 9371 22677
rect 9673 22674 9739 22677
rect 5165 22672 9739 22674
rect 5165 22616 5170 22672
rect 5226 22616 9310 22672
rect 9366 22616 9678 22672
rect 9734 22616 9739 22672
rect 5165 22614 9739 22616
rect 5165 22611 5231 22614
rect 9305 22611 9371 22614
rect 9673 22611 9739 22614
rect 3693 22538 3759 22541
rect 16297 22538 16363 22541
rect 3693 22536 16363 22538
rect 3693 22480 3698 22536
rect 3754 22480 16302 22536
rect 16358 22480 16363 22536
rect 3693 22478 16363 22480
rect 3693 22475 3759 22478
rect 16297 22475 16363 22478
rect 2405 22402 2471 22405
rect 8477 22402 8543 22405
rect 2405 22400 8543 22402
rect 2405 22344 2410 22400
rect 2466 22344 8482 22400
rect 8538 22344 8543 22400
rect 2405 22342 8543 22344
rect 2405 22339 2471 22342
rect 8477 22339 8543 22342
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3049 22266 3115 22269
rect 0 22264 3115 22266
rect 0 22208 3054 22264
rect 3110 22208 3115 22264
rect 0 22206 3115 22208
rect 0 22176 480 22206
rect 3049 22203 3115 22206
rect 2405 22130 2471 22133
rect 9397 22130 9463 22133
rect 2405 22128 9463 22130
rect 2405 22072 2410 22128
rect 2466 22072 9402 22128
rect 9458 22072 9463 22128
rect 2405 22070 9463 22072
rect 2405 22067 2471 22070
rect 9397 22067 9463 22070
rect 9765 22130 9831 22133
rect 15377 22130 15443 22133
rect 9765 22128 15443 22130
rect 9765 22072 9770 22128
rect 9826 22072 15382 22128
rect 15438 22072 15443 22128
rect 9765 22070 15443 22072
rect 9765 22067 9831 22070
rect 15377 22067 15443 22070
rect 3693 21994 3759 21997
rect 10777 21994 10843 21997
rect 3693 21992 10843 21994
rect 3693 21936 3698 21992
rect 3754 21936 10782 21992
rect 10838 21936 10843 21992
rect 3693 21934 10843 21936
rect 3693 21931 3759 21934
rect 10777 21931 10843 21934
rect 5993 21858 6059 21861
rect 11329 21858 11395 21861
rect 5993 21856 11395 21858
rect 5993 21800 5998 21856
rect 6054 21800 11334 21856
rect 11390 21800 11395 21856
rect 5993 21798 11395 21800
rect 5993 21795 6059 21798
rect 11329 21795 11395 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 8293 21722 8359 21725
rect 13445 21722 13511 21725
rect 8293 21720 13511 21722
rect 8293 21664 8298 21720
rect 8354 21664 13450 21720
rect 13506 21664 13511 21720
rect 8293 21662 13511 21664
rect 8293 21659 8359 21662
rect 13445 21659 13511 21662
rect 0 21586 480 21616
rect 1393 21586 1459 21589
rect 0 21584 1459 21586
rect 0 21528 1398 21584
rect 1454 21528 1459 21584
rect 0 21526 1459 21528
rect 0 21496 480 21526
rect 1393 21523 1459 21526
rect 12893 21586 12959 21589
rect 15285 21586 15351 21589
rect 12893 21584 15351 21586
rect 12893 21528 12898 21584
rect 12954 21528 15290 21584
rect 15346 21528 15351 21584
rect 12893 21526 15351 21528
rect 12893 21523 12959 21526
rect 15285 21523 15351 21526
rect 3509 21450 3575 21453
rect 5533 21450 5599 21453
rect 3509 21448 5599 21450
rect 3509 21392 3514 21448
rect 3570 21392 5538 21448
rect 5594 21392 5599 21448
rect 3509 21390 5599 21392
rect 3509 21387 3575 21390
rect 5533 21387 5599 21390
rect 9305 21450 9371 21453
rect 10133 21450 10199 21453
rect 11237 21450 11303 21453
rect 9305 21448 11303 21450
rect 9305 21392 9310 21448
rect 9366 21392 10138 21448
rect 10194 21392 11242 21448
rect 11298 21392 11303 21448
rect 9305 21390 11303 21392
rect 9305 21387 9371 21390
rect 10133 21387 10199 21390
rect 11237 21387 11303 21390
rect 2957 21314 3023 21317
rect 6453 21314 6519 21317
rect 2957 21312 6519 21314
rect 2957 21256 2962 21312
rect 3018 21256 6458 21312
rect 6514 21256 6519 21312
rect 2957 21254 6519 21256
rect 2957 21251 3023 21254
rect 6453 21251 6519 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 5441 21178 5507 21181
rect 1350 21176 5507 21178
rect 1350 21120 5446 21176
rect 5502 21120 5507 21176
rect 1350 21118 5507 21120
rect 0 21042 480 21072
rect 1350 21042 1410 21118
rect 5441 21115 5507 21118
rect 0 20982 1410 21042
rect 1945 21042 2011 21045
rect 11881 21042 11947 21045
rect 1945 21040 11947 21042
rect 1945 20984 1950 21040
rect 2006 20984 11886 21040
rect 11942 20984 11947 21040
rect 1945 20982 11947 20984
rect 0 20952 480 20982
rect 1945 20979 2011 20982
rect 11881 20979 11947 20982
rect 2681 20906 2747 20909
rect 8017 20906 8083 20909
rect 2681 20904 8083 20906
rect 2681 20848 2686 20904
rect 2742 20848 8022 20904
rect 8078 20848 8083 20904
rect 2681 20846 8083 20848
rect 2681 20843 2747 20846
rect 8017 20843 8083 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 8201 20634 8267 20637
rect 10409 20634 10475 20637
rect 8201 20632 10475 20634
rect 8201 20576 8206 20632
rect 8262 20576 10414 20632
rect 10470 20576 10475 20632
rect 8201 20574 10475 20576
rect 8201 20571 8267 20574
rect 10409 20571 10475 20574
rect 2405 20498 2471 20501
rect 15193 20498 15259 20501
rect 2405 20496 15259 20498
rect 2405 20440 2410 20496
rect 2466 20440 15198 20496
rect 15254 20440 15259 20496
rect 2405 20438 15259 20440
rect 2405 20435 2471 20438
rect 15193 20435 15259 20438
rect 0 20362 480 20392
rect 2865 20362 2931 20365
rect 0 20360 2931 20362
rect 0 20304 2870 20360
rect 2926 20304 2931 20360
rect 0 20302 2931 20304
rect 0 20272 480 20302
rect 2865 20299 2931 20302
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 4061 20090 4127 20093
rect 8385 20090 8451 20093
rect 4061 20088 8451 20090
rect 4061 20032 4066 20088
rect 4122 20032 8390 20088
rect 8446 20032 8451 20088
rect 4061 20030 8451 20032
rect 4061 20027 4127 20030
rect 8385 20027 8451 20030
rect 4153 19954 4219 19957
rect 11053 19954 11119 19957
rect 4153 19952 11119 19954
rect 4153 19896 4158 19952
rect 4214 19896 11058 19952
rect 11114 19896 11119 19952
rect 4153 19894 11119 19896
rect 4153 19891 4219 19894
rect 11053 19891 11119 19894
rect 0 19818 480 19848
rect 3969 19818 4035 19821
rect 0 19816 4035 19818
rect 0 19760 3974 19816
rect 4030 19760 4035 19816
rect 0 19758 4035 19760
rect 0 19728 480 19758
rect 3969 19755 4035 19758
rect 5073 19818 5139 19821
rect 10041 19818 10107 19821
rect 5073 19816 10107 19818
rect 5073 19760 5078 19816
rect 5134 19760 10046 19816
rect 10102 19760 10107 19816
rect 5073 19758 10107 19760
rect 5073 19755 5139 19758
rect 10041 19755 10107 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 11881 19546 11947 19549
rect 14457 19546 14523 19549
rect 11881 19544 14523 19546
rect 11881 19488 11886 19544
rect 11942 19488 14462 19544
rect 14518 19488 14523 19544
rect 11881 19486 14523 19488
rect 11881 19483 11947 19486
rect 14457 19483 14523 19486
rect 2037 19410 2103 19413
rect 2957 19410 3023 19413
rect 2037 19408 3023 19410
rect 2037 19352 2042 19408
rect 2098 19352 2962 19408
rect 3018 19352 3023 19408
rect 2037 19350 3023 19352
rect 2037 19347 2103 19350
rect 2957 19347 3023 19350
rect 1945 19274 2011 19277
rect 4613 19274 4679 19277
rect 1945 19272 4679 19274
rect 1945 19216 1950 19272
rect 2006 19216 4618 19272
rect 4674 19216 4679 19272
rect 1945 19214 4679 19216
rect 1945 19211 2011 19214
rect 4613 19211 4679 19214
rect 4981 19274 5047 19277
rect 15285 19274 15351 19277
rect 4981 19272 15351 19274
rect 4981 19216 4986 19272
rect 5042 19216 15290 19272
rect 15346 19216 15351 19272
rect 4981 19214 15351 19216
rect 4981 19211 5047 19214
rect 15285 19211 15351 19214
rect 0 19138 480 19168
rect 4061 19138 4127 19141
rect 0 19136 4127 19138
rect 0 19080 4066 19136
rect 4122 19080 4127 19136
rect 0 19078 4127 19080
rect 0 19048 480 19078
rect 4061 19075 4127 19078
rect 9765 19138 9831 19141
rect 9990 19138 9996 19140
rect 9765 19136 9996 19138
rect 9765 19080 9770 19136
rect 9826 19080 9996 19136
rect 9765 19078 9996 19080
rect 9765 19075 9831 19078
rect 9990 19076 9996 19078
rect 10060 19076 10066 19140
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 4889 19002 4955 19005
rect 9765 19002 9831 19005
rect 4889 19000 9831 19002
rect 4889 18944 4894 19000
rect 4950 18944 9770 19000
rect 9826 18944 9831 19000
rect 4889 18942 9831 18944
rect 4889 18939 4955 18942
rect 9765 18939 9831 18942
rect 841 18866 907 18869
rect 2865 18866 2931 18869
rect 841 18864 2931 18866
rect 841 18808 846 18864
rect 902 18808 2870 18864
rect 2926 18808 2931 18864
rect 841 18806 2931 18808
rect 841 18803 907 18806
rect 2865 18803 2931 18806
rect 8385 18866 8451 18869
rect 15745 18866 15811 18869
rect 8385 18864 15811 18866
rect 8385 18808 8390 18864
rect 8446 18808 15750 18864
rect 15806 18808 15811 18864
rect 8385 18806 15811 18808
rect 8385 18803 8451 18806
rect 15745 18803 15811 18806
rect 7649 18730 7715 18733
rect 9397 18730 9463 18733
rect 13629 18730 13695 18733
rect 7649 18728 13695 18730
rect 7649 18672 7654 18728
rect 7710 18672 9402 18728
rect 9458 18672 13634 18728
rect 13690 18672 13695 18728
rect 7649 18670 13695 18672
rect 7649 18667 7715 18670
rect 9397 18667 9463 18670
rect 13629 18667 13695 18670
rect 0 18594 480 18624
rect 4245 18594 4311 18597
rect 0 18592 4311 18594
rect 0 18536 4250 18592
rect 4306 18536 4311 18592
rect 0 18534 4311 18536
rect 0 18504 480 18534
rect 4245 18531 4311 18534
rect 9990 18532 9996 18596
rect 10060 18594 10066 18596
rect 10961 18594 11027 18597
rect 10060 18592 11027 18594
rect 10060 18536 10966 18592
rect 11022 18536 11027 18592
rect 10060 18534 11027 18536
rect 10060 18532 10066 18534
rect 10961 18531 11027 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 6821 18458 6887 18461
rect 8753 18458 8819 18461
rect 6821 18456 8819 18458
rect 6821 18400 6826 18456
rect 6882 18400 8758 18456
rect 8814 18400 8819 18456
rect 6821 18398 8819 18400
rect 6821 18395 6887 18398
rect 8753 18395 8819 18398
rect 2773 18186 2839 18189
rect 8385 18186 8451 18189
rect 2773 18184 8451 18186
rect 2773 18128 2778 18184
rect 2834 18128 8390 18184
rect 8446 18128 8451 18184
rect 2773 18126 8451 18128
rect 2773 18123 2839 18126
rect 8385 18123 8451 18126
rect 8661 18186 8727 18189
rect 27613 18186 27679 18189
rect 8661 18184 27679 18186
rect 8661 18128 8666 18184
rect 8722 18128 27618 18184
rect 27674 18128 27679 18184
rect 8661 18126 27679 18128
rect 8661 18123 8727 18126
rect 27613 18123 27679 18126
rect 3693 18050 3759 18053
rect 6545 18050 6611 18053
rect 3693 18048 6611 18050
rect 3693 17992 3698 18048
rect 3754 17992 6550 18048
rect 6606 17992 6611 18048
rect 3693 17990 6611 17992
rect 3693 17987 3759 17990
rect 6545 17987 6611 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 4245 17914 4311 17917
rect 0 17912 4311 17914
rect 0 17856 4250 17912
rect 4306 17856 4311 17912
rect 0 17854 4311 17856
rect 0 17824 480 17854
rect 4245 17851 4311 17854
rect 4061 17778 4127 17781
rect 8477 17778 8543 17781
rect 4061 17776 8543 17778
rect 4061 17720 4066 17776
rect 4122 17720 8482 17776
rect 8538 17720 8543 17776
rect 4061 17718 8543 17720
rect 4061 17715 4127 17718
rect 8477 17715 8543 17718
rect 3877 17642 3943 17645
rect 13997 17642 14063 17645
rect 3877 17640 14063 17642
rect 3877 17584 3882 17640
rect 3938 17584 14002 17640
rect 14058 17584 14063 17640
rect 3877 17582 14063 17584
rect 3877 17579 3943 17582
rect 13997 17579 14063 17582
rect 2589 17506 2655 17509
rect 5073 17506 5139 17509
rect 2589 17504 5139 17506
rect 2589 17448 2594 17504
rect 2650 17448 5078 17504
rect 5134 17448 5139 17504
rect 2589 17446 5139 17448
rect 2589 17443 2655 17446
rect 5073 17443 5139 17446
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 1577 17370 1643 17373
rect 0 17368 1643 17370
rect 0 17312 1582 17368
rect 1638 17312 1643 17368
rect 0 17310 1643 17312
rect 0 17280 480 17310
rect 1577 17307 1643 17310
rect 2589 17370 2655 17373
rect 3785 17370 3851 17373
rect 2589 17368 3851 17370
rect 2589 17312 2594 17368
rect 2650 17312 3790 17368
rect 3846 17312 3851 17368
rect 2589 17310 3851 17312
rect 2589 17307 2655 17310
rect 3785 17307 3851 17310
rect 5901 17234 5967 17237
rect 8569 17234 8635 17237
rect 5901 17232 8635 17234
rect 5901 17176 5906 17232
rect 5962 17176 8574 17232
rect 8630 17176 8635 17232
rect 5901 17174 8635 17176
rect 5901 17171 5967 17174
rect 8569 17171 8635 17174
rect 7649 17098 7715 17101
rect 12709 17098 12775 17101
rect 7649 17096 12775 17098
rect 7649 17040 7654 17096
rect 7710 17040 12714 17096
rect 12770 17040 12775 17096
rect 7649 17038 12775 17040
rect 7649 17035 7715 17038
rect 12709 17035 12775 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 1485 16690 1551 16693
rect 0 16688 1551 16690
rect 0 16632 1490 16688
rect 1546 16632 1551 16688
rect 0 16630 1551 16632
rect 0 16600 480 16630
rect 1485 16627 1551 16630
rect 12157 16690 12223 16693
rect 14917 16690 14983 16693
rect 12157 16688 14983 16690
rect 12157 16632 12162 16688
rect 12218 16632 14922 16688
rect 14978 16632 14983 16688
rect 12157 16630 14983 16632
rect 12157 16627 12223 16630
rect 14917 16627 14983 16630
rect 1577 16554 1643 16557
rect 9305 16554 9371 16557
rect 1577 16552 9371 16554
rect 1577 16496 1582 16552
rect 1638 16496 9310 16552
rect 9366 16496 9371 16552
rect 1577 16494 9371 16496
rect 1577 16491 1643 16494
rect 9305 16491 9371 16494
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 5993 16282 6059 16285
rect 9029 16282 9095 16285
rect 5993 16280 9095 16282
rect 5993 16224 5998 16280
rect 6054 16224 9034 16280
rect 9090 16224 9095 16280
rect 5993 16222 9095 16224
rect 5993 16219 6059 16222
rect 9029 16219 9095 16222
rect 0 16146 480 16176
rect 1669 16146 1735 16149
rect 0 16144 1735 16146
rect 0 16088 1674 16144
rect 1730 16088 1735 16144
rect 0 16086 1735 16088
rect 0 16056 480 16086
rect 1669 16083 1735 16086
rect 10685 16146 10751 16149
rect 12617 16146 12683 16149
rect 10685 16144 12683 16146
rect 10685 16088 10690 16144
rect 10746 16088 12622 16144
rect 12678 16088 12683 16144
rect 10685 16086 12683 16088
rect 10685 16083 10751 16086
rect 12617 16083 12683 16086
rect 1577 16010 1643 16013
rect 15285 16010 15351 16013
rect 1577 16008 15351 16010
rect 1577 15952 1582 16008
rect 1638 15952 15290 16008
rect 15346 15952 15351 16008
rect 1577 15950 15351 15952
rect 1577 15947 1643 15950
rect 15285 15947 15351 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15466 480 15496
rect 1853 15466 1919 15469
rect 0 15464 1919 15466
rect 0 15408 1858 15464
rect 1914 15408 1919 15464
rect 0 15406 1919 15408
rect 0 15376 480 15406
rect 1853 15403 1919 15406
rect 8385 15330 8451 15333
rect 11973 15330 12039 15333
rect 8385 15328 12039 15330
rect 8385 15272 8390 15328
rect 8446 15272 11978 15328
rect 12034 15272 12039 15328
rect 8385 15270 12039 15272
rect 8385 15267 8451 15270
rect 11973 15267 12039 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3693 15058 3759 15061
rect 1350 15056 3759 15058
rect 1350 15000 3698 15056
rect 3754 15000 3759 15056
rect 1350 14998 3759 15000
rect 0 14922 480 14952
rect 1350 14922 1410 14998
rect 3693 14995 3759 14998
rect 3969 15058 4035 15061
rect 16113 15058 16179 15061
rect 3969 15056 16179 15058
rect 3969 15000 3974 15056
rect 4030 15000 16118 15056
rect 16174 15000 16179 15056
rect 3969 14998 16179 15000
rect 3969 14995 4035 14998
rect 16113 14995 16179 14998
rect 0 14862 1410 14922
rect 3693 14922 3759 14925
rect 8477 14922 8543 14925
rect 3693 14920 8543 14922
rect 3693 14864 3698 14920
rect 3754 14864 8482 14920
rect 8538 14864 8543 14920
rect 3693 14862 8543 14864
rect 0 14832 480 14862
rect 3693 14859 3759 14862
rect 8477 14859 8543 14862
rect 9581 14922 9647 14925
rect 11053 14922 11119 14925
rect 9581 14920 11119 14922
rect 9581 14864 9586 14920
rect 9642 14864 11058 14920
rect 11114 14864 11119 14920
rect 9581 14862 11119 14864
rect 9581 14859 9647 14862
rect 11053 14859 11119 14862
rect 11881 14786 11947 14789
rect 14089 14786 14155 14789
rect 11881 14784 14155 14786
rect 11881 14728 11886 14784
rect 11942 14728 14094 14784
rect 14150 14728 14155 14784
rect 11881 14726 14155 14728
rect 11881 14723 11947 14726
rect 14089 14723 14155 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1393 14650 1459 14653
rect 4429 14650 4495 14653
rect 1393 14648 4495 14650
rect 1393 14592 1398 14648
rect 1454 14592 4434 14648
rect 4490 14592 4495 14648
rect 1393 14590 4495 14592
rect 1393 14587 1459 14590
rect 4429 14587 4495 14590
rect 3877 14514 3943 14517
rect 4981 14514 5047 14517
rect 5717 14514 5783 14517
rect 3877 14512 5783 14514
rect 3877 14456 3882 14512
rect 3938 14456 4986 14512
rect 5042 14456 5722 14512
rect 5778 14456 5783 14512
rect 3877 14454 5783 14456
rect 3877 14451 3943 14454
rect 4981 14451 5047 14454
rect 5717 14451 5783 14454
rect 0 14378 480 14408
rect 4153 14378 4219 14381
rect 0 14376 4219 14378
rect 0 14320 4158 14376
rect 4214 14320 4219 14376
rect 0 14318 4219 14320
rect 0 14288 480 14318
rect 4153 14315 4219 14318
rect 12893 14378 12959 14381
rect 15377 14378 15443 14381
rect 12893 14376 15443 14378
rect 12893 14320 12898 14376
rect 12954 14320 15382 14376
rect 15438 14320 15443 14376
rect 12893 14318 15443 14320
rect 12893 14315 12959 14318
rect 15377 14315 15443 14318
rect 9213 14242 9279 14245
rect 11697 14242 11763 14245
rect 9213 14240 11763 14242
rect 9213 14184 9218 14240
rect 9274 14184 11702 14240
rect 11758 14184 11763 14240
rect 9213 14182 11763 14184
rect 9213 14179 9279 14182
rect 11697 14179 11763 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 6821 14106 6887 14109
rect 9029 14106 9095 14109
rect 27520 14106 28000 14136
rect 6821 14104 9095 14106
rect 6821 14048 6826 14104
rect 6882 14048 9034 14104
rect 9090 14048 9095 14104
rect 6821 14046 9095 14048
rect 6821 14043 6887 14046
rect 9029 14043 9095 14046
rect 24902 14046 28000 14106
rect 6821 13970 6887 13973
rect 14549 13970 14615 13973
rect 24902 13970 24962 14046
rect 27520 14016 28000 14046
rect 6821 13968 14474 13970
rect 6821 13912 6826 13968
rect 6882 13912 14474 13968
rect 6821 13910 14474 13912
rect 6821 13907 6887 13910
rect 4429 13834 4495 13837
rect 10133 13834 10199 13837
rect 4429 13832 10199 13834
rect 4429 13776 4434 13832
rect 4490 13776 10138 13832
rect 10194 13776 10199 13832
rect 4429 13774 10199 13776
rect 14414 13834 14474 13910
rect 14549 13968 24962 13970
rect 14549 13912 14554 13968
rect 14610 13912 24962 13968
rect 14549 13910 24962 13912
rect 14549 13907 14615 13910
rect 15469 13834 15535 13837
rect 14414 13832 15535 13834
rect 14414 13776 15474 13832
rect 15530 13776 15535 13832
rect 14414 13774 15535 13776
rect 4429 13771 4495 13774
rect 10133 13771 10199 13774
rect 15469 13771 15535 13774
rect 0 13698 480 13728
rect 6177 13698 6243 13701
rect 0 13696 6243 13698
rect 0 13640 6182 13696
rect 6238 13640 6243 13696
rect 0 13638 6243 13640
rect 0 13608 480 13638
rect 6177 13635 6243 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4153 13426 4219 13429
rect 13997 13426 14063 13429
rect 4153 13424 14063 13426
rect 4153 13368 4158 13424
rect 4214 13368 14002 13424
rect 14058 13368 14063 13424
rect 4153 13366 14063 13368
rect 4153 13363 4219 13366
rect 13997 13363 14063 13366
rect 5165 13290 5231 13293
rect 7741 13290 7807 13293
rect 5165 13288 7807 13290
rect 5165 13232 5170 13288
rect 5226 13232 7746 13288
rect 7802 13232 7807 13288
rect 5165 13230 7807 13232
rect 5165 13227 5231 13230
rect 7741 13227 7807 13230
rect 0 13154 480 13184
rect 1761 13154 1827 13157
rect 0 13152 1827 13154
rect 0 13096 1766 13152
rect 1822 13096 1827 13152
rect 0 13094 1827 13096
rect 0 13064 480 13094
rect 1761 13091 1827 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 4797 12882 4863 12885
rect 7005 12882 7071 12885
rect 8201 12882 8267 12885
rect 4797 12880 8267 12882
rect 4797 12824 4802 12880
rect 4858 12824 7010 12880
rect 7066 12824 8206 12880
rect 8262 12824 8267 12880
rect 4797 12822 8267 12824
rect 4797 12819 4863 12822
rect 7005 12819 7071 12822
rect 8201 12819 8267 12822
rect 9581 12882 9647 12885
rect 13813 12882 13879 12885
rect 9581 12880 13879 12882
rect 9581 12824 9586 12880
rect 9642 12824 13818 12880
rect 13874 12824 13879 12880
rect 9581 12822 13879 12824
rect 9581 12819 9647 12822
rect 13813 12819 13879 12822
rect 4337 12746 4403 12749
rect 8845 12746 8911 12749
rect 4337 12744 8911 12746
rect 4337 12688 4342 12744
rect 4398 12688 8850 12744
rect 8906 12688 8911 12744
rect 4337 12686 8911 12688
rect 4337 12683 4403 12686
rect 8845 12683 8911 12686
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 2497 12474 2563 12477
rect 0 12472 2563 12474
rect 0 12416 2502 12472
rect 2558 12416 2563 12472
rect 0 12414 2563 12416
rect 0 12384 480 12414
rect 2497 12411 2563 12414
rect 2681 12474 2747 12477
rect 10133 12474 10199 12477
rect 2681 12472 10199 12474
rect 2681 12416 2686 12472
rect 2742 12416 10138 12472
rect 10194 12416 10199 12472
rect 2681 12414 10199 12416
rect 2681 12411 2747 12414
rect 10133 12411 10199 12414
rect 5901 12338 5967 12341
rect 6269 12338 6335 12341
rect 5901 12336 6335 12338
rect 5901 12280 5906 12336
rect 5962 12280 6274 12336
rect 6330 12280 6335 12336
rect 5901 12278 6335 12280
rect 5901 12275 5967 12278
rect 6269 12275 6335 12278
rect 6545 12338 6611 12341
rect 8293 12338 8359 12341
rect 6545 12336 8359 12338
rect 6545 12280 6550 12336
rect 6606 12280 8298 12336
rect 8354 12280 8359 12336
rect 6545 12278 8359 12280
rect 6545 12275 6611 12278
rect 8293 12275 8359 12278
rect 10869 12338 10935 12341
rect 13537 12338 13603 12341
rect 10869 12336 13603 12338
rect 10869 12280 10874 12336
rect 10930 12280 13542 12336
rect 13598 12280 13603 12336
rect 10869 12278 13603 12280
rect 10869 12275 10935 12278
rect 13537 12275 13603 12278
rect 13721 12338 13787 12341
rect 20897 12338 20963 12341
rect 13721 12336 20963 12338
rect 13721 12280 13726 12336
rect 13782 12280 20902 12336
rect 20958 12280 20963 12336
rect 13721 12278 20963 12280
rect 13721 12275 13787 12278
rect 20897 12275 20963 12278
rect 5165 12202 5231 12205
rect 8109 12202 8175 12205
rect 5165 12200 8175 12202
rect 5165 12144 5170 12200
rect 5226 12144 8114 12200
rect 8170 12144 8175 12200
rect 5165 12142 8175 12144
rect 5165 12139 5231 12142
rect 8109 12139 8175 12142
rect 8293 12202 8359 12205
rect 12341 12202 12407 12205
rect 8293 12200 9506 12202
rect 8293 12144 8298 12200
rect 8354 12168 9506 12200
rect 9630 12200 12407 12202
rect 9630 12168 12346 12200
rect 8354 12144 12346 12168
rect 12402 12144 12407 12200
rect 8293 12142 12407 12144
rect 8293 12139 8359 12142
rect 9446 12108 9690 12142
rect 12341 12139 12407 12142
rect 9584 12040 9690 12108
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 2865 11930 2931 11933
rect 0 11928 2931 11930
rect 0 11872 2870 11928
rect 2926 11872 2931 11928
rect 0 11870 2931 11872
rect 0 11840 480 11870
rect 2865 11867 2931 11870
rect 2497 11794 2563 11797
rect 4889 11794 4955 11797
rect 2497 11792 4955 11794
rect 2497 11736 2502 11792
rect 2558 11736 4894 11792
rect 4950 11736 4955 11792
rect 2497 11734 4955 11736
rect 2497 11731 2563 11734
rect 4889 11731 4955 11734
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 0 11250 480 11280
rect 1761 11250 1827 11253
rect 0 11248 1827 11250
rect 0 11192 1766 11248
rect 1822 11192 1827 11248
rect 0 11190 1827 11192
rect 0 11160 480 11190
rect 1761 11187 1827 11190
rect 7833 11114 7899 11117
rect 19517 11114 19583 11117
rect 7833 11112 19583 11114
rect 7833 11056 7838 11112
rect 7894 11056 19522 11112
rect 19578 11056 19583 11112
rect 7833 11054 19583 11056
rect 7833 11051 7899 11054
rect 19517 11051 19583 11054
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 0 10706 480 10736
rect 3693 10706 3759 10709
rect 0 10704 3759 10706
rect 0 10648 3698 10704
rect 3754 10648 3759 10704
rect 0 10646 3759 10648
rect 0 10616 480 10646
rect 3693 10643 3759 10646
rect 3969 10706 4035 10709
rect 18321 10706 18387 10709
rect 3969 10704 18387 10706
rect 3969 10648 3974 10704
rect 4030 10648 18326 10704
rect 18382 10648 18387 10704
rect 3969 10646 18387 10648
rect 3969 10643 4035 10646
rect 18321 10643 18387 10646
rect 1485 10570 1551 10573
rect 18045 10570 18111 10573
rect 1485 10568 18111 10570
rect 1485 10512 1490 10568
rect 1546 10512 18050 10568
rect 18106 10512 18111 10568
rect 1485 10510 18111 10512
rect 1485 10507 1551 10510
rect 18045 10507 18111 10510
rect 3969 10434 4035 10437
rect 5165 10434 5231 10437
rect 3969 10432 5231 10434
rect 3969 10376 3974 10432
rect 4030 10376 5170 10432
rect 5226 10376 5231 10432
rect 3969 10374 5231 10376
rect 3969 10371 4035 10374
rect 5165 10371 5231 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 6637 10162 6703 10165
rect 19517 10162 19583 10165
rect 6637 10160 19583 10162
rect 6637 10104 6642 10160
rect 6698 10104 19522 10160
rect 19578 10104 19583 10160
rect 6637 10102 19583 10104
rect 6637 10099 6703 10102
rect 19517 10099 19583 10102
rect 0 10026 480 10056
rect 4521 10026 4587 10029
rect 0 10024 4587 10026
rect 0 9968 4526 10024
rect 4582 9968 4587 10024
rect 0 9966 4587 9968
rect 0 9936 480 9966
rect 4521 9963 4587 9966
rect 4705 10026 4771 10029
rect 7741 10026 7807 10029
rect 4705 10024 7807 10026
rect 4705 9968 4710 10024
rect 4766 9968 7746 10024
rect 7802 9968 7807 10024
rect 4705 9966 7807 9968
rect 4705 9963 4771 9966
rect 7741 9963 7807 9966
rect 9673 10026 9739 10029
rect 20897 10026 20963 10029
rect 9673 10024 20963 10026
rect 9673 9968 9678 10024
rect 9734 9968 20902 10024
rect 20958 9968 20963 10024
rect 9673 9966 20963 9968
rect 9673 9963 9739 9966
rect 20897 9963 20963 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 4337 9754 4403 9757
rect 3374 9752 4403 9754
rect 3374 9696 4342 9752
rect 4398 9696 4403 9752
rect 3374 9694 4403 9696
rect 2773 9618 2839 9621
rect 3049 9618 3115 9621
rect 3374 9620 3434 9694
rect 4337 9691 4403 9694
rect 2773 9616 3115 9618
rect 2773 9560 2778 9616
rect 2834 9560 3054 9616
rect 3110 9560 3115 9616
rect 2773 9558 3115 9560
rect 2773 9555 2839 9558
rect 3049 9555 3115 9558
rect 3366 9556 3372 9620
rect 3436 9556 3442 9620
rect 0 9482 480 9512
rect 3233 9482 3299 9485
rect 16665 9482 16731 9485
rect 0 9422 1410 9482
rect 0 9392 480 9422
rect 1350 9346 1410 9422
rect 3233 9480 16731 9482
rect 3233 9424 3238 9480
rect 3294 9424 16670 9480
rect 16726 9424 16731 9480
rect 3233 9422 16731 9424
rect 3233 9419 3299 9422
rect 16665 9419 16731 9422
rect 7649 9346 7715 9349
rect 1350 9344 7715 9346
rect 1350 9288 7654 9344
rect 7710 9288 7715 9344
rect 1350 9286 7715 9288
rect 7649 9283 7715 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 9765 8938 9831 8941
rect 4846 8936 9831 8938
rect 4846 8880 9770 8936
rect 9826 8880 9831 8936
rect 4846 8878 9831 8880
rect 0 8802 480 8832
rect 4846 8802 4906 8878
rect 9765 8875 9831 8878
rect 0 8742 4906 8802
rect 0 8712 480 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 2589 8530 2655 8533
rect 10961 8530 11027 8533
rect 2589 8528 11027 8530
rect 2589 8472 2594 8528
rect 2650 8472 10966 8528
rect 11022 8472 11027 8528
rect 2589 8470 11027 8472
rect 2589 8467 2655 8470
rect 10961 8467 11027 8470
rect 0 8258 480 8288
rect 0 8198 2514 8258
rect 0 8168 480 8198
rect 2454 7986 2514 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 10777 7986 10843 7989
rect 2454 7984 10843 7986
rect 2454 7928 10782 7984
rect 10838 7928 10843 7984
rect 2454 7926 10843 7928
rect 10777 7923 10843 7926
rect 4061 7850 4127 7853
rect 17401 7850 17467 7853
rect 4061 7848 17467 7850
rect 4061 7792 4066 7848
rect 4122 7792 17406 7848
rect 17462 7792 17467 7848
rect 4061 7790 17467 7792
rect 4061 7787 4127 7790
rect 17401 7787 17467 7790
rect 5610 7648 5930 7649
rect 0 7578 480 7608
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 0 7518 1410 7578
rect 0 7488 480 7518
rect 1350 7306 1410 7518
rect 22185 7306 22251 7309
rect 1350 7304 22251 7306
rect 1350 7248 22190 7304
rect 22246 7248 22251 7304
rect 1350 7246 22251 7248
rect 22185 7243 22251 7246
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 0 6974 2698 7034
rect 0 6944 480 6974
rect 2638 6898 2698 6974
rect 22737 6898 22803 6901
rect 2638 6896 22803 6898
rect 2638 6840 22742 6896
rect 22798 6840 22803 6896
rect 2638 6838 22803 6840
rect 22737 6835 22803 6838
rect 3417 6762 3483 6765
rect 7925 6762 7991 6765
rect 3417 6760 7991 6762
rect 3417 6704 3422 6760
rect 3478 6704 7930 6760
rect 7986 6704 7991 6760
rect 3417 6702 7991 6704
rect 3417 6699 3483 6702
rect 7925 6699 7991 6702
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 23657 6354 23723 6357
rect 0 6352 23723 6354
rect 0 6296 23662 6352
rect 23718 6296 23723 6352
rect 0 6294 23723 6296
rect 0 6264 480 6294
rect 23657 6291 23723 6294
rect 2957 6218 3023 6221
rect 9029 6218 9095 6221
rect 2957 6216 9095 6218
rect 2957 6160 2962 6216
rect 3018 6160 9034 6216
rect 9090 6160 9095 6216
rect 2957 6158 9095 6160
rect 2957 6155 3023 6158
rect 9029 6155 9095 6158
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 0 5810 480 5840
rect 23933 5810 23999 5813
rect 0 5808 23999 5810
rect 0 5752 23938 5808
rect 23994 5752 23999 5808
rect 0 5750 23999 5752
rect 0 5720 480 5750
rect 23933 5747 23999 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 24485 5266 24551 5269
rect 2638 5264 24551 5266
rect 2638 5208 24490 5264
rect 24546 5208 24551 5264
rect 2638 5206 24551 5208
rect 0 5130 480 5160
rect 2638 5130 2698 5206
rect 24485 5203 24551 5206
rect 0 5070 2698 5130
rect 0 5040 480 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24761 4858 24827 4861
rect 26325 4858 26391 4861
rect 24761 4856 26391 4858
rect 24761 4800 24766 4856
rect 24822 4800 26330 4856
rect 26386 4800 26391 4856
rect 24761 4798 26391 4800
rect 24761 4795 24827 4798
rect 26325 4795 26391 4798
rect 24577 4722 24643 4725
rect 2638 4720 24643 4722
rect 2638 4664 24582 4720
rect 24638 4664 24643 4720
rect 2638 4662 24643 4664
rect 0 4586 480 4616
rect 2638 4586 2698 4662
rect 24577 4659 24643 4662
rect 0 4526 2698 4586
rect 0 4496 480 4526
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 0 3906 480 3936
rect 3877 3906 3943 3909
rect 0 3904 3943 3906
rect 0 3848 3882 3904
rect 3938 3848 3943 3904
rect 0 3846 3943 3848
rect 0 3816 480 3846
rect 3877 3843 3943 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 5441 3498 5507 3501
rect 20989 3498 21055 3501
rect 5441 3496 21055 3498
rect 5441 3440 5446 3496
rect 5502 3440 20994 3496
rect 21050 3440 21055 3496
rect 5441 3438 21055 3440
rect 5441 3435 5507 3438
rect 20989 3435 21055 3438
rect 0 3362 480 3392
rect 3325 3362 3391 3365
rect 0 3360 3391 3362
rect 0 3304 3330 3360
rect 3386 3304 3391 3360
rect 0 3302 3391 3304
rect 0 3272 480 3302
rect 3325 3299 3391 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2589 2682 2655 2685
rect 0 2680 2655 2682
rect 0 2624 2594 2680
rect 2650 2624 2655 2680
rect 0 2622 2655 2624
rect 0 2592 480 2622
rect 2589 2619 2655 2622
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 3366 2138 3372 2140
rect 0 2078 3372 2138
rect 0 2048 480 2078
rect 3366 2076 3372 2078
rect 3436 2076 3442 2140
rect 0 1458 480 1488
rect 3417 1458 3483 1461
rect 0 1456 3483 1458
rect 0 1400 3422 1456
rect 3478 1400 3483 1456
rect 0 1398 3483 1400
rect 0 1368 480 1398
rect 3417 1395 3483 1398
rect 12617 1322 12683 1325
rect 3190 1320 12683 1322
rect 3190 1264 12622 1320
rect 12678 1264 12683 1320
rect 3190 1262 12683 1264
rect 0 914 480 944
rect 3190 914 3250 1262
rect 12617 1259 12683 1262
rect 0 854 3250 914
rect 0 824 480 854
rect 0 370 480 400
rect 2957 370 3023 373
rect 0 368 3023 370
rect 0 312 2962 368
rect 3018 312 3023 368
rect 0 310 3023 312
rect 0 280 480 310
rect 2957 307 3023 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 9996 19076 10060 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 9996 18532 10060 18596
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 3372 9556 3436 9620
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 3372 2076 3436 2140
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9995 19140 10061 19141
rect 9995 19076 9996 19140
rect 10060 19076 10061 19140
rect 9995 19075 10061 19076
rect 9998 18597 10058 19075
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 9995 18596 10061 18597
rect 9995 18532 9996 18596
rect 10060 18532 10061 18596
rect 9995 18531 10061 18532
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 3374 2141 3434 9555
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 3371 2140 3437 2141
rect 3371 2076 3372 2140
rect 3436 2076 3437 2140
rect 5610 2128 5931 2144
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 3371 2075 3437 2076
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604681595
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_273
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24564 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_251
timestamp 1604681595
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1604681595
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1604681595
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1604681595
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_250
timestamp 1604681595
transform 1 0 24104 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_262
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_274
timestamp 1604681595
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_237
timestamp 1604681595
transform 1 0 22908 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__84__A
timestamp 1604681595
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1604681595
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1604681595
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 23920 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__83__A
timestamp 1604681595
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_252
timestamp 1604681595
transform 1 0 24288 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_264
timestamp 1604681595
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_272
timestamp 1604681595
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604681595
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_11
timestamp 1604681595
transform 1 0 2116 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_16
timestamp 1604681595
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1604681595
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4048 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp 1604681595
transform 1 0 3312 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_34
timestamp 1604681595
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_38
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_54
timestamp 1604681595
transform 1 0 6072 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1604681595
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_228
timestamp 1604681595
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1604681595
transform 1 0 22724 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1604681595
transform 1 0 22540 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1604681595
transform 1 0 22908 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1604681595
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_13
timestamp 1604681595
transform 1 0 2300 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1604681595
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp 1604681595
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1604681595
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1604681595
transform 1 0 5980 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1604681595
transform 1 0 7084 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_77
timestamp 1604681595
transform 1 0 8188 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604681595
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 1564 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_8
timestamp 1604681595
transform 1 0 1840 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_17
timestamp 1604681595
transform 1 0 2668 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_29
timestamp 1604681595
transform 1 0 3772 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1604681595
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_73
timestamp 1604681595
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_77
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_89
timestamp 1604681595
transform 1 0 9292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_101
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1604681595
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604681595
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_269
timestamp 1604681595
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_20
timestamp 1604681595
transform 1 0 2944 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1604681595
transform 1 0 3312 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_28
timestamp 1604681595
transform 1 0 3680 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_35
timestamp 1604681595
transform 1 0 4324 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5060 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_76
timestamp 1604681595
transform 1 0 8096 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1604681595
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1840 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_24
timestamp 1604681595
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_41
timestamp 1604681595
transform 1 0 4876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_14_49
timestamp 1604681595
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_45
timestamp 1604681595
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1604681595
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1604681595
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1604681595
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5980 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7084 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_79
timestamp 1604681595
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_85
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_103
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_115
timestamp 1604681595
transform 1 0 11684 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_121
timestamp 1604681595
transform 1 0 12236 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_106
timestamp 1604681595
transform 1 0 10856 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_118
timestamp 1604681595
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_130
timestamp 1604681595
transform 1 0 13064 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1604681595
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1604681595
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1604681595
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1604681595
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1604681595
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1472 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1604681595
transform 1 0 2300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_17
timestamp 1604681595
transform 1 0 2668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 1604681595
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_25
timestamp 1604681595
transform 1 0 3404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5612 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_47
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_51
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_55
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1604681595
transform 1 0 7452 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10396 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_97
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1604681595
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19596 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604681595
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1604681595
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1604681595
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_223
timestamp 1604681595
transform 1 0 21620 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_235
timestamp 1604681595
transform 1 0 22724 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1604681595
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1604681595
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604681595
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_46
timestamp 1604681595
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_70
timestamp 1604681595
transform 1 0 7544 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1604681595
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_113
timestamp 1604681595
transform 1 0 11500 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_137
timestamp 1604681595
transform 1 0 13708 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1604681595
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1604681595
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1604681595
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1604681595
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_12
timestamp 1604681595
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1604681595
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp 1604681595
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1604681595
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_111
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_119
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_152
timestamp 1604681595
transform 1 0 15088 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_164
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1604681595
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_190
timestamp 1604681595
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_194
timestamp 1604681595
transform 1 0 18952 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_206
timestamp 1604681595
transform 1 0 20056 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_214
timestamp 1604681595
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1604681595
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_50
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8096 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1604681595
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_81
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1604681595
transform 1 0 9200 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1604681595
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_139
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1604681595
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1604681595
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_257
timestamp 1604681595
transform 1 0 24748 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 1932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1604681595
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1604681595
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1604681595
transform 1 0 2116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_35
timestamp 1604681595
transform 1 0 4324 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1604681595
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1604681595
transform 1 0 4968 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_59
timestamp 1604681595
transform 1 0 6532 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8280 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_78
timestamp 1604681595
transform 1 0 8280 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_82
timestamp 1604681595
transform 1 0 8648 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_64
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_76
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_80
timestamp 1604681595
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_99
timestamp 1604681595
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1604681595
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_110
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_120
timestamp 1604681595
transform 1 0 12144 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_116
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_139
timestamp 1604681595
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1604681595
transform 1 0 16376 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1604681595
transform 1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_183
timestamp 1604681595
transform 1 0 17940 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_195
timestamp 1604681595
transform 1 0 19044 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1604681595
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1604681595
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1604681595
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1604681595
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1604681595
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1604681595
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_32
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1604681595
transform 1 0 11224 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1604681595
transform 1 0 10856 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1604681595
transform 1 0 11500 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_150
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_168
timestamp 1604681595
transform 1 0 16560 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_19
timestamp 1604681595
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3496 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6164 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_53
timestamp 1604681595
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 7728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_68
timestamp 1604681595
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1604681595
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1604681595
transform 1 0 13340 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1604681595
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_144
timestamp 1604681595
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1604681595
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1604681595
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1604681595
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1604681595
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_12
timestamp 1604681595
transform 1 0 2208 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_31
timestamp 1604681595
transform 1 0 3956 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_52
timestamp 1604681595
transform 1 0 5888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1604681595
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_165
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_177
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_6
timestamp 1604681595
transform 1 0 1656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_10
timestamp 1604681595
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604681595
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1604681595
transform 1 0 5244 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8004 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_66
timestamp 1604681595
transform 1 0 7176 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_70
timestamp 1604681595
transform 1 0 7544 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_73
timestamp 1604681595
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_77
timestamp 1604681595
transform 1 0 8188 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_115
timestamp 1604681595
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1604681595
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_139
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_143
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16100 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_162
timestamp 1604681595
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_169
timestamp 1604681595
transform 1 0 16652 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_181
timestamp 1604681595
transform 1 0 17756 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1604681595
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1604681595
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1604681595
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1604681595
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1564 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_14
timestamp 1604681595
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 3128 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_46
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 5704 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_83
timestamp 1604681595
transform 1 0 8740 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9108 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1604681595
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_166
timestamp 1604681595
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1604681595
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1604681595
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_269
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_35
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_50
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_46
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 5152 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5888 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_87
timestamp 1604681595
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1604681595
transform 1 0 11500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_113
timestamp 1604681595
transform 1 0 11500 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1604681595
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1604681595
transform 1 0 12236 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_117
timestamp 1604681595
transform 1 0 11868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_123
timestamp 1604681595
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12052 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 11684 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp 1604681595
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1604681595
transform 1 0 12788 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1604681595
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_140
timestamp 1604681595
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1604681595
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_160
timestamp 1604681595
transform 1 0 15824 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1604681595
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_155
timestamp 1604681595
transform 1 0 15364 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_172
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_184
timestamp 1604681595
transform 1 0 18032 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_167
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1604681595
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1604681595
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1604681595
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1604681595
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_269
timestamp 1604681595
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1604681595
transform 1 0 1656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1604681595
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4600 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1604681595
transform 1 0 4416 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_40
timestamp 1604681595
transform 1 0 4784 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 6900 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_79
timestamp 1604681595
transform 1 0 8372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_83
timestamp 1604681595
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_87
timestamp 1604681595
transform 1 0 9108 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_106
timestamp 1604681595
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_130
timestamp 1604681595
transform 1 0 13064 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_134
timestamp 1604681595
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_144
timestamp 1604681595
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1604681595
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1604681595
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1604681595
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1604681595
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1604681595
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1604681595
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1656 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_22
timestamp 1604681595
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_26
timestamp 1604681595
transform 1 0 3496 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_46
timestamp 1604681595
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_50
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_54
timestamp 1604681595
transform 1 0 6072 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1604681595
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1604681595
transform 1 0 9568 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12880 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_148
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_160
timestamp 1604681595
transform 1 0 15824 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1604681595
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1604681595
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_269
timestamp 1604681595
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_6
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_40
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5520 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_72
timestamp 1604681595
transform 1 0 7728 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_77
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1604681595
transform 1 0 12328 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1604681595
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_139
timestamp 1604681595
transform 1 0 13892 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1604681595
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_29
timestamp 1604681595
transform 1 0 3772 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_99
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_116
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_143
timestamp 1604681595
transform 1 0 14260 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 1604681595
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_160
timestamp 1604681595
transform 1 0 15824 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1604681595
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604681595
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 1564 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3312 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_26
timestamp 1604681595
transform 1 0 3496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1604681595
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1604681595
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 7360 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1604681595
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_120
timestamp 1604681595
transform 1 0 12144 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_137
timestamp 1604681595
transform 1 0 13708 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_160
timestamp 1604681595
transform 1 0 15824 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_172
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_196
timestamp 1604681595
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_208
timestamp 1604681595
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1604681595
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1604681595
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_6
timestamp 1604681595
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_16
timestamp 1604681595
transform 1 0 2576 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_12
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_10
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 2944 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_23
timestamp 1604681595
transform 1 0 3220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_38
timestamp 1604681595
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_34
timestamp 1604681595
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_52
timestamp 1604681595
transform 1 0 5888 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_48
timestamp 1604681595
transform 1 0 5520 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 5704 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_55
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6716 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_78
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1604681595
transform 1 0 8648 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_77
timestamp 1604681595
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_81
timestamp 1604681595
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10672 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_102
timestamp 1604681595
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1604681595
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_109
timestamp 1604681595
transform 1 0 11132 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1604681595
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_113
timestamp 1604681595
transform 1 0 11500 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1604681595
transform 1 0 11500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11316 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_121
timestamp 1604681595
transform 1 0 12236 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13064 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_127
timestamp 1604681595
transform 1 0 12788 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1604681595
transform 1 0 14812 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1604681595
transform 1 0 14904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_146
timestamp 1604681595
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 15272 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_157
timestamp 1604681595
transform 1 0 15548 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1604681595
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1604681595
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_220
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604681595
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604681595
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_11
timestamp 1604681595
transform 1 0 2116 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 4140 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_25
timestamp 1604681595
transform 1 0 3404 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_29
timestamp 1604681595
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_37
timestamp 1604681595
transform 1 0 4508 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_42
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 5244 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_49
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_53
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1604681595
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8740 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_66
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_79
timestamp 1604681595
transform 1 0 8372 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9292 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10304 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_85
timestamp 1604681595
transform 1 0 8924 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_102
timestamp 1604681595
transform 1 0 10488 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604681595
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14076 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_133
timestamp 1604681595
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 15640 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15088 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1604681595
transform 1 0 14904 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_154
timestamp 1604681595
transform 1 0 15272 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_161
timestamp 1604681595
transform 1 0 15916 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_173
timestamp 1604681595
transform 1 0 17020 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_181
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1604681595
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1604681595
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1604681595
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1604681595
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1604681595
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1604681595
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 2852 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_11
timestamp 1604681595
transform 1 0 2116 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 5704 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 6072 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1604681595
transform 1 0 5888 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_56
timestamp 1604681595
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7912 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_67
timestamp 1604681595
transform 1 0 7268 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_72
timestamp 1604681595
transform 1 0 7728 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_76
timestamp 1604681595
transform 1 0 8096 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9936 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_84
timestamp 1604681595
transform 1 0 8832 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_88
timestamp 1604681595
transform 1 0 9200 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_91
timestamp 1604681595
transform 1 0 9476 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 12144 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 11960 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_112
timestamp 1604681595
transform 1 0 11408 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_123
timestamp 1604681595
transform 1 0 12420 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12972 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_157
timestamp 1604681595
transform 1 0 15548 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1604681595
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1604681595
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_192
timestamp 1604681595
transform 1 0 18768 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_204
timestamp 1604681595
transform 1 0 19872 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1604681595
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1604681595
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1604681595
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_263
timestamp 1604681595
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2668 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_10
timestamp 1604681595
transform 1 0 2024 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_19
timestamp 1604681595
transform 1 0 2852 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3220 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_32
timestamp 1604681595
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1604681595
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 6348 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_49
timestamp 1604681595
transform 1 0 5612 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1604681595
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7084 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8280 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_76
timestamp 1604681595
transform 1 0 8096 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_80
timestamp 1604681595
transform 1 0 8464 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9200 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1604681595
transform 1 0 8832 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_103
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_107
timestamp 1604681595
transform 1 0 10948 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13064 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1604681595
transform 1 0 12788 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15732 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14720 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_146
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_150
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_157
timestamp 1604681595
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1604681595
transform 1 0 15916 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__95__A
timestamp 1604681595
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1604681595
transform 1 0 16468 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_170
timestamp 1604681595
transform 1 0 16744 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_182
timestamp 1604681595
transform 1 0 17848 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__90__A
timestamp 1604681595
transform 1 0 19320 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_196
timestamp 1604681595
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_200
timestamp 1604681595
transform 1 0 19504 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_212
timestamp 1604681595
transform 1 0 20608 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_217
timestamp 1604681595
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1604681595
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_241
timestamp 1604681595
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1604681595
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_269
timestamp 1604681595
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 2852 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1564 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2300 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1604681595
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604681595
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_48
timestamp 1604681595
transform 1 0 5520 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_59
timestamp 1604681595
transform 1 0 6532 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6900 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_81
timestamp 1604681595
transform 1 0 8556 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1604681595
transform 1 0 8924 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11868 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_111
timestamp 1604681595
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_115
timestamp 1604681595
transform 1 0 11684 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_119
timestamp 1604681595
transform 1 0 12052 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_124
timestamp 1604681595
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12880 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_144
timestamp 1604681595
transform 1 0 14352 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_152
timestamp 1604681595
transform 1 0 15088 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_160
timestamp 1604681595
transform 1 0 15824 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _95_
timestamp 1604681595
transform 1 0 16560 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_172
timestamp 1604681595
transform 1 0 16928 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_184
timestamp 1604681595
transform 1 0 18032 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 19320 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_196
timestamp 1604681595
transform 1 0 19136 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1604681595
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_221
timestamp 1604681595
transform 1 0 21436 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_233
timestamp 1604681595
transform 1 0 22540 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_245
timestamp 1604681595
transform 1 0 23644 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_257
timestamp 1604681595
transform 1 0 24748 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_269
timestamp 1604681595
transform 1 0 25852 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1656 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_10
timestamp 1604681595
transform 1 0 2024 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_12
timestamp 1604681595
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_17
timestamp 1604681595
transform 1 0 2668 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_14
timestamp 1604681595
transform 1 0 2392 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_20
timestamp 1604681595
transform 1 0 2944 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_16
timestamp 1604681595
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 2760 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 2760 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1604681595
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_26
timestamp 1604681595
transform 1 0 3496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_22
timestamp 1604681595
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3128 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_40
timestamp 1604681595
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3312 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4692 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_44
timestamp 1604681595
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 5336 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 5520 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_55
timestamp 1604681595
transform 1 0 6164 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_52
timestamp 1604681595
transform 1 0 5888 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_60
timestamp 1604681595
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6808 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6992 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7084 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 8648 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_80
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 9016 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_85
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_89
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_88
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_93
timestamp 1604681595
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9936 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10028 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_40_109
timestamp 1604681595
transform 1 0 11132 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1604681595
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 10948 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11500 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_122
timestamp 1604681595
transform 1 0 12328 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_117
timestamp 1604681595
transform 1 0 11868 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12880 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13064 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12696 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12880 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_144
timestamp 1604681595
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_126
timestamp 1604681595
transform 1 0 12696 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_139
timestamp 1604681595
transform 1 0 13892 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_148
timestamp 1604681595
transform 1 0 14720 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _99_
timestamp 1604681595
transform 1 0 15088 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _98_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1604681595
transform 1 0 15640 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_160
timestamp 1604681595
transform 1 0 15824 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_156
timestamp 1604681595
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__98__A
timestamp 1604681595
transform 1 0 16008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__99__A
timestamp 1604681595
transform 1 0 15640 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _97_
timestamp 1604681595
transform 1 0 16192 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _96_
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_170
timestamp 1604681595
transform 1 0 16744 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_172
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_168
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__96__A
timestamp 1604681595
transform 1 0 17112 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__97__A
timestamp 1604681595
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_182
timestamp 1604681595
transform 1 0 17848 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_180
timestamp 1604681595
transform 1 0 17664 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_176
timestamp 1604681595
transform 1 0 17296 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__94__A
timestamp 1604681595
transform 1 0 17480 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _94_
timestamp 1604681595
transform 1 0 17480 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _93_
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_190
timestamp 1604681595
transform 1 0 18584 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1604681595
transform 1 0 18768 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_188
timestamp 1604681595
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__91__A
timestamp 1604681595
transform 1 0 18952 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__93__A
timestamp 1604681595
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _92_
timestamp 1604681595
transform 1 0 19136 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _91_
timestamp 1604681595
transform 1 0 18768 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_208
timestamp 1604681595
transform 1 0 20240 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1604681595
transform 1 0 19504 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__92__A
timestamp 1604681595
transform 1 0 19688 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_196
timestamp 1604681595
transform 1 0 19136 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_216
timestamp 1604681595
transform 1 0 20976 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_212
timestamp 1604681595
transform 1 0 20608 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__88__A
timestamp 1604681595
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__89__A
timestamp 1604681595
transform 1 0 20792 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__87__A
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 21344 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_219
timestamp 1604681595
transform 1 0 21252 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__86__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_231
timestamp 1604681595
transform 1 0 22356 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_269
timestamp 1604681595
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_255
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_267
timestamp 1604681595
transform 1 0 25668 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2944 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4876 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_39
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_43
timestamp 1604681595
transform 1 0 5060 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_53
timestamp 1604681595
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 8372 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8188 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_71
timestamp 1604681595
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_75
timestamp 1604681595
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_83
timestamp 1604681595
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_87
timestamp 1604681595
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_91
timestamp 1604681595
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_104
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_108
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 13984 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_132
timestamp 1604681595
transform 1 0 13248 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_155
timestamp 1604681595
transform 1 0 15364 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_167
timestamp 1604681595
transform 1 0 16468 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_179
timestamp 1604681595
transform 1 0 17572 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1604681595
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1604681595
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1604681595
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1604681595
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1604681595
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_269
timestamp 1604681595
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3128 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_24
timestamp 1604681595
transform 1 0 3312 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1604681595
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_32
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5888 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_46
timestamp 1604681595
transform 1 0 5336 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_50
timestamp 1604681595
transform 1 0 5704 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_54
timestamp 1604681595
transform 1 0 6072 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 8464 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_72
timestamp 1604681595
transform 1 0 7728 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_84
timestamp 1604681595
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_92
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_98
timestamp 1604681595
transform 1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_102
timestamp 1604681595
transform 1 0 10488 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 10856 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_110
timestamp 1604681595
transform 1 0 11224 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_122
timestamp 1604681595
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 13616 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_128
timestamp 1604681595
transform 1 0 12880 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_139
timestamp 1604681595
transform 1 0 13892 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_180
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_187
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_199
timestamp 1604681595
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_211
timestamp 1604681595
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1604681595
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_242
timestamp 1604681595
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604681595
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604681595
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 14016 28000 14136 6 ccff_head
port 0 nsew default input
rlabel metal2 s 20994 0 21050 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 4802 27520 4858 28000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 10506 27520 10562 28000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 11058 27520 11114 28000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 11702 27520 11758 28000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 12254 27520 12310 28000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 12806 27520 12862 28000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 13358 27520 13414 28000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14554 27520 14610 28000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15106 27520 15162 28000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15658 27520 15714 28000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 5354 27520 5410 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 5998 27520 6054 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 6550 27520 6606 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 7102 27520 7158 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 8206 27520 8262 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8850 27520 8906 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9402 27520 9458 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 9954 27520 10010 28000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 16210 27520 16266 28000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 21914 27520 21970 28000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 22466 27520 22522 28000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 23110 27520 23166 28000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 23662 27520 23718 28000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 24214 27520 24270 28000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 16762 27520 16818 28000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 17406 27520 17462 28000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 17958 27520 18014 28000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 18510 27520 18566 28000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 19614 27520 19670 28000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 20258 27520 20314 28000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 20810 27520 20866 28000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 21362 27520 21418 28000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 84 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 85 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 86 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 87 nsew default input
rlabel metal2 s 7010 0 7066 480 6 prog_clk
port 88 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_42_
port 89 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_43_
port 90 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_44_
port 91 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_45_
port 92 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_46_
port 93 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_47_
port 94 nsew default input
rlabel metal2 s 3698 27520 3754 28000 6 top_left_grid_pin_48_
port 95 nsew default input
rlabel metal2 s 4250 27520 4306 28000 6 top_left_grid_pin_49_
port 96 nsew default input
rlabel metal2 s 27618 27520 27674 28000 6 top_right_grid_pin_1_
port 97 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 98 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 99 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
