VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cbx_1__0_
  CLASS BLOCK ;
  FOREIGN cbx_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 120.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 2.400 ;
    END
  END SC_IN_BOT
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 117.600 48.670 120.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 2.400 ;
    END
  END SC_OUT_BOT
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.210 117.600 56.490 120.000 ;
    END
  END SC_OUT_TOP
  PIN bottom_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END bottom_grid_pin_0_
  PIN bottom_grid_pin_10_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 2.400 ;
    END
  END bottom_grid_pin_10_
  PIN bottom_grid_pin_2_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END bottom_grid_pin_2_
  PIN bottom_grid_pin_4_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 2.400 ;
    END
  END bottom_grid_pin_4_
  PIN bottom_grid_pin_6_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 2.400 ;
    END
  END bottom_grid_pin_6_
  PIN bottom_grid_pin_8_
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END bottom_grid_pin_8_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 2.400 97.200 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 2.400 106.720 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 2.400 109.440 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 2.400 112.160 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 2.400 118.280 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 2.400 67.280 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 2.400 76.800 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 2.400 79.520 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 2.400 82.240 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 2.400 85.640 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 2.400 88.360 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 2.400 2.000 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 2.400 34.640 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 2.400 37.360 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 2.400 43.480 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 2.400 46.880 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 2.400 49.600 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 2.400 55.720 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 2.400 58.440 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 2.400 4.720 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 2.400 7.440 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 2.400 13.560 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 2.400 16.960 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 2.400 22.400 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 2.400 25.800 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 2.400 28.520 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 61.240 150.000 61.840 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 91.160 150.000 91.760 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 93.880 150.000 94.480 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 96.600 150.000 97.200 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 100.000 150.000 100.600 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 102.720 150.000 103.320 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 106.120 150.000 106.720 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 108.840 150.000 109.440 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 111.560 150.000 112.160 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 114.960 150.000 115.560 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 117.680 150.000 118.280 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 63.960 150.000 64.560 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 66.680 150.000 67.280 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 70.080 150.000 70.680 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 72.800 150.000 73.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 76.200 150.000 76.800 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 78.920 150.000 79.520 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 81.640 150.000 82.240 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 85.040 150.000 85.640 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 147.600 87.760 150.000 88.360 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 1.400 150.000 2.000 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 31.320 150.000 31.920 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 34.040 150.000 34.640 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 36.760 150.000 37.360 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 40.160 150.000 40.760 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 42.880 150.000 43.480 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 46.280 150.000 46.880 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 49.000 150.000 49.600 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 51.720 150.000 52.320 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 55.120 150.000 55.720 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 57.840 150.000 58.440 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 4.120 150.000 4.720 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 6.840 150.000 7.440 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 10.240 150.000 10.840 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 12.960 150.000 13.560 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 16.360 150.000 16.960 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 19.080 150.000 19.680 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 21.800 150.000 22.400 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 25.200 150.000 25.800 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 147.600 27.920 150.000 28.520 ;
    END
  END chanx_right_out[9]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_DIR[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_IN[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_IN[5]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[0]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[1]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[2]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[3]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[4]
  PIN gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 2.400 ;
    END
  END gfpga_pad_EMBEDDED_IO_SOC_OUT[5]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 2.400 ;
    END
  END prog_clk
  PIN top_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 117.600 63.850 120.000 ;
    END
  END top_width_0_height_0__pin_0_
  PIN top_width_0_height_0__pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 117.600 101.110 120.000 ;
    END
  END top_width_0_height_0__pin_10_
  PIN top_width_0_height_0__pin_11_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 145.910 117.600 146.190 120.000 ;
    END
  END top_width_0_height_0__pin_11_lower
  PIN top_width_0_height_0__pin_11_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.030 117.600 41.310 120.000 ;
    END
  END top_width_0_height_0__pin_11_upper
  PIN top_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 117.600 108.930 120.000 ;
    END
  END top_width_0_height_0__pin_1_lower
  PIN top_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 3.770 117.600 4.050 120.000 ;
    END
  END top_width_0_height_0__pin_1_upper
  PIN top_width_0_height_0__pin_2_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.930 117.600 71.210 120.000 ;
    END
  END top_width_0_height_0__pin_2_
  PIN top_width_0_height_0__pin_3_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 117.600 116.290 120.000 ;
    END
  END top_width_0_height_0__pin_3_lower
  PIN top_width_0_height_0__pin_3_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.130 117.600 11.410 120.000 ;
    END
  END top_width_0_height_0__pin_3_upper
  PIN top_width_0_height_0__pin_4_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.750 117.600 79.030 120.000 ;
    END
  END top_width_0_height_0__pin_4_
  PIN top_width_0_height_0__pin_5_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 123.370 117.600 123.650 120.000 ;
    END
  END top_width_0_height_0__pin_5_lower
  PIN top_width_0_height_0__pin_5_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.490 117.600 18.770 120.000 ;
    END
  END top_width_0_height_0__pin_5_upper
  PIN top_width_0_height_0__pin_6_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.110 117.600 86.390 120.000 ;
    END
  END top_width_0_height_0__pin_6_
  PIN top_width_0_height_0__pin_7_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 117.600 131.470 120.000 ;
    END
  END top_width_0_height_0__pin_7_lower
  PIN top_width_0_height_0__pin_7_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 117.600 26.130 120.000 ;
    END
  END top_width_0_height_0__pin_7_upper
  PIN top_width_0_height_0__pin_8_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.470 117.600 93.750 120.000 ;
    END
  END top_width_0_height_0__pin_8_
  PIN top_width_0_height_0__pin_9_lower
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.550 117.600 138.830 120.000 ;
    END
  END top_width_0_height_0__pin_9_lower
  PIN top_width_0_height_0__pin_9_upper
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.670 117.600 33.950 120.000 ;
    END
  END top_width_0_height_0__pin_9_upper
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.720 10.640 31.320 109.040 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 54.720 10.640 56.320 109.040 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 108.885 ;
      LAYER met1 ;
        RECT 5.520 2.760 144.440 111.140 ;
      LAYER met2 ;
        RECT 2.460 117.320 3.490 118.165 ;
        RECT 4.330 117.320 10.850 118.165 ;
        RECT 11.690 117.320 18.210 118.165 ;
        RECT 19.050 117.320 25.570 118.165 ;
        RECT 26.410 117.320 33.390 118.165 ;
        RECT 34.230 117.320 40.750 118.165 ;
        RECT 41.590 117.320 48.110 118.165 ;
        RECT 48.950 117.320 55.930 118.165 ;
        RECT 56.770 117.320 63.290 118.165 ;
        RECT 64.130 117.320 70.650 118.165 ;
        RECT 71.490 117.320 78.470 118.165 ;
        RECT 79.310 117.320 85.830 118.165 ;
        RECT 86.670 117.320 93.190 118.165 ;
        RECT 94.030 117.320 100.550 118.165 ;
        RECT 101.390 117.320 108.370 118.165 ;
        RECT 109.210 117.320 115.730 118.165 ;
        RECT 116.570 117.320 123.090 118.165 ;
        RECT 123.930 117.320 130.910 118.165 ;
        RECT 131.750 117.320 138.270 118.165 ;
        RECT 139.110 117.320 145.630 118.165 ;
        RECT 146.470 117.320 147.110 118.165 ;
        RECT 2.460 2.680 147.110 117.320 ;
        RECT 2.950 1.515 7.170 2.680 ;
        RECT 8.010 1.515 12.230 2.680 ;
        RECT 13.070 1.515 17.290 2.680 ;
        RECT 18.130 1.515 22.350 2.680 ;
        RECT 23.190 1.515 27.870 2.680 ;
        RECT 28.710 1.515 32.930 2.680 ;
        RECT 33.770 1.515 37.990 2.680 ;
        RECT 38.830 1.515 43.050 2.680 ;
        RECT 43.890 1.515 48.570 2.680 ;
        RECT 49.410 1.515 53.630 2.680 ;
        RECT 54.470 1.515 58.690 2.680 ;
        RECT 59.530 1.515 63.750 2.680 ;
        RECT 64.590 1.515 69.270 2.680 ;
        RECT 70.110 1.515 74.330 2.680 ;
        RECT 75.170 1.515 79.390 2.680 ;
        RECT 80.230 1.515 84.450 2.680 ;
        RECT 85.290 1.515 89.970 2.680 ;
        RECT 90.810 1.515 95.030 2.680 ;
        RECT 95.870 1.515 100.090 2.680 ;
        RECT 100.930 1.515 105.150 2.680 ;
        RECT 105.990 1.515 110.670 2.680 ;
        RECT 111.510 1.515 115.730 2.680 ;
        RECT 116.570 1.515 120.790 2.680 ;
        RECT 121.630 1.515 125.850 2.680 ;
        RECT 126.690 1.515 131.370 2.680 ;
        RECT 132.210 1.515 136.430 2.680 ;
        RECT 137.270 1.515 141.490 2.680 ;
        RECT 142.330 1.515 146.550 2.680 ;
      LAYER met3 ;
        RECT 2.800 117.280 147.200 118.145 ;
        RECT 2.400 115.960 147.600 117.280 ;
        RECT 2.800 114.560 147.200 115.960 ;
        RECT 2.400 112.560 147.600 114.560 ;
        RECT 2.800 111.160 147.200 112.560 ;
        RECT 2.400 109.840 147.600 111.160 ;
        RECT 2.800 108.440 147.200 109.840 ;
        RECT 2.400 107.120 147.600 108.440 ;
        RECT 2.800 105.720 147.200 107.120 ;
        RECT 2.400 103.720 147.600 105.720 ;
        RECT 2.800 102.320 147.200 103.720 ;
        RECT 2.400 101.000 147.600 102.320 ;
        RECT 2.800 99.600 147.200 101.000 ;
        RECT 2.400 97.600 147.600 99.600 ;
        RECT 2.800 96.200 147.200 97.600 ;
        RECT 2.400 94.880 147.600 96.200 ;
        RECT 2.800 93.480 147.200 94.880 ;
        RECT 2.400 92.160 147.600 93.480 ;
        RECT 2.800 90.760 147.200 92.160 ;
        RECT 2.400 88.760 147.600 90.760 ;
        RECT 2.800 87.360 147.200 88.760 ;
        RECT 2.400 86.040 147.600 87.360 ;
        RECT 2.800 84.640 147.200 86.040 ;
        RECT 2.400 82.640 147.600 84.640 ;
        RECT 2.800 81.240 147.200 82.640 ;
        RECT 2.400 79.920 147.600 81.240 ;
        RECT 2.800 78.520 147.200 79.920 ;
        RECT 2.400 77.200 147.600 78.520 ;
        RECT 2.800 75.800 147.200 77.200 ;
        RECT 2.400 73.800 147.600 75.800 ;
        RECT 2.800 72.400 147.200 73.800 ;
        RECT 2.400 71.080 147.600 72.400 ;
        RECT 2.800 69.680 147.200 71.080 ;
        RECT 2.400 67.680 147.600 69.680 ;
        RECT 2.800 66.280 147.200 67.680 ;
        RECT 2.400 64.960 147.600 66.280 ;
        RECT 2.800 63.560 147.200 64.960 ;
        RECT 2.400 62.240 147.600 63.560 ;
        RECT 2.800 60.840 147.200 62.240 ;
        RECT 2.400 58.840 147.600 60.840 ;
        RECT 2.800 57.440 147.200 58.840 ;
        RECT 2.400 56.120 147.600 57.440 ;
        RECT 2.800 54.720 147.200 56.120 ;
        RECT 2.400 52.720 147.600 54.720 ;
        RECT 2.800 51.320 147.200 52.720 ;
        RECT 2.400 50.000 147.600 51.320 ;
        RECT 2.800 48.600 147.200 50.000 ;
        RECT 2.400 47.280 147.600 48.600 ;
        RECT 2.800 45.880 147.200 47.280 ;
        RECT 2.400 43.880 147.600 45.880 ;
        RECT 2.800 42.480 147.200 43.880 ;
        RECT 2.400 41.160 147.600 42.480 ;
        RECT 2.800 39.760 147.200 41.160 ;
        RECT 2.400 37.760 147.600 39.760 ;
        RECT 2.800 36.360 147.200 37.760 ;
        RECT 2.400 35.040 147.600 36.360 ;
        RECT 2.800 33.640 147.200 35.040 ;
        RECT 2.400 32.320 147.600 33.640 ;
        RECT 2.800 30.920 147.200 32.320 ;
        RECT 2.400 28.920 147.600 30.920 ;
        RECT 2.800 27.520 147.200 28.920 ;
        RECT 2.400 26.200 147.600 27.520 ;
        RECT 2.800 24.800 147.200 26.200 ;
        RECT 2.400 22.800 147.600 24.800 ;
        RECT 2.800 21.400 147.200 22.800 ;
        RECT 2.400 20.080 147.600 21.400 ;
        RECT 2.800 18.680 147.200 20.080 ;
        RECT 2.400 17.360 147.600 18.680 ;
        RECT 2.800 15.960 147.200 17.360 ;
        RECT 2.400 13.960 147.600 15.960 ;
        RECT 2.800 12.560 147.200 13.960 ;
        RECT 2.400 11.240 147.600 12.560 ;
        RECT 2.800 9.840 147.200 11.240 ;
        RECT 2.400 7.840 147.600 9.840 ;
        RECT 2.800 6.440 147.200 7.840 ;
        RECT 2.400 5.120 147.600 6.440 ;
        RECT 2.800 3.720 147.200 5.120 ;
        RECT 2.400 2.400 147.600 3.720 ;
        RECT 2.800 1.535 147.200 2.400 ;
      LAYER met4 ;
        RECT 35.750 10.640 54.320 109.040 ;
        RECT 56.720 10.640 133.530 109.040 ;
      LAYER met5 ;
        RECT 35.540 41.700 133.740 43.300 ;
  END
END cbx_1__0_
END LIBRARY

