VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__0_
  CLASS BLOCK ;
  FOREIGN sb_0__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 2.400 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 137.600 137.910 140.000 ;
    END
  END ccff_tail
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 61.240 140.000 61.840 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 89.800 140.000 90.400 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 92.520 140.000 93.120 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 95.240 140.000 95.840 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 97.960 140.000 98.560 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 104.080 140.000 104.680 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 106.800 140.000 107.400 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 109.520 140.000 110.120 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 112.240 140.000 112.840 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 115.640 140.000 116.240 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 63.960 140.000 64.560 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.680 140.000 67.280 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 69.400 140.000 70.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 72.800 140.000 73.400 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 75.520 140.000 76.120 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 78.240 140.000 78.840 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.960 140.000 81.560 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 83.680 140.000 84.280 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 4.120 140.000 4.720 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 32.680 140.000 33.280 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 35.400 140.000 36.000 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 40.840 140.000 41.440 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.240 140.000 44.840 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 46.960 140.000 47.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 49.680 140.000 50.280 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 55.120 140.000 55.720 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 58.520 140.000 59.120 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 6.840 140.000 7.440 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 9.560 140.000 10.160 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 12.280 140.000 12.880 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 15.680 140.000 16.280 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 18.400 140.000 19.000 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 21.120 140.000 21.720 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 26.560 140.000 27.160 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 29.960 140.000 30.560 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 137.600 4.970 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 137.600 38.090 140.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 137.600 41.310 140.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.710 137.600 44.990 140.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 137.600 48.210 140.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 137.600 51.430 140.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 137.600 54.650 140.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 137.600 58.330 140.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 137.600 61.550 140.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.490 137.600 64.770 140.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.710 137.600 67.990 140.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 137.600 8.190 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.130 137.600 11.410 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 137.600 14.630 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 137.600 18.310 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 137.600 21.530 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.470 137.600 24.750 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 137.600 27.970 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 137.600 31.650 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 137.600 34.870 140.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 137.600 71.670 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 104.510 137.600 104.790 140.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 137.600 108.010 140.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.950 137.600 111.230 140.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.630 137.600 114.910 140.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 137.600 118.130 140.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 137.600 121.350 140.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 137.600 124.570 140.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.970 137.600 128.250 140.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 137.600 131.470 140.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.410 137.600 134.690 140.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 137.600 74.890 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.830 137.600 78.110 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 137.600 81.330 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.270 137.600 84.550 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 137.600 88.230 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.170 137.600 91.450 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 137.600 94.670 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.610 137.600 97.890 140.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 137.600 101.570 140.000 ;
    END
  END chany_top_out[9]
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END prog_clk
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 1.400 140.000 2.000 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_top_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 118.360 140.000 118.960 ;
    END
  END right_top_grid_pin_42_
  PIN right_top_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 121.080 140.000 121.680 ;
    END
  END right_top_grid_pin_43_
  PIN right_top_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 123.800 140.000 124.400 ;
    END
  END right_top_grid_pin_44_
  PIN right_top_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 126.520 140.000 127.120 ;
    END
  END right_top_grid_pin_45_
  PIN right_top_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.920 140.000 130.520 ;
    END
  END right_top_grid_pin_46_
  PIN right_top_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 132.640 140.000 133.240 ;
    END
  END right_top_grid_pin_47_
  PIN right_top_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 135.360 140.000 135.960 ;
    END
  END right_top_grid_pin_48_
  PIN right_top_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 138.080 140.000 138.680 ;
    END
  END right_top_grid_pin_49_
  PIN top_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 137.600 1.750 140.000 ;
    END
  END top_left_grid_pin_1_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 134.320 134.940 ;
      LAYER met2 ;
        RECT 2.030 137.320 4.410 138.565 ;
        RECT 5.250 137.320 7.630 138.565 ;
        RECT 8.470 137.320 10.850 138.565 ;
        RECT 11.690 137.320 14.070 138.565 ;
        RECT 14.910 137.320 17.750 138.565 ;
        RECT 18.590 137.320 20.970 138.565 ;
        RECT 21.810 137.320 24.190 138.565 ;
        RECT 25.030 137.320 27.410 138.565 ;
        RECT 28.250 137.320 31.090 138.565 ;
        RECT 31.930 137.320 34.310 138.565 ;
        RECT 35.150 137.320 37.530 138.565 ;
        RECT 38.370 137.320 40.750 138.565 ;
        RECT 41.590 137.320 44.430 138.565 ;
        RECT 45.270 137.320 47.650 138.565 ;
        RECT 48.490 137.320 50.870 138.565 ;
        RECT 51.710 137.320 54.090 138.565 ;
        RECT 54.930 137.320 57.770 138.565 ;
        RECT 58.610 137.320 60.990 138.565 ;
        RECT 61.830 137.320 64.210 138.565 ;
        RECT 65.050 137.320 67.430 138.565 ;
        RECT 68.270 137.320 71.110 138.565 ;
        RECT 71.950 137.320 74.330 138.565 ;
        RECT 75.170 137.320 77.550 138.565 ;
        RECT 78.390 137.320 80.770 138.565 ;
        RECT 81.610 137.320 83.990 138.565 ;
        RECT 84.830 137.320 87.670 138.565 ;
        RECT 88.510 137.320 90.890 138.565 ;
        RECT 91.730 137.320 94.110 138.565 ;
        RECT 94.950 137.320 97.330 138.565 ;
        RECT 98.170 137.320 101.010 138.565 ;
        RECT 101.850 137.320 104.230 138.565 ;
        RECT 105.070 137.320 107.450 138.565 ;
        RECT 108.290 137.320 110.670 138.565 ;
        RECT 111.510 137.320 114.350 138.565 ;
        RECT 115.190 137.320 117.570 138.565 ;
        RECT 118.410 137.320 120.790 138.565 ;
        RECT 121.630 137.320 124.010 138.565 ;
        RECT 124.850 137.320 127.690 138.565 ;
        RECT 128.530 137.320 130.910 138.565 ;
        RECT 131.750 137.320 134.130 138.565 ;
        RECT 134.970 137.320 137.350 138.565 ;
        RECT 1.540 2.680 137.910 137.320 ;
        RECT 1.540 1.515 69.730 2.680 ;
        RECT 70.570 1.515 137.910 2.680 ;
      LAYER met3 ;
        RECT 1.905 137.680 137.200 138.545 ;
        RECT 1.905 136.360 137.935 137.680 ;
        RECT 1.905 134.960 137.200 136.360 ;
        RECT 1.905 133.640 137.935 134.960 ;
        RECT 1.905 132.240 137.200 133.640 ;
        RECT 1.905 130.920 137.935 132.240 ;
        RECT 1.905 129.520 137.200 130.920 ;
        RECT 1.905 127.520 137.935 129.520 ;
        RECT 1.905 126.120 137.200 127.520 ;
        RECT 1.905 124.800 137.935 126.120 ;
        RECT 1.905 123.400 137.200 124.800 ;
        RECT 1.905 122.080 137.935 123.400 ;
        RECT 1.905 120.680 137.200 122.080 ;
        RECT 1.905 119.360 137.935 120.680 ;
        RECT 1.905 117.960 137.200 119.360 ;
        RECT 1.905 116.640 137.935 117.960 ;
        RECT 1.905 115.240 137.200 116.640 ;
        RECT 1.905 113.240 137.935 115.240 ;
        RECT 1.905 111.840 137.200 113.240 ;
        RECT 1.905 110.520 137.935 111.840 ;
        RECT 1.905 109.120 137.200 110.520 ;
        RECT 1.905 107.800 137.935 109.120 ;
        RECT 1.905 106.400 137.200 107.800 ;
        RECT 1.905 105.080 137.935 106.400 ;
        RECT 1.905 103.680 137.200 105.080 ;
        RECT 1.905 102.360 137.935 103.680 ;
        RECT 1.905 100.960 137.200 102.360 ;
        RECT 1.905 98.960 137.935 100.960 ;
        RECT 1.905 97.560 137.200 98.960 ;
        RECT 1.905 96.240 137.935 97.560 ;
        RECT 1.905 94.840 137.200 96.240 ;
        RECT 1.905 93.520 137.935 94.840 ;
        RECT 1.905 92.120 137.200 93.520 ;
        RECT 1.905 90.800 137.935 92.120 ;
        RECT 1.905 89.400 137.200 90.800 ;
        RECT 1.905 88.080 137.935 89.400 ;
        RECT 1.905 86.680 137.200 88.080 ;
        RECT 1.905 84.680 137.935 86.680 ;
        RECT 1.905 83.280 137.200 84.680 ;
        RECT 1.905 81.960 137.935 83.280 ;
        RECT 1.905 80.560 137.200 81.960 ;
        RECT 1.905 79.240 137.935 80.560 ;
        RECT 1.905 77.840 137.200 79.240 ;
        RECT 1.905 76.520 137.935 77.840 ;
        RECT 1.905 75.120 137.200 76.520 ;
        RECT 1.905 73.800 137.935 75.120 ;
        RECT 1.905 72.400 137.200 73.800 ;
        RECT 1.905 71.080 137.935 72.400 ;
        RECT 2.800 70.400 137.935 71.080 ;
        RECT 2.800 69.680 137.200 70.400 ;
        RECT 1.905 69.000 137.200 69.680 ;
        RECT 1.905 67.680 137.935 69.000 ;
        RECT 1.905 66.280 137.200 67.680 ;
        RECT 1.905 64.960 137.935 66.280 ;
        RECT 1.905 63.560 137.200 64.960 ;
        RECT 1.905 62.240 137.935 63.560 ;
        RECT 1.905 60.840 137.200 62.240 ;
        RECT 1.905 59.520 137.935 60.840 ;
        RECT 1.905 58.120 137.200 59.520 ;
        RECT 1.905 56.120 137.935 58.120 ;
        RECT 1.905 54.720 137.200 56.120 ;
        RECT 1.905 53.400 137.935 54.720 ;
        RECT 1.905 52.000 137.200 53.400 ;
        RECT 1.905 50.680 137.935 52.000 ;
        RECT 1.905 49.280 137.200 50.680 ;
        RECT 1.905 47.960 137.935 49.280 ;
        RECT 1.905 46.560 137.200 47.960 ;
        RECT 1.905 45.240 137.935 46.560 ;
        RECT 1.905 43.840 137.200 45.240 ;
        RECT 1.905 41.840 137.935 43.840 ;
        RECT 1.905 40.440 137.200 41.840 ;
        RECT 1.905 39.120 137.935 40.440 ;
        RECT 1.905 37.720 137.200 39.120 ;
        RECT 1.905 36.400 137.935 37.720 ;
        RECT 1.905 35.000 137.200 36.400 ;
        RECT 1.905 33.680 137.935 35.000 ;
        RECT 1.905 32.280 137.200 33.680 ;
        RECT 1.905 30.960 137.935 32.280 ;
        RECT 1.905 29.560 137.200 30.960 ;
        RECT 1.905 27.560 137.935 29.560 ;
        RECT 1.905 26.160 137.200 27.560 ;
        RECT 1.905 24.840 137.935 26.160 ;
        RECT 1.905 23.440 137.200 24.840 ;
        RECT 1.905 22.120 137.935 23.440 ;
        RECT 1.905 20.720 137.200 22.120 ;
        RECT 1.905 19.400 137.935 20.720 ;
        RECT 1.905 18.000 137.200 19.400 ;
        RECT 1.905 16.680 137.935 18.000 ;
        RECT 1.905 15.280 137.200 16.680 ;
        RECT 1.905 13.280 137.935 15.280 ;
        RECT 1.905 11.880 137.200 13.280 ;
        RECT 1.905 10.560 137.935 11.880 ;
        RECT 1.905 9.160 137.200 10.560 ;
        RECT 1.905 7.840 137.935 9.160 ;
        RECT 1.905 6.440 137.200 7.840 ;
        RECT 1.905 5.120 137.935 6.440 ;
        RECT 1.905 3.720 137.200 5.120 ;
        RECT 1.905 2.400 137.935 3.720 ;
        RECT 1.905 1.535 137.200 2.400 ;
      LAYER met4 ;
        RECT 30.055 10.640 50.985 128.080 ;
        RECT 53.385 10.640 122.985 128.080 ;
  END
END sb_0__0_
END LIBRARY

