magic
tech sky130A
magscale 1 2
timestamp 1605107892
<< locali >>
rect 14013 24055 14047 24361
rect 22201 18615 22235 18921
rect 2881 14807 2915 15045
rect 2421 13787 2455 14025
rect 6101 13855 6135 13957
rect 6043 13821 6135 13855
<< viali >>
rect 4261 25449 4295 25483
rect 7573 25449 7607 25483
rect 11621 25449 11655 25483
rect 12909 25449 12943 25483
rect 20085 25449 20119 25483
rect 23029 25449 23063 25483
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 5181 25313 5215 25347
rect 10333 25313 10367 25347
rect 11437 25313 11471 25347
rect 12725 25313 12759 25347
rect 14197 25313 14231 25347
rect 14289 25313 14323 25347
rect 16129 25313 16163 25347
rect 18705 25313 18739 25347
rect 18797 25313 18831 25347
rect 19901 25313 19935 25347
rect 21557 25313 21591 25347
rect 24593 25313 24627 25347
rect 7665 25245 7699 25279
rect 7757 25245 7791 25279
rect 14381 25245 14415 25279
rect 16221 25245 16255 25279
rect 16313 25245 16347 25279
rect 17785 25245 17819 25279
rect 18889 25245 18923 25279
rect 21649 25245 21683 25279
rect 21833 25245 21867 25279
rect 2697 25177 2731 25211
rect 5365 25177 5399 25211
rect 10517 25177 10551 25211
rect 15301 25177 15335 25211
rect 18153 25177 18187 25211
rect 24777 25177 24811 25211
rect 1593 25109 1627 25143
rect 7205 25109 7239 25143
rect 9229 25109 9263 25143
rect 13369 25109 13403 25143
rect 13829 25109 13863 25143
rect 14841 25109 14875 25143
rect 15761 25109 15795 25143
rect 18337 25109 18371 25143
rect 19717 25109 19751 25143
rect 21005 25109 21039 25143
rect 21189 25109 21223 25143
rect 3801 24905 3835 24939
rect 4905 24905 4939 24939
rect 12265 24905 12299 24939
rect 22201 24905 22235 24939
rect 24777 24905 24811 24939
rect 4261 24769 4295 24803
rect 6285 24769 6319 24803
rect 8309 24769 8343 24803
rect 9781 24769 9815 24803
rect 13645 24769 13679 24803
rect 15209 24769 15243 24803
rect 16773 24769 16807 24803
rect 17233 24769 17267 24803
rect 18613 24769 18647 24803
rect 19533 24769 19567 24803
rect 20177 24769 20211 24803
rect 21649 24769 21683 24803
rect 21741 24769 21775 24803
rect 1409 24701 1443 24735
rect 2513 24701 2547 24735
rect 3157 24701 3191 24735
rect 3617 24701 3651 24735
rect 4721 24701 4755 24735
rect 9689 24701 9723 24735
rect 11253 24701 11287 24735
rect 13461 24701 13495 24735
rect 16681 24701 16715 24735
rect 18429 24701 18463 24735
rect 21097 24701 21131 24735
rect 24593 24701 24627 24735
rect 8033 24633 8067 24667
rect 10425 24633 10459 24667
rect 13001 24633 13035 24667
rect 15117 24633 15151 24667
rect 15761 24633 15795 24667
rect 19165 24633 19199 24667
rect 19993 24633 20027 24667
rect 22569 24633 22603 24667
rect 1593 24565 1627 24599
rect 1961 24565 1995 24599
rect 2329 24565 2363 24599
rect 2697 24565 2731 24599
rect 3525 24565 3559 24599
rect 4629 24565 4663 24599
rect 5273 24565 5307 24599
rect 6561 24565 6595 24599
rect 7297 24565 7331 24599
rect 7665 24565 7699 24599
rect 8125 24565 8159 24599
rect 8769 24565 8803 24599
rect 9045 24565 9079 24599
rect 9229 24565 9263 24599
rect 9597 24565 9631 24599
rect 10701 24565 10735 24599
rect 11161 24565 11195 24599
rect 11437 24565 11471 24599
rect 11897 24565 11931 24599
rect 13093 24565 13127 24599
rect 13553 24565 13587 24599
rect 14105 24565 14139 24599
rect 14473 24565 14507 24599
rect 14657 24565 14691 24599
rect 15025 24565 15059 24599
rect 16037 24565 16071 24599
rect 16221 24565 16255 24599
rect 16589 24565 16623 24599
rect 17785 24565 17819 24599
rect 18061 24565 18095 24599
rect 18521 24565 18555 24599
rect 19625 24565 19659 24599
rect 20085 24565 20119 24599
rect 20729 24565 20763 24599
rect 21189 24565 21223 24599
rect 21557 24565 21591 24599
rect 23029 24565 23063 24599
rect 24409 24565 24443 24599
rect 25145 24565 25179 24599
rect 4261 24361 4295 24395
rect 7665 24361 7699 24395
rect 9689 24361 9723 24395
rect 14013 24361 14047 24395
rect 18613 24361 18647 24395
rect 20177 24361 20211 24395
rect 24777 24361 24811 24395
rect 9321 24293 9355 24327
rect 1409 24225 1443 24259
rect 2513 24225 2547 24259
rect 4077 24225 4111 24259
rect 4629 24225 4663 24259
rect 6000 24225 6034 24259
rect 8493 24225 8527 24259
rect 10057 24225 10091 24259
rect 11345 24225 11379 24259
rect 13001 24225 13035 24259
rect 2053 24157 2087 24191
rect 5641 24157 5675 24191
rect 5733 24157 5767 24191
rect 10149 24157 10183 24191
rect 10241 24157 10275 24191
rect 11529 24157 11563 24191
rect 13093 24157 13127 24191
rect 13185 24157 13219 24191
rect 10701 24089 10735 24123
rect 12541 24089 12575 24123
rect 21557 24293 21591 24327
rect 23121 24293 23155 24327
rect 15301 24225 15335 24259
rect 16845 24225 16879 24259
rect 19441 24225 19475 24259
rect 21465 24225 21499 24259
rect 23029 24225 23063 24259
rect 24593 24225 24627 24259
rect 14197 24157 14231 24191
rect 15485 24157 15519 24191
rect 16589 24157 16623 24191
rect 18981 24157 19015 24191
rect 19533 24157 19567 24191
rect 19625 24157 19659 24191
rect 21649 24157 21683 24191
rect 23213 24157 23247 24191
rect 21097 24089 21131 24123
rect 22477 24089 22511 24123
rect 22661 24089 22695 24123
rect 1593 24021 1627 24055
rect 2697 24021 2731 24055
rect 3709 24021 3743 24055
rect 5273 24021 5307 24055
rect 7113 24021 7147 24055
rect 8125 24021 8159 24055
rect 8677 24021 8711 24055
rect 11069 24021 11103 24055
rect 12173 24021 12207 24055
rect 12633 24021 12667 24055
rect 13921 24021 13955 24055
rect 14013 24021 14047 24055
rect 14657 24021 14691 24055
rect 15025 24021 15059 24055
rect 16037 24021 16071 24055
rect 16405 24021 16439 24055
rect 17969 24021 18003 24055
rect 19073 24021 19107 24055
rect 20453 24021 20487 24055
rect 22109 24021 22143 24055
rect 23673 24021 23707 24055
rect 2513 23817 2547 23851
rect 2973 23817 3007 23851
rect 3525 23817 3559 23851
rect 6285 23817 6319 23851
rect 9137 23817 9171 23851
rect 14565 23817 14599 23851
rect 15025 23817 15059 23851
rect 16681 23817 16715 23851
rect 17049 23817 17083 23851
rect 17509 23817 17543 23851
rect 19533 23817 19567 23851
rect 21925 23817 21959 23851
rect 22293 23817 22327 23851
rect 22661 23817 22695 23851
rect 24593 23817 24627 23851
rect 25145 23817 25179 23851
rect 3617 23749 3651 23783
rect 9321 23749 9355 23783
rect 20729 23749 20763 23783
rect 20913 23749 20947 23783
rect 1685 23681 1719 23715
rect 4169 23681 4203 23715
rect 4721 23681 4755 23715
rect 5825 23681 5859 23715
rect 9965 23681 9999 23715
rect 10701 23681 10735 23715
rect 11253 23681 11287 23715
rect 15393 23681 15427 23715
rect 16129 23681 16163 23715
rect 20453 23681 20487 23715
rect 21465 23681 21499 23715
rect 1409 23613 1443 23647
rect 3985 23613 4019 23647
rect 6837 23613 6871 23647
rect 9781 23613 9815 23647
rect 11069 23613 11103 23647
rect 12265 23613 12299 23647
rect 12449 23613 12483 23647
rect 15945 23613 15979 23647
rect 18153 23613 18187 23647
rect 21281 23613 21315 23647
rect 22477 23613 22511 23647
rect 23029 23613 23063 23647
rect 23673 23613 23707 23647
rect 24961 23613 24995 23647
rect 25513 23613 25547 23647
rect 5089 23545 5123 23579
rect 5641 23545 5675 23579
rect 7082 23545 7116 23579
rect 8769 23545 8803 23579
rect 11897 23545 11931 23579
rect 12716 23545 12750 23579
rect 15853 23545 15887 23579
rect 17877 23545 17911 23579
rect 18420 23545 18454 23579
rect 21373 23545 21407 23579
rect 23949 23545 23983 23579
rect 2145 23477 2179 23511
rect 4077 23477 4111 23511
rect 5181 23477 5215 23511
rect 5549 23477 5583 23511
rect 6653 23477 6687 23511
rect 8217 23477 8251 23511
rect 9689 23477 9723 23511
rect 10333 23477 10367 23511
rect 13829 23477 13863 23511
rect 15485 23477 15519 23511
rect 23397 23477 23431 23511
rect 5641 23273 5675 23307
rect 6193 23273 6227 23307
rect 7757 23273 7791 23307
rect 13369 23273 13403 23307
rect 16773 23273 16807 23307
rect 19165 23273 19199 23307
rect 22569 23273 22603 23307
rect 23673 23273 23707 23307
rect 25421 23273 25455 23307
rect 3709 23205 3743 23239
rect 4506 23205 4540 23239
rect 8585 23205 8619 23239
rect 10241 23205 10275 23239
rect 11704 23205 11738 23239
rect 14197 23205 14231 23239
rect 17325 23205 17359 23239
rect 20729 23205 20763 23239
rect 21456 23205 21490 23239
rect 1501 23137 1535 23171
rect 2605 23137 2639 23171
rect 2789 23137 2823 23171
rect 7113 23137 7147 23171
rect 8309 23137 8343 23171
rect 13921 23137 13955 23171
rect 14749 23137 14783 23171
rect 15117 23137 15151 23171
rect 15393 23137 15427 23171
rect 15660 23137 15694 23171
rect 17969 23137 18003 23171
rect 19625 23137 19659 23171
rect 24041 23137 24075 23171
rect 25237 23137 25271 23171
rect 1777 23069 1811 23103
rect 4261 23069 4295 23103
rect 7205 23069 7239 23103
rect 7389 23069 7423 23103
rect 8217 23069 8251 23103
rect 10333 23069 10367 23103
rect 10517 23069 10551 23103
rect 11437 23069 11471 23103
rect 18153 23069 18187 23103
rect 19717 23069 19751 23103
rect 19809 23069 19843 23103
rect 21189 23069 21223 23103
rect 23581 23069 23615 23103
rect 24133 23069 24167 23103
rect 24225 23069 24259 23103
rect 6745 23001 6779 23035
rect 13737 23001 13771 23035
rect 20269 23001 20303 23035
rect 2329 22933 2363 22967
rect 2973 22933 3007 22967
rect 6561 22933 6595 22967
rect 9413 22933 9447 22967
rect 9873 22933 9907 22967
rect 10977 22933 11011 22967
rect 11253 22933 11287 22967
rect 12817 22933 12851 22967
rect 17877 22933 17911 22967
rect 18797 22933 18831 22967
rect 19257 22933 19291 22967
rect 23121 22933 23155 22967
rect 5641 22729 5675 22763
rect 7113 22729 7147 22763
rect 10333 22729 10367 22763
rect 11897 22729 11931 22763
rect 15025 22729 15059 22763
rect 18245 22729 18279 22763
rect 19349 22729 19383 22763
rect 21189 22729 21223 22763
rect 21741 22729 21775 22763
rect 23121 22729 23155 22763
rect 25421 22729 25455 22763
rect 9965 22661 9999 22695
rect 16865 22661 16899 22695
rect 2973 22593 3007 22627
rect 9597 22593 9631 22627
rect 11437 22593 11471 22627
rect 12449 22593 12483 22627
rect 17877 22593 17911 22627
rect 18705 22593 18739 22627
rect 18889 22593 18923 22627
rect 24317 22593 24351 22627
rect 1501 22525 1535 22559
rect 5457 22525 5491 22559
rect 6009 22525 6043 22559
rect 7389 22525 7423 22559
rect 7645 22525 7679 22559
rect 10609 22525 10643 22559
rect 11161 22525 11195 22559
rect 12716 22525 12750 22559
rect 15485 22525 15519 22559
rect 19625 22525 19659 22559
rect 19809 22525 19843 22559
rect 20065 22525 20099 22559
rect 22293 22525 22327 22559
rect 23489 22525 23523 22559
rect 24133 22525 24167 22559
rect 25237 22525 25271 22559
rect 1777 22457 1811 22491
rect 2513 22457 2547 22491
rect 3218 22457 3252 22491
rect 11253 22457 11287 22491
rect 12265 22457 12299 22491
rect 15393 22457 15427 22491
rect 15752 22457 15786 22491
rect 17509 22457 17543 22491
rect 18613 22457 18647 22491
rect 22569 22457 22603 22491
rect 24041 22457 24075 22491
rect 24685 22457 24719 22491
rect 2881 22389 2915 22423
rect 4353 22389 4387 22423
rect 4905 22389 4939 22423
rect 5365 22389 5399 22423
rect 6653 22389 6687 22423
rect 8769 22389 8803 22423
rect 10793 22389 10827 22423
rect 13829 22389 13863 22423
rect 14381 22389 14415 22423
rect 22109 22389 22143 22423
rect 23673 22389 23707 22423
rect 25145 22389 25179 22423
rect 25789 22389 25823 22423
rect 2421 22185 2455 22219
rect 2789 22185 2823 22219
rect 3433 22185 3467 22219
rect 4537 22185 4571 22219
rect 6009 22185 6043 22219
rect 7573 22185 7607 22219
rect 7941 22185 7975 22219
rect 10425 22185 10459 22219
rect 11161 22185 11195 22219
rect 12357 22185 12391 22219
rect 12725 22185 12759 22219
rect 13829 22185 13863 22219
rect 15117 22185 15151 22219
rect 16681 22185 16715 22219
rect 17969 22185 18003 22219
rect 19901 22185 19935 22219
rect 20269 22185 20303 22219
rect 24133 22185 24167 22219
rect 1409 22117 1443 22151
rect 2881 22117 2915 22151
rect 4445 22117 4479 22151
rect 7389 22117 7423 22151
rect 13369 22117 13403 22151
rect 22376 22117 22410 22151
rect 24409 22117 24443 22151
rect 1961 22049 1995 22083
rect 6377 22049 6411 22083
rect 7113 22049 7147 22083
rect 8033 22049 8067 22083
rect 11897 22049 11931 22083
rect 13921 22049 13955 22083
rect 14657 22049 14691 22083
rect 15669 22049 15703 22083
rect 17049 22049 17083 22083
rect 18705 22049 18739 22083
rect 21005 22049 21039 22083
rect 24961 22049 24995 22083
rect 3065 21981 3099 22015
rect 4629 21981 4663 22015
rect 6469 21981 6503 22015
rect 6653 21981 6687 22015
rect 8125 21981 8159 22015
rect 9505 21981 9539 22015
rect 9965 21981 9999 22015
rect 10517 21981 10551 22015
rect 10701 21981 10735 22015
rect 12265 21981 12299 22015
rect 12817 21981 12851 22015
rect 13001 21981 13035 22015
rect 14197 21981 14231 22015
rect 15761 21981 15795 22015
rect 15945 21981 15979 22015
rect 17325 21981 17359 22015
rect 18797 21981 18831 22015
rect 18981 21981 19015 22015
rect 22109 21981 22143 22015
rect 25053 21981 25087 22015
rect 25237 21981 25271 22015
rect 25605 21981 25639 22015
rect 2329 21913 2363 21947
rect 4077 21913 4111 21947
rect 8953 21913 8987 21947
rect 15301 21913 15335 21947
rect 18337 21913 18371 21947
rect 21189 21913 21223 21947
rect 3801 21845 3835 21879
rect 5089 21845 5123 21879
rect 5457 21845 5491 21879
rect 5825 21845 5859 21879
rect 8677 21845 8711 21879
rect 10057 21845 10091 21879
rect 11437 21845 11471 21879
rect 16313 21845 16347 21879
rect 19441 21845 19475 21879
rect 20545 21845 20579 21879
rect 21557 21845 21591 21879
rect 22017 21845 22051 21879
rect 23489 21845 23523 21879
rect 24593 21845 24627 21879
rect 2605 21641 2639 21675
rect 4997 21641 5031 21675
rect 5365 21641 5399 21675
rect 6561 21641 6595 21675
rect 7665 21641 7699 21675
rect 9137 21641 9171 21675
rect 10149 21641 10183 21675
rect 10517 21641 10551 21675
rect 12265 21641 12299 21675
rect 12449 21641 12483 21675
rect 14013 21641 14047 21675
rect 15025 21641 15059 21675
rect 16957 21641 16991 21675
rect 17509 21641 17543 21675
rect 20177 21641 20211 21675
rect 22017 21641 22051 21675
rect 25973 21641 26007 21675
rect 17785 21573 17819 21607
rect 21925 21573 21959 21607
rect 23121 21573 23155 21607
rect 2053 21505 2087 21539
rect 2973 21505 3007 21539
rect 7757 21505 7791 21539
rect 11253 21505 11287 21539
rect 11437 21505 11471 21539
rect 12909 21505 12943 21539
rect 13001 21505 13035 21539
rect 14565 21505 14599 21539
rect 16129 21505 16163 21539
rect 22477 21505 22511 21539
rect 22661 21505 22695 21539
rect 23673 21505 23707 21539
rect 3065 21437 3099 21471
rect 3332 21437 3366 21471
rect 5549 21437 5583 21471
rect 12817 21437 12851 21471
rect 13461 21437 13495 21471
rect 16037 21437 16071 21471
rect 18797 21437 18831 21471
rect 19064 21437 19098 21471
rect 22385 21437 22419 21471
rect 23940 21437 23974 21471
rect 1961 21369 1995 21403
rect 7297 21369 7331 21403
rect 8024 21369 8058 21403
rect 9781 21369 9815 21403
rect 11161 21369 11195 21403
rect 14473 21369 14507 21403
rect 15945 21369 15979 21403
rect 16589 21369 16623 21403
rect 21557 21369 21591 21403
rect 23489 21369 23523 21403
rect 1501 21301 1535 21335
rect 1869 21301 1903 21335
rect 4445 21301 4479 21335
rect 5733 21301 5767 21335
rect 6101 21301 6135 21335
rect 10793 21301 10827 21335
rect 11897 21301 11931 21335
rect 13921 21301 13955 21335
rect 14381 21301 14415 21335
rect 15393 21301 15427 21335
rect 15577 21301 15611 21335
rect 18429 21301 18463 21335
rect 21097 21301 21131 21335
rect 25053 21301 25087 21335
rect 25697 21301 25731 21335
rect 1409 21097 1443 21131
rect 2329 21097 2363 21131
rect 2421 21097 2455 21131
rect 4629 21097 4663 21131
rect 6285 21097 6319 21131
rect 6837 21097 6871 21131
rect 7757 21097 7791 21131
rect 7849 21097 7883 21131
rect 8401 21097 8435 21131
rect 10517 21097 10551 21131
rect 11989 21097 12023 21131
rect 12909 21097 12943 21131
rect 13093 21097 13127 21131
rect 14105 21097 14139 21131
rect 15117 21097 15151 21131
rect 15577 21097 15611 21131
rect 17049 21097 17083 21131
rect 17601 21097 17635 21131
rect 19165 21097 19199 21131
rect 19901 21097 19935 21131
rect 20729 21097 20763 21131
rect 20913 21097 20947 21131
rect 22477 21097 22511 21131
rect 25421 21097 25455 21131
rect 12633 21029 12667 21063
rect 18061 21029 18095 21063
rect 18521 21029 18555 21063
rect 23029 21029 23063 21063
rect 23305 21029 23339 21063
rect 23756 21029 23790 21063
rect 2789 20961 2823 20995
rect 3433 20961 3467 20995
rect 5172 20961 5206 20995
rect 10876 20961 10910 20995
rect 13461 20961 13495 20995
rect 13553 20961 13587 20995
rect 15669 20961 15703 20995
rect 15936 20961 15970 20995
rect 18613 20961 18647 20995
rect 19717 20961 19751 20995
rect 21281 20961 21315 20995
rect 23489 20961 23523 20995
rect 2881 20893 2915 20927
rect 2973 20893 3007 20927
rect 4261 20893 4295 20927
rect 4905 20893 4939 20927
rect 7297 20893 7331 20927
rect 7941 20893 7975 20927
rect 10609 20893 10643 20927
rect 13645 20893 13679 20927
rect 18705 20893 18739 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 8861 20825 8895 20859
rect 19533 20825 19567 20859
rect 20269 20825 20303 20859
rect 1961 20757 1995 20791
rect 3893 20757 3927 20791
rect 7389 20757 7423 20791
rect 9137 20757 9171 20791
rect 9873 20757 9907 20791
rect 14473 20757 14507 20791
rect 18153 20757 18187 20791
rect 22109 20757 22143 20791
rect 24869 20757 24903 20791
rect 2605 20553 2639 20587
rect 7665 20553 7699 20587
rect 7941 20553 7975 20587
rect 10793 20553 10827 20587
rect 11897 20553 11931 20587
rect 14289 20553 14323 20587
rect 16037 20553 16071 20587
rect 16681 20553 16715 20587
rect 18337 20553 18371 20587
rect 20085 20553 20119 20587
rect 23489 20553 23523 20587
rect 6469 20485 6503 20519
rect 10333 20485 10367 20519
rect 12449 20485 12483 20519
rect 13461 20485 13495 20519
rect 17509 20485 17543 20519
rect 23673 20485 23707 20519
rect 3249 20417 3283 20451
rect 4353 20417 4387 20451
rect 5089 20417 5123 20451
rect 7113 20417 7147 20451
rect 8125 20417 8159 20451
rect 11437 20417 11471 20451
rect 13093 20417 13127 20451
rect 21557 20417 21591 20451
rect 22569 20417 22603 20451
rect 24225 20417 24259 20451
rect 1409 20349 1443 20383
rect 3065 20349 3099 20383
rect 4813 20349 4847 20383
rect 6193 20349 6227 20383
rect 6653 20349 6687 20383
rect 8392 20349 8426 20383
rect 14657 20349 14691 20383
rect 17877 20349 17911 20383
rect 18705 20349 18739 20383
rect 18972 20349 19006 20383
rect 21833 20349 21867 20383
rect 25237 20349 25271 20383
rect 25973 20349 26007 20383
rect 2421 20281 2455 20315
rect 4905 20281 4939 20315
rect 11161 20281 11195 20315
rect 12817 20281 12851 20315
rect 14924 20281 14958 20315
rect 22477 20281 22511 20315
rect 24041 20281 24075 20315
rect 25053 20281 25087 20315
rect 25513 20281 25547 20315
rect 1593 20213 1627 20247
rect 2053 20213 2087 20247
rect 2973 20213 3007 20247
rect 3617 20213 3651 20247
rect 4445 20213 4479 20247
rect 5549 20213 5583 20247
rect 5917 20213 5951 20247
rect 9505 20213 9539 20247
rect 10609 20213 10643 20247
rect 11253 20213 11287 20247
rect 12173 20213 12207 20247
rect 12909 20213 12943 20247
rect 13921 20213 13955 20247
rect 17233 20213 17267 20247
rect 17693 20213 17727 20247
rect 20913 20213 20947 20247
rect 22017 20213 22051 20247
rect 22385 20213 22419 20247
rect 23029 20213 23063 20247
rect 24133 20213 24167 20247
rect 24685 20213 24719 20247
rect 1409 20009 1443 20043
rect 3525 20009 3559 20043
rect 8401 20009 8435 20043
rect 10149 20009 10183 20043
rect 11989 20009 12023 20043
rect 12633 20009 12667 20043
rect 13553 20009 13587 20043
rect 14749 20009 14783 20043
rect 16681 20009 16715 20043
rect 19625 20009 19659 20043
rect 20729 20009 20763 20043
rect 22385 20009 22419 20043
rect 23121 20009 23155 20043
rect 23489 20009 23523 20043
rect 25145 20009 25179 20043
rect 2329 19941 2363 19975
rect 9045 19941 9079 19975
rect 10517 19941 10551 19975
rect 10876 19941 10910 19975
rect 15568 19941 15602 19975
rect 18512 19941 18546 19975
rect 24032 19941 24066 19975
rect 2789 19873 2823 19907
rect 5080 19873 5114 19907
rect 7665 19873 7699 19907
rect 9505 19873 9539 19907
rect 13461 19873 13495 19907
rect 15301 19873 15335 19907
rect 17969 19873 18003 19907
rect 18245 19873 18279 19907
rect 21005 19873 21039 19907
rect 21272 19873 21306 19907
rect 23765 19873 23799 19907
rect 2881 19805 2915 19839
rect 3065 19805 3099 19839
rect 4813 19805 4847 19839
rect 7757 19805 7791 19839
rect 7941 19805 7975 19839
rect 8769 19805 8803 19839
rect 10609 19805 10643 19839
rect 13645 19805 13679 19839
rect 1961 19737 1995 19771
rect 2421 19737 2455 19771
rect 13001 19737 13035 19771
rect 15025 19737 15059 19771
rect 17325 19737 17359 19771
rect 17785 19737 17819 19771
rect 3801 19669 3835 19703
rect 4353 19669 4387 19703
rect 4721 19669 4755 19703
rect 6193 19669 6227 19703
rect 6837 19669 6871 19703
rect 7297 19669 7331 19703
rect 9321 19669 9355 19703
rect 13093 19669 13127 19703
rect 14197 19669 14231 19703
rect 17601 19669 17635 19703
rect 20177 19669 20211 19703
rect 3709 19465 3743 19499
rect 5641 19465 5675 19499
rect 6837 19465 6871 19499
rect 11345 19465 11379 19499
rect 12449 19465 12483 19499
rect 13553 19465 13587 19499
rect 16957 19465 16991 19499
rect 19165 19465 19199 19499
rect 23765 19465 23799 19499
rect 2513 19397 2547 19431
rect 6653 19397 6687 19431
rect 10241 19397 10275 19431
rect 3341 19329 3375 19363
rect 7389 19329 7423 19363
rect 9229 19329 9263 19363
rect 9781 19329 9815 19363
rect 10885 19329 10919 19363
rect 11897 19329 11931 19363
rect 13001 19329 13035 19363
rect 14565 19329 14599 19363
rect 16221 19329 16255 19363
rect 16589 19329 16623 19363
rect 18613 19329 18647 19363
rect 20821 19329 20855 19363
rect 24317 19329 24351 19363
rect 24777 19329 24811 19363
rect 1409 19261 1443 19295
rect 4261 19261 4295 19295
rect 6285 19261 6319 19295
rect 7297 19261 7331 19295
rect 10609 19261 10643 19295
rect 12909 19261 12943 19295
rect 15025 19261 15059 19295
rect 15485 19261 15519 19295
rect 16037 19261 16071 19295
rect 18429 19261 18463 19295
rect 19625 19261 19659 19295
rect 25145 19261 25179 19295
rect 25329 19261 25363 19295
rect 26065 19261 26099 19295
rect 1685 19193 1719 19227
rect 3157 19193 3191 19227
rect 4169 19193 4203 19227
rect 4528 19193 4562 19227
rect 8585 19193 8619 19227
rect 9137 19193 9171 19227
rect 10057 19193 10091 19227
rect 14381 19193 14415 19227
rect 15945 19193 15979 19227
rect 18521 19193 18555 19227
rect 20361 19193 20395 19227
rect 21066 19193 21100 19227
rect 23121 19193 23155 19227
rect 24133 19193 24167 19227
rect 25605 19193 25639 19227
rect 2697 19125 2731 19159
rect 3065 19125 3099 19159
rect 7205 19125 7239 19159
rect 7849 19125 7883 19159
rect 8677 19125 8711 19159
rect 9045 19125 9079 19159
rect 10701 19125 10735 19159
rect 12173 19125 12207 19159
rect 12817 19125 12851 19159
rect 13829 19125 13863 19159
rect 14013 19125 14047 19159
rect 14473 19125 14507 19159
rect 15577 19125 15611 19159
rect 17417 19125 17451 19159
rect 17785 19125 17819 19159
rect 18061 19125 18095 19159
rect 19533 19125 19567 19159
rect 19809 19125 19843 19159
rect 20729 19125 20763 19159
rect 22201 19125 22235 19159
rect 23489 19125 23523 19159
rect 24225 19125 24259 19159
rect 2513 18921 2547 18955
rect 3065 18921 3099 18955
rect 5273 18921 5307 18955
rect 6469 18921 6503 18955
rect 6837 18921 6871 18955
rect 7573 18921 7607 18955
rect 9137 18921 9171 18955
rect 10241 18921 10275 18955
rect 14381 18921 14415 18955
rect 15025 18921 15059 18955
rect 15761 18921 15795 18955
rect 18245 18921 18279 18955
rect 21925 18921 21959 18955
rect 22201 18921 22235 18955
rect 22477 18921 22511 18955
rect 23489 18921 23523 18955
rect 25237 18921 25271 18955
rect 5181 18853 5215 18887
rect 6009 18853 6043 18887
rect 8493 18853 8527 18887
rect 10692 18853 10726 18887
rect 15669 18853 15703 18887
rect 16313 18853 16347 18887
rect 2421 18785 2455 18819
rect 6377 18785 6411 18819
rect 8401 18785 8435 18819
rect 13277 18785 13311 18819
rect 18153 18785 18187 18819
rect 19349 18785 19383 18819
rect 20085 18785 20119 18819
rect 20729 18785 20763 18819
rect 21281 18785 21315 18819
rect 21373 18785 21407 18819
rect 2697 18717 2731 18751
rect 4353 18717 4387 18751
rect 4721 18717 4755 18751
rect 5457 18717 5491 18751
rect 6929 18717 6963 18751
rect 7113 18717 7147 18751
rect 8585 18717 8619 18751
rect 10425 18717 10459 18751
rect 13369 18717 13403 18751
rect 13461 18717 13495 18751
rect 15853 18717 15887 18751
rect 18429 18717 18463 18751
rect 19533 18717 19567 18751
rect 21465 18717 21499 18751
rect 1961 18649 1995 18683
rect 4813 18649 4847 18683
rect 7941 18649 7975 18683
rect 16773 18649 16807 18683
rect 17141 18649 17175 18683
rect 24501 18853 24535 18887
rect 23857 18785 23891 18819
rect 25053 18785 25087 18819
rect 23949 18717 23983 18751
rect 24041 18717 24075 18751
rect 2053 18581 2087 18615
rect 3525 18581 3559 18615
rect 3893 18581 3927 18615
rect 8033 18581 8067 18615
rect 9505 18581 9539 18615
rect 9873 18581 9907 18615
rect 11805 18581 11839 18615
rect 12449 18581 12483 18615
rect 12909 18581 12943 18615
rect 14013 18581 14047 18615
rect 15301 18581 15335 18615
rect 17693 18581 17727 18615
rect 17785 18581 17819 18615
rect 18889 18581 18923 18615
rect 19257 18581 19291 18615
rect 20913 18581 20947 18615
rect 22201 18581 22235 18615
rect 22385 18581 22419 18615
rect 23305 18581 23339 18615
rect 1777 18377 1811 18411
rect 2145 18377 2179 18411
rect 4261 18377 4295 18411
rect 5181 18377 5215 18411
rect 6561 18377 6595 18411
rect 8125 18377 8159 18411
rect 9873 18377 9907 18411
rect 10517 18377 10551 18411
rect 16865 18377 16899 18411
rect 17509 18377 17543 18411
rect 17877 18377 17911 18411
rect 19809 18377 19843 18411
rect 19993 18377 20027 18411
rect 21005 18377 21039 18411
rect 22569 18377 22603 18411
rect 23121 18377 23155 18411
rect 25053 18377 25087 18411
rect 25605 18377 25639 18411
rect 5733 18241 5767 18275
rect 7389 18241 7423 18275
rect 11897 18241 11931 18275
rect 18521 18241 18555 18275
rect 18705 18241 18739 18275
rect 20545 18241 20579 18275
rect 22109 18241 22143 18275
rect 2329 18173 2363 18207
rect 8493 18173 8527 18207
rect 11253 18173 11287 18207
rect 12265 18173 12299 18207
rect 13001 18173 13035 18207
rect 15485 18173 15519 18207
rect 18429 18173 18463 18207
rect 20453 18173 20487 18207
rect 21925 18173 21959 18207
rect 23673 18173 23707 18207
rect 23929 18173 23963 18207
rect 2574 18105 2608 18139
rect 4721 18105 4755 18139
rect 5549 18105 5583 18139
rect 7205 18105 7239 18139
rect 8738 18105 8772 18139
rect 13268 18105 13302 18139
rect 14933 18105 14967 18139
rect 15752 18105 15786 18139
rect 21465 18105 21499 18139
rect 22017 18105 22051 18139
rect 3709 18037 3743 18071
rect 4997 18037 5031 18071
rect 5641 18037 5675 18071
rect 6837 18037 6871 18071
rect 7297 18037 7331 18071
rect 10793 18037 10827 18071
rect 11437 18037 11471 18071
rect 12817 18037 12851 18071
rect 14381 18037 14415 18071
rect 15393 18037 15427 18071
rect 18061 18037 18095 18071
rect 19073 18037 19107 18071
rect 19533 18037 19567 18071
rect 20361 18037 20395 18071
rect 21557 18037 21591 18071
rect 23489 18037 23523 18071
rect 1593 17833 1627 17867
rect 1869 17833 1903 17867
rect 3249 17833 3283 17867
rect 5457 17833 5491 17867
rect 6745 17833 6779 17867
rect 8033 17833 8067 17867
rect 8493 17833 8527 17867
rect 10149 17833 10183 17867
rect 12633 17833 12667 17867
rect 13553 17833 13587 17867
rect 16681 17833 16715 17867
rect 17325 17833 17359 17867
rect 18245 17833 18279 17867
rect 18797 17833 18831 17867
rect 20729 17833 20763 17867
rect 22661 17833 22695 17867
rect 23581 17833 23615 17867
rect 25053 17833 25087 17867
rect 9137 17765 9171 17799
rect 9413 17765 9447 17799
rect 11520 17765 11554 17799
rect 13185 17765 13219 17799
rect 14197 17765 14231 17799
rect 15546 17765 15580 17799
rect 17693 17765 17727 17799
rect 19165 17765 19199 17799
rect 19625 17765 19659 17799
rect 21373 17765 21407 17799
rect 23918 17765 23952 17799
rect 2237 17697 2271 17731
rect 2329 17697 2363 17731
rect 3617 17697 3651 17731
rect 4333 17697 4367 17731
rect 6561 17697 6595 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 11253 17697 11287 17731
rect 13921 17697 13955 17731
rect 15301 17697 15335 17731
rect 18153 17697 18187 17731
rect 19349 17697 19383 17731
rect 21281 17697 21315 17731
rect 22477 17697 22511 17731
rect 2421 17629 2455 17663
rect 4077 17629 4111 17663
rect 6469 17629 6503 17663
rect 8677 17629 8711 17663
rect 10333 17629 10367 17663
rect 18337 17629 18371 17663
rect 21465 17629 21499 17663
rect 23673 17629 23707 17663
rect 6101 17561 6135 17595
rect 9689 17561 9723 17595
rect 14933 17561 14967 17595
rect 17785 17561 17819 17595
rect 20913 17561 20947 17595
rect 2973 17493 3007 17527
rect 7113 17493 7147 17527
rect 7573 17493 7607 17527
rect 7941 17493 7975 17527
rect 10885 17493 10919 17527
rect 20177 17493 20211 17527
rect 21925 17493 21959 17527
rect 1961 17289 1995 17323
rect 4169 17289 4203 17323
rect 4629 17289 4663 17323
rect 4905 17289 4939 17323
rect 5089 17289 5123 17323
rect 6101 17289 6135 17323
rect 6561 17289 6595 17323
rect 9689 17289 9723 17323
rect 10241 17289 10275 17323
rect 14933 17289 14967 17323
rect 15945 17289 15979 17323
rect 17877 17289 17911 17323
rect 19993 17289 20027 17323
rect 22385 17289 22419 17323
rect 23121 17289 23155 17323
rect 23489 17289 23523 17323
rect 7021 17221 7055 17255
rect 14749 17221 14783 17255
rect 21833 17221 21867 17255
rect 23673 17221 23707 17255
rect 5641 17153 5675 17187
rect 7757 17153 7791 17187
rect 8125 17153 8159 17187
rect 11345 17153 11379 17187
rect 12449 17153 12483 17187
rect 15485 17153 15519 17187
rect 17509 17153 17543 17187
rect 18705 17153 18739 17187
rect 24317 17153 24351 17187
rect 2145 17085 2179 17119
rect 5549 17085 5583 17119
rect 6837 17085 6871 17119
rect 8309 17085 8343 17119
rect 8576 17085 8610 17119
rect 11253 17085 11287 17119
rect 15301 17085 15335 17119
rect 16497 17085 16531 17119
rect 20453 17085 20487 17119
rect 25237 17085 25271 17119
rect 25973 17085 26007 17119
rect 2412 17017 2446 17051
rect 12265 17017 12299 17051
rect 12694 17017 12728 17051
rect 15393 17017 15427 17051
rect 16773 17017 16807 17051
rect 18429 17017 18463 17051
rect 19441 17017 19475 17051
rect 20698 17017 20732 17051
rect 24041 17017 24075 17051
rect 25053 17017 25087 17051
rect 25513 17017 25547 17051
rect 3525 16949 3559 16983
rect 5457 16949 5491 16983
rect 10609 16949 10643 16983
rect 10793 16949 10827 16983
rect 11161 16949 11195 16983
rect 11897 16949 11931 16983
rect 13829 16949 13863 16983
rect 14381 16949 14415 16983
rect 16313 16949 16347 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19073 16949 19107 16983
rect 20361 16949 20395 16983
rect 24133 16949 24167 16983
rect 24685 16949 24719 16983
rect 1869 16745 1903 16779
rect 3341 16745 3375 16779
rect 5181 16745 5215 16779
rect 6745 16745 6779 16779
rect 8033 16745 8067 16779
rect 9045 16745 9079 16779
rect 9689 16745 9723 16779
rect 10149 16745 10183 16779
rect 10885 16745 10919 16779
rect 12633 16745 12667 16779
rect 14933 16745 14967 16779
rect 15301 16745 15335 16779
rect 18981 16745 19015 16779
rect 19441 16745 19475 16779
rect 19717 16745 19751 16779
rect 22293 16745 22327 16779
rect 22937 16745 22971 16779
rect 23305 16745 23339 16779
rect 25145 16745 25179 16779
rect 2329 16677 2363 16711
rect 3617 16677 3651 16711
rect 4353 16677 4387 16711
rect 7297 16677 7331 16711
rect 8493 16677 8527 16711
rect 9505 16677 9539 16711
rect 14197 16677 14231 16711
rect 15761 16677 15795 16711
rect 16773 16677 16807 16711
rect 17316 16677 17350 16711
rect 21180 16677 21214 16711
rect 1777 16609 1811 16643
rect 2237 16609 2271 16643
rect 2973 16609 3007 16643
rect 4077 16609 4111 16643
rect 5632 16609 5666 16643
rect 8401 16609 8435 16643
rect 10057 16609 10091 16643
rect 11253 16609 11287 16643
rect 11520 16609 11554 16643
rect 13461 16609 13495 16643
rect 13921 16609 13955 16643
rect 15669 16609 15703 16643
rect 17049 16609 17083 16643
rect 19533 16609 19567 16643
rect 20545 16609 20579 16643
rect 23581 16609 23615 16643
rect 23765 16609 23799 16643
rect 24032 16609 24066 16643
rect 2421 16541 2455 16575
rect 5365 16541 5399 16575
rect 8677 16541 8711 16575
rect 10241 16541 10275 16575
rect 15853 16541 15887 16575
rect 20177 16541 20211 16575
rect 20913 16541 20947 16575
rect 7941 16473 7975 16507
rect 18429 16473 18463 16507
rect 13829 16405 13863 16439
rect 16497 16405 16531 16439
rect 2513 16201 2547 16235
rect 2789 16201 2823 16235
rect 6285 16201 6319 16235
rect 6653 16201 6687 16235
rect 7113 16201 7147 16235
rect 9597 16201 9631 16235
rect 10149 16201 10183 16235
rect 10517 16201 10551 16235
rect 10793 16201 10827 16235
rect 11805 16201 11839 16235
rect 12173 16201 12207 16235
rect 14013 16201 14047 16235
rect 15393 16201 15427 16235
rect 16405 16201 16439 16235
rect 19441 16201 19475 16235
rect 20637 16201 20671 16235
rect 20913 16201 20947 16235
rect 23765 16201 23799 16235
rect 25513 16201 25547 16235
rect 7757 16133 7791 16167
rect 8033 16133 8067 16167
rect 19993 16133 20027 16167
rect 3249 16065 3283 16099
rect 3433 16065 3467 16099
rect 5733 16065 5767 16099
rect 7205 16065 7239 16099
rect 8217 16065 8251 16099
rect 11437 16065 11471 16099
rect 12909 16065 12943 16099
rect 13093 16065 13127 16099
rect 14565 16065 14599 16099
rect 15945 16065 15979 16099
rect 17049 16065 17083 16099
rect 17877 16065 17911 16099
rect 24317 16065 24351 16099
rect 24777 16065 24811 16099
rect 25145 16065 25179 16099
rect 1409 15997 1443 16031
rect 3157 15997 3191 16031
rect 5641 15997 5675 16031
rect 8484 15997 8518 16031
rect 16773 15997 16807 16031
rect 18061 15997 18095 16031
rect 18328 15997 18362 16031
rect 21097 15997 21131 16031
rect 21353 15997 21387 16031
rect 25329 15997 25363 16031
rect 25881 15997 25915 16031
rect 1685 15929 1719 15963
rect 2237 15929 2271 15963
rect 3801 15929 3835 15963
rect 4721 15929 4755 15963
rect 5549 15929 5583 15963
rect 11253 15929 11287 15963
rect 16313 15929 16347 15963
rect 16865 15929 16899 15963
rect 23029 15929 23063 15963
rect 24133 15929 24167 15963
rect 4261 15861 4295 15895
rect 4997 15861 5031 15895
rect 5181 15861 5215 15895
rect 11161 15861 11195 15895
rect 12449 15861 12483 15895
rect 12817 15861 12851 15895
rect 13461 15861 13495 15895
rect 13829 15861 13863 15895
rect 14381 15861 14415 15895
rect 14473 15861 14507 15895
rect 17509 15861 17543 15895
rect 22477 15861 22511 15895
rect 23489 15861 23523 15895
rect 24225 15861 24259 15895
rect 1961 15657 1995 15691
rect 3525 15657 3559 15691
rect 4261 15657 4295 15691
rect 4997 15657 5031 15691
rect 6009 15657 6043 15691
rect 9137 15657 9171 15691
rect 9873 15657 9907 15691
rect 10333 15657 10367 15691
rect 10793 15657 10827 15691
rect 12909 15657 12943 15691
rect 14749 15657 14783 15691
rect 18245 15657 18279 15691
rect 20913 15657 20947 15691
rect 22293 15657 22327 15691
rect 24777 15657 24811 15691
rect 7380 15589 7414 15623
rect 11130 15589 11164 15623
rect 18153 15589 18187 15623
rect 23642 15589 23676 15623
rect 2329 15521 2363 15555
rect 4077 15521 4111 15555
rect 5365 15521 5399 15555
rect 5917 15521 5951 15555
rect 7113 15521 7147 15555
rect 9505 15521 9539 15555
rect 13737 15521 13771 15555
rect 15669 15521 15703 15555
rect 16028 15521 16062 15555
rect 18613 15521 18647 15555
rect 20729 15521 20763 15555
rect 21281 15521 21315 15555
rect 22661 15521 22695 15555
rect 2421 15453 2455 15487
rect 2513 15453 2547 15487
rect 6101 15453 6135 15487
rect 10885 15453 10919 15487
rect 13829 15453 13863 15487
rect 13921 15453 13955 15487
rect 14381 15453 14415 15487
rect 15761 15453 15795 15487
rect 18705 15453 18739 15487
rect 18889 15453 18923 15487
rect 19809 15453 19843 15487
rect 21373 15453 21407 15487
rect 21557 15453 21591 15487
rect 23397 15453 23431 15487
rect 4629 15385 4663 15419
rect 5549 15385 5583 15419
rect 12265 15385 12299 15419
rect 17141 15385 17175 15419
rect 1685 15317 1719 15351
rect 3249 15317 3283 15351
rect 5181 15317 5215 15351
rect 6929 15317 6963 15351
rect 8493 15317 8527 15351
rect 13185 15317 13219 15351
rect 13369 15317 13403 15351
rect 17693 15317 17727 15351
rect 19349 15317 19383 15351
rect 19625 15317 19659 15351
rect 20361 15317 20395 15351
rect 21925 15317 21959 15351
rect 22477 15317 22511 15351
rect 23305 15317 23339 15351
rect 3065 15113 3099 15147
rect 5181 15113 5215 15147
rect 5549 15113 5583 15147
rect 7941 15113 7975 15147
rect 8861 15113 8895 15147
rect 10977 15113 11011 15147
rect 11805 15113 11839 15147
rect 12449 15113 12483 15147
rect 13553 15113 13587 15147
rect 15945 15113 15979 15147
rect 17877 15113 17911 15147
rect 20361 15113 20395 15147
rect 20913 15113 20947 15147
rect 21925 15113 21959 15147
rect 22661 15113 22695 15147
rect 23029 15113 23063 15147
rect 23765 15113 23799 15147
rect 24777 15113 24811 15147
rect 25513 15113 25547 15147
rect 2605 15045 2639 15079
rect 2881 15045 2915 15079
rect 4537 15045 4571 15079
rect 14013 15045 14047 15079
rect 22385 15045 22419 15079
rect 2237 14977 2271 15011
rect 1961 14841 1995 14875
rect 7389 14977 7423 15011
rect 8401 14977 8435 15011
rect 9505 14977 9539 15011
rect 13001 14977 13035 15011
rect 14565 14977 14599 15011
rect 15025 14977 15059 15011
rect 15669 14977 15703 15011
rect 16865 14977 16899 15011
rect 17049 14977 17083 15011
rect 20085 14977 20119 15011
rect 21465 14977 21499 15011
rect 24409 14977 24443 15011
rect 3157 14909 3191 14943
rect 5641 14909 5675 14943
rect 6653 14909 6687 14943
rect 7205 14909 7239 14943
rect 9597 14909 9631 14943
rect 9864 14909 9898 14943
rect 12265 14909 12299 14943
rect 12909 14909 12943 14943
rect 16313 14909 16347 14943
rect 16773 14909 16807 14943
rect 18061 14909 18095 14943
rect 18328 14909 18362 14943
rect 21281 14909 21315 14943
rect 22477 14909 22511 14943
rect 25329 14909 25363 14943
rect 25881 14909 25915 14943
rect 3402 14841 3436 14875
rect 6285 14841 6319 14875
rect 13829 14841 13863 14875
rect 14473 14841 14507 14875
rect 24225 14841 24259 14875
rect 25145 14841 25179 14875
rect 1593 14773 1627 14807
rect 2053 14773 2087 14807
rect 2881 14773 2915 14807
rect 5825 14773 5859 14807
rect 6837 14773 6871 14807
rect 7297 14773 7331 14807
rect 8217 14773 8251 14807
rect 12817 14773 12851 14807
rect 14381 14773 14415 14807
rect 16129 14773 16163 14807
rect 16405 14773 16439 14807
rect 17417 14773 17451 14807
rect 19441 14773 19475 14807
rect 20821 14773 20855 14807
rect 21373 14773 21407 14807
rect 23489 14773 23523 14807
rect 24133 14773 24167 14807
rect 3893 14569 3927 14603
rect 4537 14569 4571 14603
rect 5273 14569 5307 14603
rect 5641 14569 5675 14603
rect 8217 14569 8251 14603
rect 8769 14569 8803 14603
rect 9045 14569 9079 14603
rect 9413 14569 9447 14603
rect 10977 14569 11011 14603
rect 12725 14569 12759 14603
rect 13093 14569 13127 14603
rect 18889 14569 18923 14603
rect 22293 14569 22327 14603
rect 22845 14569 22879 14603
rect 23397 14569 23431 14603
rect 4629 14501 4663 14535
rect 6000 14501 6034 14535
rect 7665 14501 7699 14535
rect 10149 14501 10183 14535
rect 11621 14501 11655 14535
rect 14105 14501 14139 14535
rect 19625 14501 19659 14535
rect 20729 14501 20763 14535
rect 24409 14501 24443 14535
rect 1768 14433 1802 14467
rect 8033 14433 8067 14467
rect 10057 14433 10091 14467
rect 11529 14433 11563 14467
rect 13185 14433 13219 14467
rect 14473 14433 14507 14467
rect 15568 14433 15602 14467
rect 17693 14433 17727 14467
rect 18153 14433 18187 14467
rect 19349 14433 19383 14467
rect 21180 14433 21214 14467
rect 23765 14433 23799 14467
rect 24961 14433 24995 14467
rect 1501 14365 1535 14399
rect 4721 14365 4755 14399
rect 5733 14365 5767 14399
rect 11805 14365 11839 14399
rect 13277 14365 13311 14399
rect 15301 14365 15335 14399
rect 18245 14365 18279 14399
rect 18429 14365 18463 14399
rect 20913 14365 20947 14399
rect 23857 14365 23891 14399
rect 24041 14365 24075 14399
rect 25237 14365 25271 14399
rect 3525 14297 3559 14331
rect 17233 14297 17267 14331
rect 17785 14297 17819 14331
rect 2881 14229 2915 14263
rect 4169 14229 4203 14263
rect 7113 14229 7147 14263
rect 11161 14229 11195 14263
rect 12541 14229 12575 14263
rect 13829 14229 13863 14263
rect 14933 14229 14967 14263
rect 16681 14229 16715 14263
rect 19165 14229 19199 14263
rect 20085 14229 20119 14263
rect 23305 14229 23339 14263
rect 2237 14025 2271 14059
rect 2421 14025 2455 14059
rect 4721 14025 4755 14059
rect 6561 14025 6595 14059
rect 8217 14025 8251 14059
rect 10241 14025 10275 14059
rect 12449 14025 12483 14059
rect 13829 14025 13863 14059
rect 14657 14025 14691 14059
rect 15853 14025 15887 14059
rect 16405 14025 16439 14059
rect 18245 14025 18279 14059
rect 20177 14025 20211 14059
rect 20821 14025 20855 14059
rect 21281 14025 21315 14059
rect 22293 14025 22327 14059
rect 1409 13821 1443 13855
rect 1685 13821 1719 13855
rect 2605 13957 2639 13991
rect 5181 13957 5215 13991
rect 6101 13957 6135 13991
rect 6837 13957 6871 13991
rect 7849 13957 7883 13991
rect 12265 13957 12299 13991
rect 14841 13957 14875 13991
rect 17417 13957 17451 13991
rect 17877 13957 17911 13991
rect 22661 13957 22695 13991
rect 5089 13889 5123 13923
rect 5733 13889 5767 13923
rect 7297 13889 7331 13923
rect 7389 13889 7423 13923
rect 8769 13889 8803 13923
rect 11897 13889 11931 13923
rect 13093 13889 13127 13923
rect 15301 13889 15335 13923
rect 15485 13889 15519 13923
rect 16865 13889 16899 13923
rect 16957 13889 16991 13923
rect 18613 13889 18647 13923
rect 21741 13889 21775 13923
rect 21925 13889 21959 13923
rect 24225 13889 24259 13923
rect 24685 13889 24719 13923
rect 25053 13889 25087 13923
rect 25421 13889 25455 13923
rect 2697 13821 2731 13855
rect 2964 13821 2998 13855
rect 5549 13821 5583 13855
rect 5641 13821 5675 13855
rect 6009 13821 6043 13855
rect 6193 13821 6227 13855
rect 8861 13821 8895 13855
rect 9117 13821 9151 13855
rect 10885 13821 10919 13855
rect 12909 13821 12943 13855
rect 14197 13821 14231 13855
rect 16313 13821 16347 13855
rect 18797 13821 18831 13855
rect 19053 13821 19087 13855
rect 23121 13821 23155 13855
rect 24133 13821 24167 13855
rect 25237 13821 25271 13855
rect 25973 13821 26007 13855
rect 2421 13753 2455 13787
rect 7205 13753 7239 13787
rect 11345 13753 11379 13787
rect 16773 13753 16807 13787
rect 23397 13753 23431 13787
rect 24041 13753 24075 13787
rect 4077 13685 4111 13719
rect 11253 13685 11287 13719
rect 12817 13685 12851 13719
rect 13553 13685 13587 13719
rect 15209 13685 15243 13719
rect 21189 13685 21223 13719
rect 21649 13685 21683 13719
rect 23673 13685 23707 13719
rect 2053 13481 2087 13515
rect 3157 13481 3191 13515
rect 4261 13481 4295 13515
rect 4629 13481 4663 13515
rect 7481 13481 7515 13515
rect 8033 13481 8067 13515
rect 8401 13481 8435 13515
rect 8493 13481 8527 13515
rect 9045 13481 9079 13515
rect 9413 13481 9447 13515
rect 9781 13481 9815 13515
rect 14841 13481 14875 13515
rect 16681 13481 16715 13515
rect 17233 13481 17267 13515
rect 19901 13481 19935 13515
rect 20729 13481 20763 13515
rect 21925 13481 21959 13515
rect 22661 13481 22695 13515
rect 23489 13481 23523 13515
rect 25053 13481 25087 13515
rect 5816 13413 5850 13447
rect 7941 13413 7975 13447
rect 15546 13413 15580 13447
rect 18214 13413 18248 13447
rect 21373 13413 21407 13447
rect 23918 13413 23952 13447
rect 2421 13345 2455 13379
rect 2513 13345 2547 13379
rect 4077 13345 4111 13379
rect 10241 13345 10275 13379
rect 10508 13345 10542 13379
rect 12725 13345 12759 13379
rect 15301 13345 15335 13379
rect 21281 13345 21315 13379
rect 22477 13345 22511 13379
rect 23029 13345 23063 13379
rect 2605 13277 2639 13311
rect 5549 13277 5583 13311
rect 8585 13277 8619 13311
rect 17969 13277 18003 13311
rect 21465 13277 21499 13311
rect 23673 13277 23707 13311
rect 3709 13209 3743 13243
rect 6929 13209 6963 13243
rect 14013 13209 14047 13243
rect 19349 13209 19383 13243
rect 20913 13209 20947 13243
rect 1685 13141 1719 13175
rect 5273 13141 5307 13175
rect 11621 13141 11655 13175
rect 12541 13141 12575 13175
rect 17877 13141 17911 13175
rect 1961 12937 1995 12971
rect 3433 12937 3467 12971
rect 3617 12937 3651 12971
rect 4629 12937 4663 12971
rect 6193 12937 6227 12971
rect 6653 12937 6687 12971
rect 9137 12937 9171 12971
rect 10241 12937 10275 12971
rect 10793 12937 10827 12971
rect 13277 12937 13311 12971
rect 17785 12937 17819 12971
rect 18153 12937 18187 12971
rect 20821 12937 20855 12971
rect 21281 12937 21315 12971
rect 22753 12937 22787 12971
rect 3157 12869 3191 12903
rect 5181 12869 5215 12903
rect 8769 12869 8803 12903
rect 9873 12869 9907 12903
rect 19165 12869 19199 12903
rect 21189 12869 21223 12903
rect 2697 12801 2731 12835
rect 4077 12801 4111 12835
rect 4261 12801 4295 12835
rect 5825 12801 5859 12835
rect 9321 12801 9355 12835
rect 11253 12801 11287 12835
rect 11437 12801 11471 12835
rect 11805 12801 11839 12835
rect 13001 12801 13035 12835
rect 13921 12801 13955 12835
rect 14289 12801 14323 12835
rect 16957 12801 16991 12835
rect 18797 12801 18831 12835
rect 20269 12801 20303 12835
rect 21741 12801 21775 12835
rect 21925 12801 21959 12835
rect 22293 12801 22327 12835
rect 23397 12801 23431 12835
rect 2421 12733 2455 12767
rect 4997 12733 5031 12767
rect 5641 12733 5675 12767
rect 6837 12733 6871 12767
rect 7093 12733 7127 12767
rect 10517 12733 10551 12767
rect 12817 12733 12851 12767
rect 13645 12733 13679 12767
rect 18521 12733 18555 12767
rect 20177 12733 20211 12767
rect 23857 12733 23891 12767
rect 3985 12665 4019 12699
rect 13737 12665 13771 12699
rect 14534 12665 14568 12699
rect 17509 12665 17543 12699
rect 18613 12665 18647 12699
rect 23121 12665 23155 12699
rect 24124 12665 24158 12699
rect 2053 12597 2087 12631
rect 2513 12597 2547 12631
rect 5549 12597 5583 12631
rect 8217 12597 8251 12631
rect 10333 12597 10367 12631
rect 11161 12597 11195 12631
rect 12173 12597 12207 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 15669 12597 15703 12631
rect 16221 12597 16255 12631
rect 16589 12597 16623 12631
rect 19533 12597 19567 12631
rect 19717 12597 19751 12631
rect 20085 12597 20119 12631
rect 21649 12597 21683 12631
rect 25237 12597 25271 12631
rect 1409 12393 1443 12427
rect 2421 12393 2455 12427
rect 3709 12393 3743 12427
rect 4077 12393 4111 12427
rect 5549 12393 5583 12427
rect 7389 12393 7423 12427
rect 8493 12393 8527 12427
rect 9413 12393 9447 12427
rect 10793 12393 10827 12427
rect 12357 12393 12391 12427
rect 13461 12393 13495 12427
rect 15301 12393 15335 12427
rect 18429 12393 18463 12427
rect 18889 12393 18923 12427
rect 20729 12393 20763 12427
rect 21649 12393 21683 12427
rect 22753 12393 22787 12427
rect 4537 12325 4571 12359
rect 5917 12325 5951 12359
rect 6837 12325 6871 12359
rect 7849 12325 7883 12359
rect 10149 12325 10183 12359
rect 13001 12325 13035 12359
rect 13921 12325 13955 12359
rect 18245 12325 18279 12359
rect 23940 12325 23974 12359
rect 2789 12257 2823 12291
rect 2881 12257 2915 12291
rect 4445 12257 4479 12291
rect 7757 12257 7791 12291
rect 10517 12257 10551 12291
rect 11244 12257 11278 12291
rect 13829 12257 13863 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 16681 12257 16715 12291
rect 17233 12257 17267 12291
rect 17325 12257 17359 12291
rect 18797 12257 18831 12291
rect 21465 12257 21499 12291
rect 22569 12257 22603 12291
rect 2973 12189 3007 12223
rect 4721 12189 4755 12223
rect 8033 12189 8067 12223
rect 10977 12189 11011 12223
rect 13369 12189 13403 12223
rect 14013 12189 14047 12223
rect 15853 12189 15887 12223
rect 17417 12189 17451 12223
rect 18981 12189 19015 12223
rect 23673 12189 23707 12223
rect 14933 12121 14967 12155
rect 16865 12121 16899 12155
rect 2145 12053 2179 12087
rect 5181 12053 5215 12087
rect 14473 12053 14507 12087
rect 16313 12053 16347 12087
rect 19809 12053 19843 12087
rect 21281 12053 21315 12087
rect 23213 12053 23247 12087
rect 23581 12053 23615 12087
rect 25053 12053 25087 12087
rect 1593 11849 1627 11883
rect 2329 11849 2363 11883
rect 3525 11849 3559 11883
rect 5457 11849 5491 11883
rect 7481 11849 7515 11883
rect 7849 11849 7883 11883
rect 8125 11849 8159 11883
rect 10701 11849 10735 11883
rect 12449 11849 12483 11883
rect 13829 11849 13863 11883
rect 14565 11849 14599 11883
rect 16129 11849 16163 11883
rect 18429 11849 18463 11883
rect 21281 11849 21315 11883
rect 21557 11849 21591 11883
rect 21925 11849 21959 11883
rect 22293 11849 22327 11883
rect 22661 11849 22695 11883
rect 23489 11849 23523 11883
rect 23949 11849 23983 11883
rect 25697 11849 25731 11883
rect 4077 11781 4111 11815
rect 25329 11781 25363 11815
rect 3157 11713 3191 11747
rect 4721 11713 4755 11747
rect 10333 11713 10367 11747
rect 11253 11713 11287 11747
rect 11345 11713 11379 11747
rect 13093 11713 13127 11747
rect 14289 11713 14323 11747
rect 15209 11713 15243 11747
rect 16589 11713 16623 11747
rect 16773 11713 16807 11747
rect 18521 11713 18555 11747
rect 19533 11713 19567 11747
rect 24593 11713 24627 11747
rect 1409 11645 1443 11679
rect 2973 11645 3007 11679
rect 5089 11645 5123 11679
rect 14933 11645 14967 11679
rect 15945 11645 15979 11679
rect 21373 11645 21407 11679
rect 22477 11645 22511 11679
rect 25513 11645 25547 11679
rect 26065 11645 26099 11679
rect 2053 11577 2087 11611
rect 2881 11577 2915 11611
rect 4537 11577 4571 11611
rect 9965 11577 9999 11611
rect 11161 11577 11195 11611
rect 12817 11577 12851 11611
rect 13553 11577 13587 11611
rect 15025 11577 15059 11611
rect 16497 11577 16531 11611
rect 19349 11577 19383 11611
rect 24409 11577 24443 11611
rect 24961 11577 24995 11611
rect 2513 11509 2547 11543
rect 3985 11509 4019 11543
rect 4445 11509 4479 11543
rect 10793 11509 10827 11543
rect 11805 11509 11839 11543
rect 12265 11509 12299 11543
rect 12909 11509 12943 11543
rect 15577 11509 15611 11543
rect 17141 11509 17175 11543
rect 17601 11509 17635 11543
rect 18981 11509 19015 11543
rect 23029 11509 23063 11543
rect 24317 11509 24351 11543
rect 1685 11305 1719 11339
rect 2421 11305 2455 11339
rect 2513 11305 2547 11339
rect 3341 11305 3375 11339
rect 3709 11305 3743 11339
rect 4353 11305 4387 11339
rect 11069 11305 11103 11339
rect 12081 11305 12115 11339
rect 12541 11305 12575 11339
rect 14013 11305 14047 11339
rect 14749 11305 14783 11339
rect 15301 11305 15335 11339
rect 16865 11305 16899 11339
rect 18613 11305 18647 11339
rect 20913 11305 20947 11339
rect 22109 11305 22143 11339
rect 23213 11305 23247 11339
rect 24777 11305 24811 11339
rect 2973 11237 3007 11271
rect 11897 11237 11931 11271
rect 13093 11237 13127 11271
rect 15117 11237 15151 11271
rect 16405 11237 16439 11271
rect 16773 11237 16807 11271
rect 18521 11237 18555 11271
rect 2053 11169 2087 11203
rect 4629 11169 4663 11203
rect 12449 11169 12483 11203
rect 13553 11169 13587 11203
rect 15669 11169 15703 11203
rect 17233 11169 17267 11203
rect 21925 11169 21959 11203
rect 23029 11169 23063 11203
rect 24593 11169 24627 11203
rect 12725 11101 12759 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 17325 11101 17359 11135
rect 17509 11101 17543 11135
rect 24409 11101 24443 11135
rect 11621 11033 11655 11067
rect 13645 11033 13679 11067
rect 17969 11033 18003 11067
rect 10885 10965 10919 10999
rect 23949 10965 23983 10999
rect 2145 10761 2179 10795
rect 2421 10761 2455 10795
rect 2789 10761 2823 10795
rect 12725 10761 12759 10795
rect 13369 10761 13403 10795
rect 14841 10761 14875 10795
rect 15393 10761 15427 10795
rect 16405 10761 16439 10795
rect 17693 10761 17727 10795
rect 21925 10761 21959 10795
rect 23121 10761 23155 10795
rect 24777 10761 24811 10795
rect 25145 10761 25179 10795
rect 1685 10693 1719 10727
rect 3157 10693 3191 10727
rect 13645 10693 13679 10727
rect 11805 10625 11839 10659
rect 14381 10625 14415 10659
rect 15853 10625 15887 10659
rect 16037 10625 16071 10659
rect 22569 10625 22603 10659
rect 14289 10557 14323 10591
rect 24593 10557 24627 10591
rect 12817 10489 12851 10523
rect 14197 10489 14231 10523
rect 12173 10421 12207 10455
rect 13829 10421 13863 10455
rect 15301 10421 15335 10455
rect 15761 10421 15795 10455
rect 16865 10421 16899 10455
rect 17325 10421 17359 10455
rect 24409 10421 24443 10455
rect 12725 10217 12759 10251
rect 13093 10217 13127 10251
rect 13185 10217 13219 10251
rect 14933 10217 14967 10251
rect 15301 10217 15335 10251
rect 16129 10217 16163 10251
rect 22477 10217 22511 10251
rect 24777 10217 24811 10251
rect 13921 10149 13955 10183
rect 15853 10149 15887 10183
rect 14289 10081 14323 10115
rect 23489 10081 23523 10115
rect 24593 10081 24627 10115
rect 13369 10013 13403 10047
rect 14565 9945 14599 9979
rect 23673 9945 23707 9979
rect 13461 9673 13495 9707
rect 15393 9673 15427 9707
rect 23857 9673 23891 9707
rect 12817 9605 12851 9639
rect 14197 9605 14231 9639
rect 15761 9605 15795 9639
rect 25145 9605 25179 9639
rect 13185 9537 13219 9571
rect 14105 9537 14139 9571
rect 14657 9537 14691 9571
rect 14749 9537 14783 9571
rect 24409 9537 24443 9571
rect 14565 9469 14599 9503
rect 24593 9469 24627 9503
rect 24777 9333 24811 9367
rect 14197 9129 14231 9163
rect 24777 9129 24811 9163
rect 24593 8993 24627 9027
rect 24133 8585 24167 8619
rect 24961 8585 24995 8619
rect 23949 8381 23983 8415
rect 24501 8381 24535 8415
rect 24685 5865 24719 5899
rect 24501 5729 24535 5763
rect 24593 5321 24627 5355
rect 24133 4777 24167 4811
rect 24593 4709 24627 4743
rect 24501 4641 24535 4675
rect 24685 4573 24719 4607
rect 24133 4233 24167 4267
rect 24869 4097 24903 4131
rect 24593 3893 24627 3927
rect 11989 2601 12023 2635
rect 12449 2601 12483 2635
rect 14013 2601 14047 2635
rect 12878 2533 12912 2567
rect 12633 2465 12667 2499
rect 18337 2465 18371 2499
rect 18521 2329 18555 2363
rect 18981 2261 19015 2295
rect 24225 2261 24259 2295
<< metal1 >>
rect 3326 26256 3332 26308
rect 3384 26296 3390 26308
rect 4890 26296 4896 26308
rect 3384 26268 4896 26296
rect 3384 26256 3390 26268
rect 4890 26256 4896 26268
rect 4948 26256 4954 26308
rect 12986 25780 12992 25832
rect 13044 25820 13050 25832
rect 20898 25820 20904 25832
rect 13044 25792 20904 25820
rect 13044 25780 13050 25792
rect 20898 25780 20904 25792
rect 20956 25780 20962 25832
rect 11606 25712 11612 25764
rect 11664 25752 11670 25764
rect 20346 25752 20352 25764
rect 11664 25724 20352 25752
rect 11664 25712 11670 25724
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 3050 25644 3056 25696
rect 3108 25684 3114 25696
rect 7834 25684 7840 25696
rect 3108 25656 7840 25684
rect 3108 25644 3114 25656
rect 7834 25644 7840 25656
rect 7892 25644 7898 25696
rect 9490 25644 9496 25696
rect 9548 25684 9554 25696
rect 22922 25684 22928 25696
rect 9548 25656 22928 25684
rect 9548 25644 9554 25656
rect 22922 25644 22928 25656
rect 22980 25644 22986 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 4154 25440 4160 25492
rect 4212 25480 4218 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 4212 25452 4261 25480
rect 4212 25440 4218 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 7561 25483 7619 25489
rect 7561 25449 7573 25483
rect 7607 25480 7619 25483
rect 7650 25480 7656 25492
rect 7607 25452 7656 25480
rect 7607 25449 7619 25452
rect 7561 25443 7619 25449
rect 7650 25440 7656 25452
rect 7708 25440 7714 25492
rect 11606 25480 11612 25492
rect 11567 25452 11612 25480
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 12897 25483 12955 25489
rect 12897 25449 12909 25483
rect 12943 25480 12955 25483
rect 16482 25480 16488 25492
rect 12943 25452 16488 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 16482 25440 16488 25452
rect 16540 25440 16546 25492
rect 17034 25440 17040 25492
rect 17092 25480 17098 25492
rect 20073 25483 20131 25489
rect 20073 25480 20085 25483
rect 17092 25452 20085 25480
rect 17092 25440 17098 25452
rect 20073 25449 20085 25452
rect 20119 25449 20131 25483
rect 20073 25443 20131 25449
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 27614 25480 27620 25492
rect 23063 25452 27620 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 27614 25440 27620 25452
rect 27672 25440 27678 25492
rect 7466 25372 7472 25424
rect 7524 25412 7530 25424
rect 7524 25384 7788 25412
rect 7524 25372 7530 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 1443 25316 1716 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 1688 25152 1716 25316
rect 2222 25304 2228 25356
rect 2280 25344 2286 25356
rect 2501 25347 2559 25353
rect 2501 25344 2513 25347
rect 2280 25316 2513 25344
rect 2280 25304 2286 25316
rect 2501 25313 2513 25316
rect 2547 25313 2559 25347
rect 2501 25307 2559 25313
rect 3510 25304 3516 25356
rect 3568 25344 3574 25356
rect 4065 25347 4123 25353
rect 4065 25344 4077 25347
rect 3568 25316 4077 25344
rect 3568 25304 3574 25316
rect 4065 25313 4077 25316
rect 4111 25313 4123 25347
rect 4065 25307 4123 25313
rect 5074 25304 5080 25356
rect 5132 25344 5138 25356
rect 5169 25347 5227 25353
rect 5169 25344 5181 25347
rect 5132 25316 5181 25344
rect 5132 25304 5138 25316
rect 5169 25313 5181 25316
rect 5215 25313 5227 25347
rect 5169 25307 5227 25313
rect 6270 25236 6276 25288
rect 6328 25276 6334 25288
rect 7760 25285 7788 25384
rect 7834 25372 7840 25424
rect 7892 25412 7898 25424
rect 24302 25412 24308 25424
rect 7892 25384 14320 25412
rect 7892 25372 7898 25384
rect 14292 25356 14320 25384
rect 14568 25384 24308 25412
rect 10318 25344 10324 25356
rect 10279 25316 10324 25344
rect 10318 25304 10324 25316
rect 10376 25304 10382 25356
rect 11330 25304 11336 25356
rect 11388 25344 11394 25356
rect 11425 25347 11483 25353
rect 11425 25344 11437 25347
rect 11388 25316 11437 25344
rect 11388 25304 11394 25316
rect 11425 25313 11437 25316
rect 11471 25313 11483 25347
rect 12710 25344 12716 25356
rect 12671 25316 12716 25344
rect 11425 25307 11483 25313
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 14090 25304 14096 25356
rect 14148 25344 14154 25356
rect 14185 25347 14243 25353
rect 14185 25344 14197 25347
rect 14148 25316 14197 25344
rect 14148 25304 14154 25316
rect 14185 25313 14197 25316
rect 14231 25313 14243 25347
rect 14185 25307 14243 25313
rect 14274 25304 14280 25356
rect 14332 25344 14338 25356
rect 14332 25316 14377 25344
rect 14332 25304 14338 25316
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 6328 25248 7665 25276
rect 6328 25236 6334 25248
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 7745 25279 7803 25285
rect 7745 25245 7757 25279
rect 7791 25245 7803 25279
rect 7745 25239 7803 25245
rect 13998 25236 14004 25288
rect 14056 25276 14062 25288
rect 14369 25279 14427 25285
rect 14369 25276 14381 25279
rect 14056 25248 14381 25276
rect 14056 25236 14062 25248
rect 14369 25245 14381 25248
rect 14415 25245 14427 25279
rect 14369 25239 14427 25245
rect 2685 25211 2743 25217
rect 2685 25177 2697 25211
rect 2731 25208 2743 25211
rect 2774 25208 2780 25220
rect 2731 25180 2780 25208
rect 2731 25177 2743 25180
rect 2685 25171 2743 25177
rect 2774 25168 2780 25180
rect 2832 25168 2838 25220
rect 5353 25211 5411 25217
rect 5353 25177 5365 25211
rect 5399 25208 5411 25211
rect 10505 25211 10563 25217
rect 5399 25180 9536 25208
rect 5399 25177 5411 25180
rect 5353 25171 5411 25177
rect 1578 25140 1584 25152
rect 1539 25112 1584 25140
rect 1578 25100 1584 25112
rect 1636 25100 1642 25152
rect 1670 25100 1676 25152
rect 1728 25100 1734 25152
rect 2958 25100 2964 25152
rect 3016 25140 3022 25152
rect 7193 25143 7251 25149
rect 7193 25140 7205 25143
rect 3016 25112 7205 25140
rect 3016 25100 3022 25112
rect 7193 25109 7205 25112
rect 7239 25109 7251 25143
rect 7193 25103 7251 25109
rect 9122 25100 9128 25152
rect 9180 25140 9186 25152
rect 9217 25143 9275 25149
rect 9217 25140 9229 25143
rect 9180 25112 9229 25140
rect 9180 25100 9186 25112
rect 9217 25109 9229 25112
rect 9263 25109 9275 25143
rect 9508 25140 9536 25180
rect 10505 25177 10517 25211
rect 10551 25208 10563 25211
rect 12986 25208 12992 25220
rect 10551 25180 12992 25208
rect 10551 25177 10563 25180
rect 10505 25171 10563 25177
rect 12986 25168 12992 25180
rect 13044 25168 13050 25220
rect 13188 25180 13952 25208
rect 13188 25140 13216 25180
rect 13354 25140 13360 25152
rect 9508 25112 13216 25140
rect 13315 25112 13360 25140
rect 9217 25103 9275 25109
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 13814 25140 13820 25152
rect 13775 25112 13820 25140
rect 13814 25100 13820 25112
rect 13872 25100 13878 25152
rect 13924 25140 13952 25180
rect 14568 25140 14596 25384
rect 24302 25372 24308 25384
rect 24360 25372 24366 25424
rect 16117 25347 16175 25353
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 16390 25344 16396 25356
rect 16163 25316 16396 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 17862 25304 17868 25356
rect 17920 25344 17926 25356
rect 18693 25347 18751 25353
rect 18693 25344 18705 25347
rect 17920 25316 18705 25344
rect 17920 25304 17926 25316
rect 18693 25313 18705 25316
rect 18739 25313 18751 25347
rect 18693 25307 18751 25313
rect 18785 25347 18843 25353
rect 18785 25313 18797 25347
rect 18831 25344 18843 25347
rect 19150 25344 19156 25356
rect 18831 25316 19156 25344
rect 18831 25313 18843 25316
rect 18785 25307 18843 25313
rect 19150 25304 19156 25316
rect 19208 25304 19214 25356
rect 19889 25347 19947 25353
rect 19889 25313 19901 25347
rect 19935 25344 19947 25347
rect 20438 25344 20444 25356
rect 19935 25316 20444 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 20438 25304 20444 25316
rect 20496 25304 20502 25356
rect 21542 25344 21548 25356
rect 21503 25316 21548 25344
rect 21542 25304 21548 25316
rect 21600 25304 21606 25356
rect 24581 25347 24639 25353
rect 24581 25313 24593 25347
rect 24627 25344 24639 25347
rect 25038 25344 25044 25356
rect 24627 25316 25044 25344
rect 24627 25313 24639 25316
rect 24581 25307 24639 25313
rect 25038 25304 25044 25316
rect 25096 25304 25102 25356
rect 16206 25276 16212 25288
rect 16167 25248 16212 25276
rect 16206 25236 16212 25248
rect 16264 25236 16270 25288
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 17773 25279 17831 25285
rect 17773 25245 17785 25279
rect 17819 25276 17831 25279
rect 18874 25276 18880 25288
rect 17819 25248 18736 25276
rect 18835 25248 18880 25276
rect 17819 25245 17831 25248
rect 17773 25239 17831 25245
rect 15289 25211 15347 25217
rect 15289 25177 15301 25211
rect 15335 25208 15347 25211
rect 15930 25208 15936 25220
rect 15335 25180 15936 25208
rect 15335 25177 15347 25180
rect 15289 25171 15347 25177
rect 15930 25168 15936 25180
rect 15988 25208 15994 25220
rect 16316 25208 16344 25239
rect 16758 25208 16764 25220
rect 15988 25180 16764 25208
rect 15988 25168 15994 25180
rect 16758 25168 16764 25180
rect 16816 25168 16822 25220
rect 18141 25211 18199 25217
rect 18141 25177 18153 25211
rect 18187 25208 18199 25211
rect 18598 25208 18604 25220
rect 18187 25180 18604 25208
rect 18187 25177 18199 25180
rect 18141 25171 18199 25177
rect 18598 25168 18604 25180
rect 18656 25168 18662 25220
rect 18708 25208 18736 25248
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 21174 25236 21180 25288
rect 21232 25276 21238 25288
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 21232 25248 21649 25276
rect 21232 25236 21238 25248
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 21637 25239 21695 25245
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25276 21879 25279
rect 23014 25276 23020 25288
rect 21867 25248 23020 25276
rect 21867 25245 21879 25248
rect 21821 25239 21879 25245
rect 23014 25236 23020 25248
rect 23072 25236 23078 25288
rect 18966 25208 18972 25220
rect 18708 25180 18972 25208
rect 18966 25168 18972 25180
rect 19024 25208 19030 25220
rect 24762 25208 24768 25220
rect 19024 25180 21220 25208
rect 24723 25180 24768 25208
rect 19024 25168 19030 25180
rect 14826 25140 14832 25152
rect 13924 25112 14596 25140
rect 14787 25112 14832 25140
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15746 25140 15752 25152
rect 15707 25112 15752 25140
rect 15746 25100 15752 25112
rect 15804 25100 15810 25152
rect 17034 25100 17040 25152
rect 17092 25140 17098 25152
rect 18325 25143 18383 25149
rect 18325 25140 18337 25143
rect 17092 25112 18337 25140
rect 17092 25100 17098 25112
rect 18325 25109 18337 25112
rect 18371 25109 18383 25143
rect 18325 25103 18383 25109
rect 19705 25143 19763 25149
rect 19705 25109 19717 25143
rect 19751 25140 19763 25143
rect 20070 25140 20076 25152
rect 19751 25112 20076 25140
rect 19751 25109 19763 25112
rect 19705 25103 19763 25109
rect 20070 25100 20076 25112
rect 20128 25100 20134 25152
rect 20993 25143 21051 25149
rect 20993 25109 21005 25143
rect 21039 25140 21051 25143
rect 21082 25140 21088 25152
rect 21039 25112 21088 25140
rect 21039 25109 21051 25112
rect 20993 25103 21051 25109
rect 21082 25100 21088 25112
rect 21140 25100 21146 25152
rect 21192 25149 21220 25180
rect 24762 25168 24768 25180
rect 24820 25168 24826 25220
rect 21177 25143 21235 25149
rect 21177 25109 21189 25143
rect 21223 25109 21235 25143
rect 21177 25103 21235 25109
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3786 24936 3792 24948
rect 3747 24908 3792 24936
rect 3786 24896 3792 24908
rect 3844 24896 3850 24948
rect 4890 24936 4896 24948
rect 4851 24908 4896 24936
rect 4890 24896 4896 24908
rect 4948 24896 4954 24948
rect 12250 24936 12256 24948
rect 12163 24908 12256 24936
rect 12250 24896 12256 24908
rect 12308 24936 12314 24948
rect 12308 24908 13676 24936
rect 12308 24896 12314 24908
rect 7650 24868 7656 24880
rect 6840 24840 7656 24868
rect 4249 24803 4307 24809
rect 4249 24769 4261 24803
rect 4295 24800 4307 24803
rect 4890 24800 4896 24812
rect 4295 24772 4896 24800
rect 4295 24769 4307 24772
rect 4249 24763 4307 24769
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 2038 24732 2044 24744
rect 1443 24704 2044 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 2038 24692 2044 24704
rect 2096 24692 2102 24744
rect 2501 24735 2559 24741
rect 2501 24701 2513 24735
rect 2547 24732 2559 24735
rect 3145 24735 3203 24741
rect 3145 24732 3157 24735
rect 2547 24704 3157 24732
rect 2547 24701 2559 24704
rect 2501 24695 2559 24701
rect 3145 24701 3157 24704
rect 3191 24732 3203 24735
rect 3418 24732 3424 24744
rect 3191 24704 3424 24732
rect 3191 24701 3203 24704
rect 3145 24695 3203 24701
rect 3418 24692 3424 24704
rect 3476 24692 3482 24744
rect 3605 24735 3663 24741
rect 3605 24701 3617 24735
rect 3651 24732 3663 24735
rect 4264 24732 4292 24763
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 6273 24803 6331 24809
rect 6273 24769 6285 24803
rect 6319 24800 6331 24803
rect 6840 24800 6868 24840
rect 7650 24828 7656 24840
rect 7708 24828 7714 24880
rect 9122 24828 9128 24880
rect 9180 24868 9186 24880
rect 9180 24840 9812 24868
rect 9180 24828 9186 24840
rect 9784 24809 9812 24840
rect 6319 24772 6868 24800
rect 8297 24803 8355 24809
rect 6319 24769 6331 24772
rect 6273 24763 6331 24769
rect 8297 24769 8309 24803
rect 8343 24800 8355 24803
rect 9769 24803 9827 24809
rect 8343 24772 8800 24800
rect 8343 24769 8355 24772
rect 8297 24763 8355 24769
rect 3651 24704 4292 24732
rect 4709 24735 4767 24741
rect 3651 24701 3663 24704
rect 3605 24695 3663 24701
rect 4709 24701 4721 24735
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 4724 24608 4752 24695
rect 8021 24667 8079 24673
rect 8021 24633 8033 24667
rect 8067 24664 8079 24667
rect 8202 24664 8208 24676
rect 8067 24636 8208 24664
rect 8067 24633 8079 24636
rect 8021 24627 8079 24633
rect 8202 24624 8208 24636
rect 8260 24624 8266 24676
rect 8772 24608 8800 24772
rect 9769 24769 9781 24803
rect 9815 24769 9827 24803
rect 9769 24763 9827 24769
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 13538 24800 13544 24812
rect 12584 24772 13544 24800
rect 12584 24760 12590 24772
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 13648 24809 13676 24908
rect 18782 24896 18788 24948
rect 18840 24936 18846 24948
rect 21542 24936 21548 24948
rect 18840 24908 21548 24936
rect 18840 24896 18846 24908
rect 21542 24896 21548 24908
rect 21600 24936 21606 24948
rect 22189 24939 22247 24945
rect 22189 24936 22201 24939
rect 21600 24908 22201 24936
rect 21600 24896 21606 24908
rect 22189 24905 22201 24908
rect 22235 24905 22247 24939
rect 22189 24899 22247 24905
rect 24670 24896 24676 24948
rect 24728 24936 24734 24948
rect 24765 24939 24823 24945
rect 24765 24936 24777 24939
rect 24728 24908 24777 24936
rect 24728 24896 24734 24908
rect 24765 24905 24777 24908
rect 24811 24905 24823 24939
rect 24765 24899 24823 24905
rect 15746 24828 15752 24880
rect 15804 24868 15810 24880
rect 20898 24868 20904 24880
rect 15804 24840 20904 24868
rect 15804 24828 15810 24840
rect 20898 24828 20904 24840
rect 20956 24828 20962 24880
rect 21082 24828 21088 24880
rect 21140 24868 21146 24880
rect 21910 24868 21916 24880
rect 21140 24840 21916 24868
rect 21140 24828 21146 24840
rect 13633 24803 13691 24809
rect 13633 24769 13645 24803
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 14458 24760 14464 24812
rect 14516 24800 14522 24812
rect 15197 24803 15255 24809
rect 15197 24800 15209 24803
rect 14516 24772 15209 24800
rect 14516 24760 14522 24772
rect 15197 24769 15209 24772
rect 15243 24769 15255 24803
rect 16758 24800 16764 24812
rect 16719 24772 16764 24800
rect 15197 24763 15255 24769
rect 16758 24760 16764 24772
rect 16816 24800 16822 24812
rect 17221 24803 17279 24809
rect 17221 24800 17233 24803
rect 16816 24772 17233 24800
rect 16816 24760 16822 24772
rect 17221 24769 17233 24772
rect 17267 24769 17279 24803
rect 18598 24800 18604 24812
rect 18559 24772 18604 24800
rect 17221 24763 17279 24769
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 19521 24803 19579 24809
rect 19521 24769 19533 24803
rect 19567 24800 19579 24803
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 19567 24772 20177 24800
rect 19567 24769 19579 24772
rect 19521 24763 19579 24769
rect 20165 24769 20177 24772
rect 20211 24800 20223 24803
rect 20346 24800 20352 24812
rect 20211 24772 20352 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20990 24760 20996 24812
rect 21048 24800 21054 24812
rect 21744 24809 21772 24840
rect 21910 24828 21916 24840
rect 21968 24828 21974 24880
rect 21637 24803 21695 24809
rect 21637 24800 21649 24803
rect 21048 24772 21649 24800
rect 21048 24760 21054 24772
rect 21637 24769 21649 24772
rect 21683 24769 21695 24803
rect 21637 24763 21695 24769
rect 21729 24803 21787 24809
rect 21729 24769 21741 24803
rect 21775 24769 21787 24803
rect 21729 24763 21787 24769
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22738 24800 22744 24812
rect 22152 24772 22744 24800
rect 22152 24760 22158 24772
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 9582 24692 9588 24744
rect 9640 24732 9646 24744
rect 9677 24735 9735 24741
rect 9677 24732 9689 24735
rect 9640 24704 9689 24732
rect 9640 24692 9646 24704
rect 9677 24701 9689 24704
rect 9723 24701 9735 24735
rect 11241 24735 11299 24741
rect 11241 24732 11253 24735
rect 9677 24695 9735 24701
rect 11164 24704 11253 24732
rect 9490 24664 9496 24676
rect 9048 24636 9496 24664
rect 9048 24608 9076 24636
rect 9490 24624 9496 24636
rect 9548 24664 9554 24676
rect 9548 24636 9628 24664
rect 9548 24624 9554 24636
rect 1394 24556 1400 24608
rect 1452 24596 1458 24608
rect 1581 24599 1639 24605
rect 1581 24596 1593 24599
rect 1452 24568 1593 24596
rect 1452 24556 1458 24568
rect 1581 24565 1593 24568
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 1670 24556 1676 24608
rect 1728 24596 1734 24608
rect 1949 24599 2007 24605
rect 1949 24596 1961 24599
rect 1728 24568 1961 24596
rect 1728 24556 1734 24568
rect 1949 24565 1961 24568
rect 1995 24565 2007 24599
rect 1949 24559 2007 24565
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2317 24599 2375 24605
rect 2317 24596 2329 24599
rect 2280 24568 2329 24596
rect 2280 24556 2286 24568
rect 2317 24565 2329 24568
rect 2363 24565 2375 24599
rect 2682 24596 2688 24608
rect 2643 24568 2688 24596
rect 2317 24559 2375 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 3510 24596 3516 24608
rect 3471 24568 3516 24596
rect 3510 24556 3516 24568
rect 3568 24556 3574 24608
rect 4617 24599 4675 24605
rect 4617 24565 4629 24599
rect 4663 24596 4675 24599
rect 4706 24596 4712 24608
rect 4663 24568 4712 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5074 24556 5080 24608
rect 5132 24596 5138 24608
rect 5261 24599 5319 24605
rect 5261 24596 5273 24599
rect 5132 24568 5273 24596
rect 5132 24556 5138 24568
rect 5261 24565 5273 24568
rect 5307 24565 5319 24599
rect 5261 24559 5319 24565
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 6549 24599 6607 24605
rect 6549 24596 6561 24599
rect 6328 24568 6561 24596
rect 6328 24556 6334 24568
rect 6549 24565 6561 24568
rect 6595 24565 6607 24599
rect 6549 24559 6607 24565
rect 7285 24599 7343 24605
rect 7285 24565 7297 24599
rect 7331 24596 7343 24599
rect 7466 24596 7472 24608
rect 7331 24568 7472 24596
rect 7331 24565 7343 24568
rect 7285 24559 7343 24565
rect 7466 24556 7472 24568
rect 7524 24556 7530 24608
rect 7650 24596 7656 24608
rect 7611 24568 7656 24596
rect 7650 24556 7656 24568
rect 7708 24556 7714 24608
rect 8110 24596 8116 24608
rect 8071 24568 8116 24596
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8754 24596 8760 24608
rect 8715 24568 8760 24596
rect 8754 24556 8760 24568
rect 8812 24556 8818 24608
rect 9030 24596 9036 24608
rect 8991 24568 9036 24596
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 9214 24596 9220 24608
rect 9175 24568 9220 24596
rect 9214 24556 9220 24568
rect 9272 24556 9278 24608
rect 9600 24605 9628 24636
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 10413 24667 10471 24673
rect 10413 24664 10425 24667
rect 10376 24636 10425 24664
rect 10376 24624 10382 24636
rect 10413 24633 10425 24636
rect 10459 24664 10471 24667
rect 10778 24664 10784 24676
rect 10459 24636 10784 24664
rect 10459 24633 10471 24636
rect 10413 24627 10471 24633
rect 10778 24624 10784 24636
rect 10836 24624 10842 24676
rect 11164 24608 11192 24704
rect 11241 24701 11253 24704
rect 11287 24701 11299 24735
rect 13354 24732 13360 24744
rect 11241 24695 11299 24701
rect 12912 24704 13360 24732
rect 12066 24624 12072 24676
rect 12124 24664 12130 24676
rect 12912 24664 12940 24704
rect 13354 24692 13360 24704
rect 13412 24732 13418 24744
rect 13449 24735 13507 24741
rect 13449 24732 13461 24735
rect 13412 24704 13461 24732
rect 13412 24692 13418 24704
rect 13449 24701 13461 24704
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 15838 24692 15844 24744
rect 15896 24732 15902 24744
rect 16669 24735 16727 24741
rect 16669 24732 16681 24735
rect 15896 24704 16681 24732
rect 15896 24692 15902 24704
rect 16669 24701 16681 24704
rect 16715 24732 16727 24735
rect 17678 24732 17684 24744
rect 16715 24704 17684 24732
rect 16715 24701 16727 24704
rect 16669 24695 16727 24701
rect 17678 24692 17684 24704
rect 17736 24692 17742 24744
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24732 18475 24735
rect 18966 24732 18972 24744
rect 18463 24704 18972 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 18966 24692 18972 24704
rect 19024 24692 19030 24744
rect 21085 24735 21143 24741
rect 21085 24701 21097 24735
rect 21131 24732 21143 24735
rect 21174 24732 21180 24744
rect 21131 24704 21180 24732
rect 21131 24701 21143 24704
rect 21085 24695 21143 24701
rect 21174 24692 21180 24704
rect 21232 24692 21238 24744
rect 22186 24692 22192 24744
rect 22244 24732 22250 24744
rect 23198 24732 23204 24744
rect 22244 24704 23204 24732
rect 22244 24692 22250 24704
rect 23198 24692 23204 24704
rect 23256 24692 23262 24744
rect 24581 24735 24639 24741
rect 24581 24732 24593 24735
rect 24412 24704 24593 24732
rect 12124 24636 12940 24664
rect 12989 24667 13047 24673
rect 12124 24624 12130 24636
rect 12989 24633 13001 24667
rect 13035 24664 13047 24667
rect 13035 24636 13492 24664
rect 13035 24633 13047 24636
rect 12989 24627 13047 24633
rect 13464 24608 13492 24636
rect 14826 24624 14832 24676
rect 14884 24664 14890 24676
rect 15105 24667 15163 24673
rect 15105 24664 15117 24667
rect 14884 24636 15117 24664
rect 14884 24624 14890 24636
rect 15105 24633 15117 24636
rect 15151 24633 15163 24667
rect 15105 24627 15163 24633
rect 15749 24667 15807 24673
rect 15749 24633 15761 24667
rect 15795 24664 15807 24667
rect 16390 24664 16396 24676
rect 15795 24636 16396 24664
rect 15795 24633 15807 24636
rect 15749 24627 15807 24633
rect 16390 24624 16396 24636
rect 16448 24624 16454 24676
rect 19150 24664 19156 24676
rect 19111 24636 19156 24664
rect 19150 24624 19156 24636
rect 19208 24624 19214 24676
rect 19981 24667 20039 24673
rect 19981 24633 19993 24667
rect 20027 24664 20039 24667
rect 20162 24664 20168 24676
rect 20027 24636 20168 24664
rect 20027 24633 20039 24636
rect 19981 24627 20039 24633
rect 20162 24624 20168 24636
rect 20220 24664 20226 24676
rect 22557 24667 22615 24673
rect 22557 24664 22569 24667
rect 20220 24636 21220 24664
rect 20220 24624 20226 24636
rect 9585 24599 9643 24605
rect 9585 24565 9597 24599
rect 9631 24565 9643 24599
rect 10686 24596 10692 24608
rect 10647 24568 10692 24596
rect 9585 24559 9643 24565
rect 10686 24556 10692 24568
rect 10744 24556 10750 24608
rect 11146 24596 11152 24608
rect 11107 24568 11152 24596
rect 11146 24556 11152 24568
rect 11204 24556 11210 24608
rect 11422 24596 11428 24608
rect 11383 24568 11428 24596
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 11885 24599 11943 24605
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 12710 24596 12716 24608
rect 11931 24568 12716 24596
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 13081 24599 13139 24605
rect 13081 24565 13093 24599
rect 13127 24596 13139 24599
rect 13354 24596 13360 24608
rect 13127 24568 13360 24596
rect 13127 24565 13139 24568
rect 13081 24559 13139 24565
rect 13354 24556 13360 24568
rect 13412 24556 13418 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 13504 24568 13553 24596
rect 13504 24556 13510 24568
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 13541 24559 13599 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14274 24556 14280 24608
rect 14332 24596 14338 24608
rect 14461 24599 14519 24605
rect 14461 24596 14473 24599
rect 14332 24568 14473 24596
rect 14332 24556 14338 24568
rect 14461 24565 14473 24568
rect 14507 24565 14519 24599
rect 14461 24559 14519 24565
rect 14550 24556 14556 24608
rect 14608 24596 14614 24608
rect 14645 24599 14703 24605
rect 14645 24596 14657 24599
rect 14608 24568 14657 24596
rect 14608 24556 14614 24568
rect 14645 24565 14657 24568
rect 14691 24565 14703 24599
rect 14645 24559 14703 24565
rect 14734 24556 14740 24608
rect 14792 24596 14798 24608
rect 15013 24599 15071 24605
rect 15013 24596 15025 24599
rect 14792 24568 15025 24596
rect 14792 24556 14798 24568
rect 15013 24565 15025 24568
rect 15059 24565 15071 24599
rect 15013 24559 15071 24565
rect 15838 24556 15844 24608
rect 15896 24596 15902 24608
rect 16025 24599 16083 24605
rect 16025 24596 16037 24599
rect 15896 24568 16037 24596
rect 15896 24556 15902 24568
rect 16025 24565 16037 24568
rect 16071 24565 16083 24599
rect 16025 24559 16083 24565
rect 16114 24556 16120 24608
rect 16172 24596 16178 24608
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 16172 24568 16221 24596
rect 16172 24556 16178 24568
rect 16209 24565 16221 24568
rect 16255 24565 16267 24599
rect 16209 24559 16267 24565
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 16577 24599 16635 24605
rect 16577 24596 16589 24599
rect 16356 24568 16589 24596
rect 16356 24556 16362 24568
rect 16577 24565 16589 24568
rect 16623 24565 16635 24599
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 16577 24559 16635 24565
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18509 24599 18567 24605
rect 18509 24565 18521 24599
rect 18555 24596 18567 24599
rect 18966 24596 18972 24608
rect 18555 24568 18972 24596
rect 18555 24565 18567 24568
rect 18509 24559 18567 24565
rect 18966 24556 18972 24568
rect 19024 24556 19030 24608
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19576 24568 19625 24596
rect 19576 24556 19582 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 20070 24596 20076 24608
rect 20031 24568 20076 24596
rect 19613 24559 19671 24565
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20717 24599 20775 24605
rect 20717 24565 20729 24599
rect 20763 24596 20775 24599
rect 20990 24596 20996 24608
rect 20763 24568 20996 24596
rect 20763 24565 20775 24568
rect 20717 24559 20775 24565
rect 20990 24556 20996 24568
rect 21048 24556 21054 24608
rect 21192 24605 21220 24636
rect 21560 24636 22569 24664
rect 21177 24599 21235 24605
rect 21177 24565 21189 24599
rect 21223 24565 21235 24599
rect 21177 24559 21235 24565
rect 21358 24556 21364 24608
rect 21416 24596 21422 24608
rect 21560 24605 21588 24636
rect 22557 24633 22569 24636
rect 22603 24633 22615 24667
rect 22557 24627 22615 24633
rect 21545 24599 21603 24605
rect 21545 24596 21557 24599
rect 21416 24568 21557 24596
rect 21416 24556 21422 24568
rect 21545 24565 21557 24568
rect 21591 24565 21603 24599
rect 23014 24596 23020 24608
rect 22927 24568 23020 24596
rect 21545 24559 21603 24565
rect 23014 24556 23020 24568
rect 23072 24596 23078 24608
rect 23198 24596 23204 24608
rect 23072 24568 23204 24596
rect 23072 24556 23078 24568
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 23474 24556 23480 24608
rect 23532 24596 23538 24608
rect 24412 24605 24440 24704
rect 24581 24701 24593 24704
rect 24627 24701 24639 24735
rect 24581 24695 24639 24701
rect 24397 24599 24455 24605
rect 24397 24596 24409 24599
rect 23532 24568 24409 24596
rect 23532 24556 23538 24568
rect 24397 24565 24409 24568
rect 24443 24565 24455 24599
rect 24397 24559 24455 24565
rect 24854 24556 24860 24608
rect 24912 24596 24918 24608
rect 25038 24596 25044 24608
rect 24912 24568 25044 24596
rect 24912 24556 24918 24568
rect 25038 24556 25044 24568
rect 25096 24596 25102 24608
rect 25133 24599 25191 24605
rect 25133 24596 25145 24599
rect 25096 24568 25145 24596
rect 25096 24556 25102 24568
rect 25133 24565 25145 24568
rect 25179 24565 25191 24599
rect 25133 24559 25191 24565
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 290 24352 296 24404
rect 348 24392 354 24404
rect 1302 24392 1308 24404
rect 348 24364 1308 24392
rect 348 24352 354 24364
rect 1302 24352 1308 24364
rect 1360 24352 1366 24404
rect 4154 24352 4160 24404
rect 4212 24392 4218 24404
rect 4249 24395 4307 24401
rect 4249 24392 4261 24395
rect 4212 24364 4261 24392
rect 4212 24352 4218 24364
rect 4249 24361 4261 24364
rect 4295 24361 4307 24395
rect 4249 24355 4307 24361
rect 6362 24352 6368 24404
rect 6420 24392 6426 24404
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 6420 24364 7665 24392
rect 6420 24352 6426 24364
rect 7653 24361 7665 24364
rect 7699 24392 7711 24395
rect 8110 24392 8116 24404
rect 7699 24364 8116 24392
rect 7699 24361 7711 24364
rect 7653 24355 7711 24361
rect 8110 24352 8116 24364
rect 8168 24352 8174 24404
rect 9674 24392 9680 24404
rect 9635 24364 9680 24392
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 13998 24392 14004 24404
rect 13959 24364 14004 24392
rect 13998 24352 14004 24364
rect 14056 24352 14062 24404
rect 18414 24352 18420 24404
rect 18472 24392 18478 24404
rect 18601 24395 18659 24401
rect 18601 24392 18613 24395
rect 18472 24364 18613 24392
rect 18472 24352 18478 24364
rect 18601 24361 18613 24364
rect 18647 24392 18659 24395
rect 18874 24392 18880 24404
rect 18647 24364 18880 24392
rect 18647 24361 18659 24364
rect 18601 24355 18659 24361
rect 18874 24352 18880 24364
rect 18932 24352 18938 24404
rect 20162 24392 20168 24404
rect 20123 24364 20168 24392
rect 20162 24352 20168 24364
rect 20220 24352 20226 24404
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 24946 24352 24952 24404
rect 25004 24392 25010 24404
rect 25958 24392 25964 24404
rect 25004 24364 25964 24392
rect 25004 24352 25010 24364
rect 25958 24352 25964 24364
rect 26016 24352 26022 24404
rect 9309 24327 9367 24333
rect 9309 24293 9321 24327
rect 9355 24324 9367 24327
rect 9582 24324 9588 24336
rect 9355 24296 9588 24324
rect 9355 24293 9367 24296
rect 9309 24287 9367 24293
rect 9582 24284 9588 24296
rect 9640 24284 9646 24336
rect 17678 24284 17684 24336
rect 17736 24324 17742 24336
rect 21545 24327 21603 24333
rect 21545 24324 21557 24327
rect 17736 24296 21557 24324
rect 17736 24284 17742 24296
rect 21545 24293 21557 24296
rect 21591 24324 21603 24327
rect 21818 24324 21824 24336
rect 21591 24296 21824 24324
rect 21591 24293 21603 24296
rect 21545 24287 21603 24293
rect 21818 24284 21824 24296
rect 21876 24284 21882 24336
rect 22278 24284 22284 24336
rect 22336 24324 22342 24336
rect 23109 24327 23167 24333
rect 23109 24324 23121 24327
rect 22336 24296 23121 24324
rect 22336 24284 22342 24296
rect 23109 24293 23121 24296
rect 23155 24293 23167 24327
rect 23109 24287 23167 24293
rect 1397 24259 1455 24265
rect 1397 24225 1409 24259
rect 1443 24256 1455 24259
rect 1946 24256 1952 24268
rect 1443 24228 1952 24256
rect 1443 24225 1455 24228
rect 1397 24219 1455 24225
rect 1946 24216 1952 24228
rect 2004 24216 2010 24268
rect 2498 24256 2504 24268
rect 2459 24228 2504 24256
rect 2498 24216 2504 24228
rect 2556 24216 2562 24268
rect 3786 24216 3792 24268
rect 3844 24256 3850 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 3844 24228 4077 24256
rect 3844 24216 3850 24228
rect 4065 24225 4077 24228
rect 4111 24256 4123 24259
rect 4617 24259 4675 24265
rect 4617 24256 4629 24259
rect 4111 24228 4629 24256
rect 4111 24225 4123 24228
rect 4065 24219 4123 24225
rect 4617 24225 4629 24228
rect 4663 24225 4675 24259
rect 4617 24219 4675 24225
rect 5988 24259 6046 24265
rect 5988 24225 6000 24259
rect 6034 24256 6046 24259
rect 6362 24256 6368 24268
rect 6034 24228 6368 24256
rect 6034 24225 6046 24228
rect 5988 24219 6046 24225
rect 6362 24216 6368 24228
rect 6420 24216 6426 24268
rect 8478 24256 8484 24268
rect 8439 24228 8484 24256
rect 8478 24216 8484 24228
rect 8536 24216 8542 24268
rect 9858 24216 9864 24268
rect 9916 24256 9922 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9916 24228 10057 24256
rect 9916 24216 9922 24228
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 10045 24219 10103 24225
rect 11333 24259 11391 24265
rect 11333 24225 11345 24259
rect 11379 24256 11391 24259
rect 12989 24259 13047 24265
rect 11379 24228 12204 24256
rect 11379 24225 11391 24228
rect 11333 24219 11391 24225
rect 2038 24188 2044 24200
rect 1999 24160 2044 24188
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24188 5687 24191
rect 5721 24191 5779 24197
rect 5721 24188 5733 24191
rect 5675 24160 5733 24188
rect 5675 24157 5687 24160
rect 5629 24151 5687 24157
rect 5721 24157 5733 24160
rect 5767 24157 5779 24191
rect 5721 24151 5779 24157
rect 1486 24012 1492 24064
rect 1544 24052 1550 24064
rect 1581 24055 1639 24061
rect 1581 24052 1593 24055
rect 1544 24024 1593 24052
rect 1544 24012 1550 24024
rect 1581 24021 1593 24024
rect 1627 24021 1639 24055
rect 1581 24015 1639 24021
rect 2685 24055 2743 24061
rect 2685 24021 2697 24055
rect 2731 24052 2743 24055
rect 2774 24052 2780 24064
rect 2731 24024 2780 24052
rect 2731 24021 2743 24024
rect 2685 24015 2743 24021
rect 2774 24012 2780 24024
rect 2832 24012 2838 24064
rect 3602 24012 3608 24064
rect 3660 24052 3666 24064
rect 3697 24055 3755 24061
rect 3697 24052 3709 24055
rect 3660 24024 3709 24052
rect 3660 24012 3666 24024
rect 3697 24021 3709 24024
rect 3743 24052 3755 24055
rect 4154 24052 4160 24064
rect 3743 24024 4160 24052
rect 3743 24021 3755 24024
rect 3697 24015 3755 24021
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 5258 24052 5264 24064
rect 5219 24024 5264 24052
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 5736 24052 5764 24151
rect 9950 24148 9956 24200
rect 10008 24188 10014 24200
rect 10137 24191 10195 24197
rect 10137 24188 10149 24191
rect 10008 24160 10149 24188
rect 10008 24148 10014 24160
rect 10137 24157 10149 24160
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24157 10287 24191
rect 11514 24188 11520 24200
rect 11475 24160 11520 24188
rect 10229 24151 10287 24157
rect 10042 24080 10048 24132
rect 10100 24120 10106 24132
rect 10244 24120 10272 24151
rect 11514 24148 11520 24160
rect 11572 24148 11578 24200
rect 10689 24123 10747 24129
rect 10689 24120 10701 24123
rect 10100 24092 10701 24120
rect 10100 24080 10106 24092
rect 10689 24089 10701 24092
rect 10735 24089 10747 24123
rect 10689 24083 10747 24089
rect 6086 24052 6092 24064
rect 5736 24024 6092 24052
rect 6086 24012 6092 24024
rect 6144 24012 6150 24064
rect 6822 24012 6828 24064
rect 6880 24052 6886 24064
rect 7101 24055 7159 24061
rect 7101 24052 7113 24055
rect 6880 24024 7113 24052
rect 6880 24012 6886 24024
rect 7101 24021 7113 24024
rect 7147 24021 7159 24055
rect 7101 24015 7159 24021
rect 8113 24055 8171 24061
rect 8113 24021 8125 24055
rect 8159 24052 8171 24055
rect 8202 24052 8208 24064
rect 8159 24024 8208 24052
rect 8159 24021 8171 24024
rect 8113 24015 8171 24021
rect 8202 24012 8208 24024
rect 8260 24012 8266 24064
rect 8662 24052 8668 24064
rect 8623 24024 8668 24052
rect 8662 24012 8668 24024
rect 8720 24012 8726 24064
rect 11054 24052 11060 24064
rect 11015 24024 11060 24052
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 12176 24061 12204 24228
rect 12989 24225 13001 24259
rect 13035 24256 13047 24259
rect 13354 24256 13360 24268
rect 13035 24228 13360 24256
rect 13035 24225 13047 24228
rect 12989 24219 13047 24225
rect 13354 24216 13360 24228
rect 13412 24216 13418 24268
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 16666 24216 16672 24268
rect 16724 24256 16730 24268
rect 16833 24259 16891 24265
rect 16833 24256 16845 24259
rect 16724 24228 16845 24256
rect 16724 24216 16730 24228
rect 16833 24225 16845 24228
rect 16879 24225 16891 24259
rect 19426 24256 19432 24268
rect 19387 24228 19432 24256
rect 16833 24219 16891 24225
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 20714 24216 20720 24268
rect 20772 24256 20778 24268
rect 21453 24259 21511 24265
rect 21453 24256 21465 24259
rect 20772 24228 21465 24256
rect 20772 24216 20778 24228
rect 21453 24225 21465 24228
rect 21499 24225 21511 24259
rect 23014 24256 23020 24268
rect 22975 24228 23020 24256
rect 21453 24219 21511 24225
rect 23014 24216 23020 24228
rect 23072 24216 23078 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 13081 24191 13139 24197
rect 13081 24188 13093 24191
rect 13004 24160 13093 24188
rect 13004 24132 13032 24160
rect 13081 24157 13093 24160
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 14185 24191 14243 24197
rect 14185 24157 14197 24191
rect 14231 24188 14243 24191
rect 14642 24188 14648 24200
rect 14231 24160 14648 24188
rect 14231 24157 14243 24160
rect 14185 24151 14243 24157
rect 12529 24123 12587 24129
rect 12529 24089 12541 24123
rect 12575 24120 12587 24123
rect 12802 24120 12808 24132
rect 12575 24092 12808 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 12802 24080 12808 24092
rect 12860 24080 12866 24132
rect 12986 24080 12992 24132
rect 13044 24080 13050 24132
rect 12161 24055 12219 24061
rect 12161 24021 12173 24055
rect 12207 24052 12219 24055
rect 12342 24052 12348 24064
rect 12207 24024 12348 24052
rect 12207 24021 12219 24024
rect 12161 24015 12219 24021
rect 12342 24012 12348 24024
rect 12400 24012 12406 24064
rect 12618 24052 12624 24064
rect 12579 24024 12624 24052
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12820 24052 12848 24080
rect 13188 24052 13216 24151
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 15470 24188 15476 24200
rect 15431 24160 15476 24188
rect 15470 24148 15476 24160
rect 15528 24148 15534 24200
rect 16574 24188 16580 24200
rect 16535 24160 16580 24188
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 18966 24188 18972 24200
rect 18927 24160 18972 24188
rect 18966 24148 18972 24160
rect 19024 24148 19030 24200
rect 19518 24188 19524 24200
rect 19479 24160 19524 24188
rect 19518 24148 19524 24160
rect 19576 24148 19582 24200
rect 19610 24148 19616 24200
rect 19668 24188 19674 24200
rect 19668 24160 19713 24188
rect 19668 24148 19674 24160
rect 21634 24148 21640 24200
rect 21692 24188 21698 24200
rect 23198 24188 23204 24200
rect 21692 24160 21737 24188
rect 23159 24160 23204 24188
rect 21692 24148 21698 24160
rect 23198 24148 23204 24160
rect 23256 24148 23262 24200
rect 21085 24123 21143 24129
rect 21085 24089 21097 24123
rect 21131 24120 21143 24123
rect 21266 24120 21272 24132
rect 21131 24092 21272 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 21266 24080 21272 24092
rect 21324 24120 21330 24132
rect 22465 24123 22523 24129
rect 22465 24120 22477 24123
rect 21324 24092 22477 24120
rect 21324 24080 21330 24092
rect 22465 24089 22477 24092
rect 22511 24089 22523 24123
rect 22646 24120 22652 24132
rect 22607 24092 22652 24120
rect 22465 24083 22523 24089
rect 22646 24080 22652 24092
rect 22704 24080 22710 24132
rect 12820 24024 13216 24052
rect 13909 24055 13967 24061
rect 13909 24021 13921 24055
rect 13955 24052 13967 24055
rect 13998 24052 14004 24064
rect 13955 24024 14004 24052
rect 13955 24021 13967 24024
rect 13909 24015 13967 24021
rect 13998 24012 14004 24024
rect 14056 24012 14062 24064
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 14645 24055 14703 24061
rect 14645 24052 14657 24055
rect 14516 24024 14657 24052
rect 14516 24012 14522 24024
rect 14645 24021 14657 24024
rect 14691 24021 14703 24055
rect 14645 24015 14703 24021
rect 14734 24012 14740 24064
rect 14792 24052 14798 24064
rect 15013 24055 15071 24061
rect 15013 24052 15025 24055
rect 14792 24024 15025 24052
rect 14792 24012 14798 24024
rect 15013 24021 15025 24024
rect 15059 24021 15071 24055
rect 15013 24015 15071 24021
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 16025 24055 16083 24061
rect 16025 24052 16037 24055
rect 15620 24024 16037 24052
rect 15620 24012 15626 24024
rect 16025 24021 16037 24024
rect 16071 24052 16083 24055
rect 16206 24052 16212 24064
rect 16071 24024 16212 24052
rect 16071 24021 16083 24024
rect 16025 24015 16083 24021
rect 16206 24012 16212 24024
rect 16264 24012 16270 24064
rect 16298 24012 16304 24064
rect 16356 24052 16362 24064
rect 16393 24055 16451 24061
rect 16393 24052 16405 24055
rect 16356 24024 16405 24052
rect 16356 24012 16362 24024
rect 16393 24021 16405 24024
rect 16439 24021 16451 24055
rect 17954 24052 17960 24064
rect 17915 24024 17960 24052
rect 16393 24015 16451 24021
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 19058 24052 19064 24064
rect 19019 24024 19064 24052
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 20438 24052 20444 24064
rect 20399 24024 20444 24052
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 22097 24055 22155 24061
rect 22097 24052 22109 24055
rect 21416 24024 22109 24052
rect 21416 24012 21422 24024
rect 22097 24021 22109 24024
rect 22143 24021 22155 24055
rect 23658 24052 23664 24064
rect 23619 24024 23664 24052
rect 22097 24015 22155 24021
rect 23658 24012 23664 24024
rect 23716 24012 23722 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 2498 23848 2504 23860
rect 2459 23820 2504 23848
rect 2498 23808 2504 23820
rect 2556 23808 2562 23860
rect 2958 23848 2964 23860
rect 2919 23820 2964 23848
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 3513 23851 3571 23857
rect 3513 23817 3525 23851
rect 3559 23848 3571 23851
rect 3970 23848 3976 23860
rect 3559 23820 3976 23848
rect 3559 23817 3571 23820
rect 3513 23811 3571 23817
rect 3970 23808 3976 23820
rect 4028 23808 4034 23860
rect 6273 23851 6331 23857
rect 6273 23817 6285 23851
rect 6319 23848 6331 23851
rect 6362 23848 6368 23860
rect 6319 23820 6368 23848
rect 6319 23817 6331 23820
rect 6273 23811 6331 23817
rect 3605 23783 3663 23789
rect 3605 23749 3617 23783
rect 3651 23780 3663 23783
rect 4522 23780 4528 23792
rect 3651 23752 4528 23780
rect 3651 23749 3663 23752
rect 3605 23743 3663 23749
rect 4522 23740 4528 23752
rect 4580 23740 4586 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23712 1731 23715
rect 3786 23712 3792 23724
rect 1719 23684 3792 23712
rect 1719 23681 1731 23684
rect 1673 23675 1731 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4154 23712 4160 23724
rect 4115 23684 4160 23712
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 5626 23712 5632 23724
rect 4755 23684 5632 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 5626 23672 5632 23684
rect 5684 23712 5690 23724
rect 5813 23715 5871 23721
rect 5813 23712 5825 23715
rect 5684 23684 5825 23712
rect 5684 23672 5690 23684
rect 5813 23681 5825 23684
rect 5859 23712 5871 23715
rect 6288 23712 6316 23811
rect 6362 23808 6368 23820
rect 6420 23808 6426 23860
rect 9030 23808 9036 23860
rect 9088 23848 9094 23860
rect 9125 23851 9183 23857
rect 9125 23848 9137 23851
rect 9088 23820 9137 23848
rect 9088 23808 9094 23820
rect 9125 23817 9137 23820
rect 9171 23848 9183 23851
rect 11330 23848 11336 23860
rect 9171 23820 11336 23848
rect 9171 23817 9183 23820
rect 9125 23811 9183 23817
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 13814 23808 13820 23860
rect 13872 23848 13878 23860
rect 14553 23851 14611 23857
rect 14553 23848 14565 23851
rect 13872 23820 14565 23848
rect 13872 23808 13878 23820
rect 14553 23817 14565 23820
rect 14599 23817 14611 23851
rect 14553 23811 14611 23817
rect 15013 23851 15071 23857
rect 15013 23817 15025 23851
rect 15059 23848 15071 23851
rect 15286 23848 15292 23860
rect 15059 23820 15292 23848
rect 15059 23817 15071 23820
rect 15013 23811 15071 23817
rect 8294 23740 8300 23792
rect 8352 23780 8358 23792
rect 9309 23783 9367 23789
rect 9309 23780 9321 23783
rect 8352 23752 9321 23780
rect 8352 23740 8358 23752
rect 9309 23749 9321 23752
rect 9355 23749 9367 23783
rect 9309 23743 9367 23749
rect 5859 23684 6316 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 8754 23672 8760 23724
rect 8812 23712 8818 23724
rect 9953 23715 10011 23721
rect 9953 23712 9965 23715
rect 8812 23684 9965 23712
rect 8812 23672 8818 23684
rect 9953 23681 9965 23684
rect 9999 23712 10011 23715
rect 10689 23715 10747 23721
rect 10689 23712 10701 23715
rect 9999 23684 10701 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 10689 23681 10701 23684
rect 10735 23681 10747 23715
rect 10689 23675 10747 23681
rect 10778 23672 10784 23724
rect 10836 23712 10842 23724
rect 11241 23715 11299 23721
rect 11241 23712 11253 23715
rect 10836 23684 11253 23712
rect 10836 23672 10842 23684
rect 11241 23681 11253 23684
rect 11287 23681 11299 23715
rect 11241 23675 11299 23681
rect 1397 23647 1455 23653
rect 1397 23613 1409 23647
rect 1443 23644 1455 23647
rect 2958 23644 2964 23656
rect 1443 23616 2964 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 2958 23604 2964 23616
rect 3016 23604 3022 23656
rect 3970 23604 3976 23656
rect 4028 23644 4034 23656
rect 4028 23616 4073 23644
rect 4028 23604 4034 23616
rect 6086 23604 6092 23656
rect 6144 23644 6150 23656
rect 6825 23647 6883 23653
rect 6825 23644 6837 23647
rect 6144 23616 6837 23644
rect 6144 23604 6150 23616
rect 6825 23613 6837 23616
rect 6871 23613 6883 23647
rect 6825 23607 6883 23613
rect 7650 23604 7656 23656
rect 7708 23644 7714 23656
rect 8018 23644 8024 23656
rect 7708 23616 8024 23644
rect 7708 23604 7714 23616
rect 8018 23604 8024 23616
rect 8076 23604 8082 23656
rect 9674 23604 9680 23656
rect 9732 23644 9738 23656
rect 9769 23647 9827 23653
rect 9769 23644 9781 23647
rect 9732 23616 9781 23644
rect 9732 23604 9738 23616
rect 9769 23613 9781 23616
rect 9815 23613 9827 23647
rect 11054 23644 11060 23656
rect 11015 23616 11060 23644
rect 9769 23607 9827 23613
rect 11054 23604 11060 23616
rect 11112 23604 11118 23656
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23644 12311 23647
rect 12299 23616 12388 23644
rect 12299 23613 12311 23616
rect 12253 23607 12311 23613
rect 3510 23536 3516 23588
rect 3568 23576 3574 23588
rect 5077 23579 5135 23585
rect 5077 23576 5089 23579
rect 3568 23548 5089 23576
rect 3568 23536 3574 23548
rect 5077 23545 5089 23548
rect 5123 23576 5135 23579
rect 5629 23579 5687 23585
rect 5629 23576 5641 23579
rect 5123 23548 5641 23576
rect 5123 23545 5135 23548
rect 5077 23539 5135 23545
rect 5629 23545 5641 23548
rect 5675 23576 5687 23579
rect 6362 23576 6368 23588
rect 5675 23548 6368 23576
rect 5675 23545 5687 23548
rect 5629 23539 5687 23545
rect 6362 23536 6368 23548
rect 6420 23536 6426 23588
rect 7070 23579 7128 23585
rect 7070 23576 7082 23579
rect 6840 23548 7082 23576
rect 6840 23520 6868 23548
rect 7070 23545 7082 23548
rect 7116 23545 7128 23579
rect 7070 23539 7128 23545
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8757 23579 8815 23585
rect 8757 23576 8769 23579
rect 7892 23548 8769 23576
rect 7892 23536 7898 23548
rect 8757 23545 8769 23548
rect 8803 23576 8815 23579
rect 9858 23576 9864 23588
rect 8803 23548 9864 23576
rect 8803 23545 8815 23548
rect 8757 23539 8815 23545
rect 9858 23536 9864 23548
rect 9916 23536 9922 23588
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12360 23576 12388 23616
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 14568 23644 14596 23811
rect 15286 23808 15292 23820
rect 15344 23808 15350 23860
rect 16666 23848 16672 23860
rect 16627 23820 16672 23848
rect 16666 23808 16672 23820
rect 16724 23808 16730 23860
rect 17034 23848 17040 23860
rect 16995 23820 17040 23848
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 17494 23848 17500 23860
rect 17455 23820 17500 23848
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 19521 23851 19579 23857
rect 19521 23817 19533 23851
rect 19567 23848 19579 23851
rect 19610 23848 19616 23860
rect 19567 23820 19616 23848
rect 19567 23817 19579 23820
rect 19521 23811 19579 23817
rect 19610 23808 19616 23820
rect 19668 23808 19674 23860
rect 21818 23808 21824 23860
rect 21876 23848 21882 23860
rect 21913 23851 21971 23857
rect 21913 23848 21925 23851
rect 21876 23820 21925 23848
rect 21876 23808 21882 23820
rect 21913 23817 21925 23820
rect 21959 23817 21971 23851
rect 22278 23848 22284 23860
rect 22239 23820 22284 23848
rect 21913 23811 21971 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 22649 23851 22707 23857
rect 22649 23817 22661 23851
rect 22695 23848 22707 23851
rect 22830 23848 22836 23860
rect 22695 23820 22836 23848
rect 22695 23817 22707 23820
rect 22649 23811 22707 23817
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 24118 23808 24124 23860
rect 24176 23848 24182 23860
rect 24581 23851 24639 23857
rect 24581 23848 24593 23851
rect 24176 23820 24593 23848
rect 24176 23808 24182 23820
rect 24581 23817 24593 23820
rect 24627 23817 24639 23851
rect 25130 23848 25136 23860
rect 25091 23820 25136 23848
rect 24581 23811 24639 23817
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 20714 23780 20720 23792
rect 20675 23752 20720 23780
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 20901 23783 20959 23789
rect 20901 23749 20913 23783
rect 20947 23780 20959 23783
rect 23658 23780 23664 23792
rect 20947 23752 23664 23780
rect 20947 23749 20959 23752
rect 20901 23743 20959 23749
rect 15381 23715 15439 23721
rect 15381 23681 15393 23715
rect 15427 23712 15439 23715
rect 16117 23715 16175 23721
rect 16117 23712 16129 23715
rect 15427 23684 16129 23712
rect 15427 23681 15439 23684
rect 15381 23675 15439 23681
rect 16117 23681 16129 23684
rect 16163 23712 16175 23715
rect 16666 23712 16672 23724
rect 16163 23684 16672 23712
rect 16163 23681 16175 23684
rect 16117 23675 16175 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 21453 23715 21511 23721
rect 21453 23712 21465 23715
rect 20487 23684 21465 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 21453 23681 21465 23684
rect 21499 23712 21511 23715
rect 22002 23712 22008 23724
rect 21499 23684 22008 23712
rect 21499 23681 21511 23684
rect 21453 23675 21511 23681
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 15933 23647 15991 23653
rect 15933 23644 15945 23647
rect 12492 23616 12537 23644
rect 14568 23616 15945 23644
rect 12492 23604 12498 23616
rect 15933 23613 15945 23616
rect 15979 23613 15991 23647
rect 15933 23607 15991 23613
rect 18046 23604 18052 23656
rect 18104 23644 18110 23656
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 18104 23616 18153 23644
rect 18104 23604 18110 23616
rect 18141 23613 18153 23616
rect 18187 23613 18199 23647
rect 18141 23607 18199 23613
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 21082 23644 21088 23656
rect 20956 23616 21088 23644
rect 20956 23604 20962 23616
rect 21082 23604 21088 23616
rect 21140 23604 21146 23656
rect 21266 23644 21272 23656
rect 21227 23616 21272 23644
rect 21266 23604 21272 23616
rect 21324 23604 21330 23656
rect 22462 23644 22468 23656
rect 22423 23616 22468 23644
rect 22462 23604 22468 23616
rect 22520 23644 22526 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22520 23616 23029 23644
rect 22520 23604 22526 23616
rect 23017 23613 23029 23616
rect 23063 23613 23075 23647
rect 23584 23644 23612 23752
rect 23658 23740 23664 23752
rect 23716 23740 23722 23792
rect 23661 23647 23719 23653
rect 23661 23644 23673 23647
rect 23584 23616 23673 23644
rect 23017 23607 23075 23613
rect 23661 23613 23673 23616
rect 23707 23613 23719 23647
rect 23661 23607 23719 23613
rect 24854 23604 24860 23656
rect 24912 23644 24918 23656
rect 24949 23647 25007 23653
rect 24949 23644 24961 23647
rect 24912 23616 24961 23644
rect 24912 23604 24918 23616
rect 24949 23613 24961 23616
rect 24995 23644 25007 23647
rect 25501 23647 25559 23653
rect 25501 23644 25513 23647
rect 24995 23616 25513 23644
rect 24995 23613 25007 23616
rect 24949 23607 25007 23613
rect 25501 23613 25513 23616
rect 25547 23613 25559 23647
rect 25501 23607 25559 23613
rect 12704 23579 12762 23585
rect 12704 23576 12716 23579
rect 11931 23548 12296 23576
rect 12360 23548 12716 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 1946 23468 1952 23520
rect 2004 23508 2010 23520
rect 2133 23511 2191 23517
rect 2133 23508 2145 23511
rect 2004 23480 2145 23508
rect 2004 23468 2010 23480
rect 2133 23477 2145 23480
rect 2179 23477 2191 23511
rect 2133 23471 2191 23477
rect 3694 23468 3700 23520
rect 3752 23508 3758 23520
rect 4065 23511 4123 23517
rect 4065 23508 4077 23511
rect 3752 23480 4077 23508
rect 3752 23468 3758 23480
rect 4065 23477 4077 23480
rect 4111 23477 4123 23511
rect 5166 23508 5172 23520
rect 5127 23480 5172 23508
rect 4065 23471 4123 23477
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5316 23480 5549 23508
rect 5316 23468 5322 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 5537 23471 5595 23477
rect 6641 23511 6699 23517
rect 6641 23477 6653 23511
rect 6687 23508 6699 23511
rect 6822 23508 6828 23520
rect 6687 23480 6828 23508
rect 6687 23477 6699 23480
rect 6641 23471 6699 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 7374 23468 7380 23520
rect 7432 23508 7438 23520
rect 8205 23511 8263 23517
rect 8205 23508 8217 23511
rect 7432 23480 8217 23508
rect 7432 23468 7438 23480
rect 8205 23477 8217 23480
rect 8251 23477 8263 23511
rect 8205 23471 8263 23477
rect 9030 23468 9036 23520
rect 9088 23508 9094 23520
rect 9677 23511 9735 23517
rect 9677 23508 9689 23511
rect 9088 23480 9689 23508
rect 9088 23468 9094 23480
rect 9677 23477 9689 23480
rect 9723 23477 9735 23511
rect 9677 23471 9735 23477
rect 9950 23468 9956 23520
rect 10008 23508 10014 23520
rect 10321 23511 10379 23517
rect 10321 23508 10333 23511
rect 10008 23480 10333 23508
rect 10008 23468 10014 23480
rect 10321 23477 10333 23480
rect 10367 23477 10379 23511
rect 12268 23508 12296 23548
rect 12704 23545 12716 23548
rect 12750 23576 12762 23579
rect 12802 23576 12808 23588
rect 12750 23548 12808 23576
rect 12750 23545 12762 23548
rect 12704 23539 12762 23545
rect 12802 23536 12808 23548
rect 12860 23536 12866 23588
rect 14182 23536 14188 23588
rect 14240 23576 14246 23588
rect 15654 23576 15660 23588
rect 14240 23548 15660 23576
rect 14240 23536 14246 23548
rect 15654 23536 15660 23548
rect 15712 23536 15718 23588
rect 15841 23579 15899 23585
rect 15841 23545 15853 23579
rect 15887 23576 15899 23579
rect 17034 23576 17040 23588
rect 15887 23548 17040 23576
rect 15887 23545 15899 23548
rect 15841 23539 15899 23545
rect 17034 23536 17040 23548
rect 17092 23536 17098 23588
rect 17865 23579 17923 23585
rect 17865 23545 17877 23579
rect 17911 23576 17923 23579
rect 17954 23576 17960 23588
rect 17911 23548 17960 23576
rect 17911 23545 17923 23548
rect 17865 23539 17923 23545
rect 17954 23536 17960 23548
rect 18012 23576 18018 23588
rect 18408 23579 18466 23585
rect 18408 23576 18420 23579
rect 18012 23548 18420 23576
rect 18012 23536 18018 23548
rect 18408 23545 18420 23548
rect 18454 23576 18466 23579
rect 18966 23576 18972 23588
rect 18454 23548 18972 23576
rect 18454 23545 18466 23548
rect 18408 23539 18466 23545
rect 18966 23536 18972 23548
rect 19024 23536 19030 23588
rect 21358 23576 21364 23588
rect 21319 23548 21364 23576
rect 21358 23536 21364 23548
rect 21416 23536 21422 23588
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 23937 23579 23995 23585
rect 23937 23576 23949 23579
rect 23532 23548 23949 23576
rect 23532 23536 23538 23548
rect 23937 23545 23949 23548
rect 23983 23545 23995 23579
rect 23937 23539 23995 23545
rect 12986 23508 12992 23520
rect 12268 23480 12992 23508
rect 10321 23471 10379 23477
rect 12986 23468 12992 23480
rect 13044 23468 13050 23520
rect 13814 23508 13820 23520
rect 13775 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 15470 23508 15476 23520
rect 15431 23480 15476 23508
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 23014 23468 23020 23520
rect 23072 23508 23078 23520
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 23072 23480 23397 23508
rect 23072 23468 23078 23480
rect 23385 23477 23397 23480
rect 23431 23508 23443 23511
rect 23842 23508 23848 23520
rect 23431 23480 23848 23508
rect 23431 23477 23443 23480
rect 23385 23471 23443 23477
rect 23842 23468 23848 23480
rect 23900 23468 23906 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 5626 23304 5632 23316
rect 5587 23276 5632 23304
rect 5626 23264 5632 23276
rect 5684 23264 5690 23316
rect 6086 23264 6092 23316
rect 6144 23304 6150 23316
rect 6181 23307 6239 23313
rect 6181 23304 6193 23307
rect 6144 23276 6193 23304
rect 6144 23264 6150 23276
rect 6181 23273 6193 23276
rect 6227 23304 6239 23307
rect 7282 23304 7288 23316
rect 6227 23276 7288 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 7282 23264 7288 23276
rect 7340 23304 7346 23316
rect 7745 23307 7803 23313
rect 7745 23304 7757 23307
rect 7340 23276 7757 23304
rect 7340 23264 7346 23276
rect 7745 23273 7757 23276
rect 7791 23273 7803 23307
rect 7745 23267 7803 23273
rect 9582 23264 9588 23316
rect 9640 23304 9646 23316
rect 10962 23304 10968 23316
rect 9640 23276 9812 23304
rect 9640 23264 9646 23276
rect 3694 23236 3700 23248
rect 3655 23208 3700 23236
rect 3694 23196 3700 23208
rect 3752 23196 3758 23248
rect 4246 23196 4252 23248
rect 4304 23236 4310 23248
rect 4494 23239 4552 23245
rect 4494 23236 4506 23239
rect 4304 23208 4506 23236
rect 4304 23196 4310 23208
rect 4494 23205 4506 23208
rect 4540 23205 4552 23239
rect 8570 23236 8576 23248
rect 8531 23208 8576 23236
rect 4494 23199 4552 23205
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 9784 23236 9812 23276
rect 10336 23276 10968 23304
rect 10336 23248 10364 23276
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 13354 23304 13360 23316
rect 13315 23276 13360 23304
rect 13354 23264 13360 23276
rect 13412 23264 13418 23316
rect 16666 23264 16672 23316
rect 16724 23304 16730 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 16724 23276 16773 23304
rect 16724 23264 16730 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 16761 23267 16819 23273
rect 19153 23307 19211 23313
rect 19153 23273 19165 23307
rect 19199 23304 19211 23307
rect 19518 23304 19524 23316
rect 19199 23276 19524 23304
rect 19199 23273 19211 23276
rect 19153 23267 19211 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 22094 23264 22100 23316
rect 22152 23304 22158 23316
rect 22370 23304 22376 23316
rect 22152 23276 22376 23304
rect 22152 23264 22158 23276
rect 22370 23264 22376 23276
rect 22428 23304 22434 23316
rect 22557 23307 22615 23313
rect 22557 23304 22569 23307
rect 22428 23276 22569 23304
rect 22428 23264 22434 23276
rect 22557 23273 22569 23276
rect 22603 23273 22615 23307
rect 23658 23304 23664 23316
rect 23619 23276 23664 23304
rect 22557 23267 22615 23273
rect 23658 23264 23664 23276
rect 23716 23264 23722 23316
rect 25409 23307 25467 23313
rect 25409 23273 25421 23307
rect 25455 23304 25467 23307
rect 25682 23304 25688 23316
rect 25455 23276 25688 23304
rect 25455 23273 25467 23276
rect 25409 23267 25467 23273
rect 25682 23264 25688 23276
rect 25740 23264 25746 23316
rect 10226 23236 10232 23248
rect 9784 23208 10232 23236
rect 10226 23196 10232 23208
rect 10284 23196 10290 23248
rect 10318 23196 10324 23248
rect 10376 23196 10382 23248
rect 11692 23239 11750 23245
rect 11692 23236 11704 23239
rect 10520 23208 11704 23236
rect 1489 23171 1547 23177
rect 1489 23137 1501 23171
rect 1535 23168 1547 23171
rect 2590 23168 2596 23180
rect 1535 23140 2596 23168
rect 1535 23137 1547 23140
rect 1489 23131 1547 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 2777 23171 2835 23177
rect 2777 23137 2789 23171
rect 2823 23168 2835 23171
rect 3326 23168 3332 23180
rect 2823 23140 3332 23168
rect 2823 23137 2835 23140
rect 2777 23131 2835 23137
rect 3326 23128 3332 23140
rect 3384 23128 3390 23180
rect 6546 23128 6552 23180
rect 6604 23168 6610 23180
rect 7101 23171 7159 23177
rect 7101 23168 7113 23171
rect 6604 23140 7113 23168
rect 6604 23128 6610 23140
rect 7101 23137 7113 23140
rect 7147 23137 7159 23171
rect 7101 23131 7159 23137
rect 8297 23171 8355 23177
rect 8297 23137 8309 23171
rect 8343 23168 8355 23171
rect 8662 23168 8668 23180
rect 8343 23140 8668 23168
rect 8343 23137 8355 23140
rect 8297 23131 8355 23137
rect 8662 23128 8668 23140
rect 8720 23128 8726 23180
rect 1762 23100 1768 23112
rect 1723 23072 1768 23100
rect 1762 23060 1768 23072
rect 1820 23060 1826 23112
rect 2958 23060 2964 23112
rect 3016 23100 3022 23112
rect 4249 23103 4307 23109
rect 4249 23100 4261 23103
rect 3016 23072 4261 23100
rect 3016 23060 3022 23072
rect 4249 23069 4261 23072
rect 4295 23069 4307 23103
rect 4249 23063 4307 23069
rect 6638 23060 6644 23112
rect 6696 23100 6702 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 6696 23072 7205 23100
rect 6696 23060 6702 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7374 23100 7380 23112
rect 7335 23072 7380 23100
rect 7193 23063 7251 23069
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 8202 23100 8208 23112
rect 8163 23072 8208 23100
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 9858 23060 9864 23112
rect 9916 23100 9922 23112
rect 10318 23100 10324 23112
rect 9916 23072 10324 23100
rect 9916 23060 9922 23072
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 10520 23109 10548 23208
rect 11692 23205 11704 23208
rect 11738 23236 11750 23239
rect 11882 23236 11888 23248
rect 11738 23208 11888 23236
rect 11738 23205 11750 23208
rect 11692 23199 11750 23205
rect 11882 23196 11888 23208
rect 11940 23236 11946 23248
rect 12250 23236 12256 23248
rect 11940 23208 12256 23236
rect 11940 23196 11946 23208
rect 12250 23196 12256 23208
rect 12308 23196 12314 23248
rect 12710 23196 12716 23248
rect 12768 23236 12774 23248
rect 14185 23239 14243 23245
rect 14185 23236 14197 23239
rect 12768 23208 14197 23236
rect 12768 23196 12774 23208
rect 14185 23205 14197 23208
rect 14231 23205 14243 23239
rect 16574 23236 16580 23248
rect 14185 23199 14243 23205
rect 15396 23208 16580 23236
rect 13906 23168 13912 23180
rect 13867 23140 13912 23168
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 15396 23177 15424 23208
rect 16574 23196 16580 23208
rect 16632 23236 16638 23248
rect 17313 23239 17371 23245
rect 17313 23236 17325 23239
rect 16632 23208 17325 23236
rect 16632 23196 16638 23208
rect 17313 23205 17325 23208
rect 17359 23205 17371 23239
rect 17313 23199 17371 23205
rect 20717 23239 20775 23245
rect 20717 23205 20729 23239
rect 20763 23236 20775 23239
rect 21444 23239 21502 23245
rect 21444 23236 21456 23239
rect 20763 23208 21456 23236
rect 20763 23205 20775 23208
rect 20717 23199 20775 23205
rect 21444 23205 21456 23208
rect 21490 23236 21502 23239
rect 21634 23236 21640 23248
rect 21490 23208 21640 23236
rect 21490 23205 21502 23208
rect 21444 23199 21502 23205
rect 15654 23177 15660 23180
rect 14737 23171 14795 23177
rect 14737 23137 14749 23171
rect 14783 23168 14795 23171
rect 15105 23171 15163 23177
rect 15105 23168 15117 23171
rect 14783 23140 15117 23168
rect 14783 23137 14795 23140
rect 14737 23131 14795 23137
rect 15105 23137 15117 23140
rect 15151 23168 15163 23171
rect 15381 23171 15439 23177
rect 15381 23168 15393 23171
rect 15151 23140 15393 23168
rect 15151 23137 15163 23140
rect 15105 23131 15163 23137
rect 15381 23137 15393 23140
rect 15427 23137 15439 23171
rect 15648 23168 15660 23177
rect 15567 23140 15660 23168
rect 15381 23131 15439 23137
rect 15648 23131 15660 23140
rect 15712 23168 15718 23180
rect 16850 23168 16856 23180
rect 15712 23140 16856 23168
rect 15654 23128 15660 23131
rect 15712 23128 15718 23140
rect 16850 23128 16856 23140
rect 16908 23128 16914 23180
rect 17954 23168 17960 23180
rect 17867 23140 17960 23168
rect 17954 23128 17960 23140
rect 18012 23168 18018 23180
rect 19058 23168 19064 23180
rect 18012 23140 19064 23168
rect 18012 23128 18018 23140
rect 19058 23128 19064 23140
rect 19116 23128 19122 23180
rect 19610 23168 19616 23180
rect 19571 23140 19616 23168
rect 19610 23128 19616 23140
rect 19668 23128 19674 23180
rect 20254 23168 20260 23180
rect 19812 23140 20260 23168
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23069 10563 23103
rect 11425 23103 11483 23109
rect 11425 23100 11437 23103
rect 10505 23063 10563 23069
rect 11256 23072 11437 23100
rect 6730 23032 6736 23044
rect 6691 23004 6736 23032
rect 6730 22992 6736 23004
rect 6788 22992 6794 23044
rect 2317 22967 2375 22973
rect 2317 22933 2329 22967
rect 2363 22964 2375 22967
rect 2406 22964 2412 22976
rect 2363 22936 2412 22964
rect 2363 22933 2375 22936
rect 2317 22927 2375 22933
rect 2406 22924 2412 22936
rect 2464 22924 2470 22976
rect 2866 22924 2872 22976
rect 2924 22964 2930 22976
rect 2961 22967 3019 22973
rect 2961 22964 2973 22967
rect 2924 22936 2973 22964
rect 2924 22924 2930 22936
rect 2961 22933 2973 22936
rect 3007 22933 3019 22967
rect 6546 22964 6552 22976
rect 6507 22936 6552 22964
rect 2961 22927 3019 22933
rect 6546 22924 6552 22936
rect 6604 22924 6610 22976
rect 9398 22964 9404 22976
rect 9359 22936 9404 22964
rect 9398 22924 9404 22936
rect 9456 22924 9462 22976
rect 9858 22964 9864 22976
rect 9819 22936 9864 22964
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 10962 22964 10968 22976
rect 10923 22936 10968 22964
rect 10962 22924 10968 22936
rect 11020 22924 11026 22976
rect 11146 22924 11152 22976
rect 11204 22964 11210 22976
rect 11256 22973 11284 23072
rect 11425 23069 11437 23072
rect 11471 23069 11483 23103
rect 18138 23100 18144 23112
rect 18099 23072 18144 23100
rect 11425 23063 11483 23069
rect 18138 23060 18144 23072
rect 18196 23060 18202 23112
rect 19702 23100 19708 23112
rect 19663 23072 19708 23100
rect 19702 23060 19708 23072
rect 19760 23060 19766 23112
rect 19812 23109 19840 23140
rect 20254 23128 20260 23140
rect 20312 23168 20318 23180
rect 20732 23168 20760 23199
rect 21634 23196 21640 23208
rect 21692 23196 21698 23248
rect 21910 23196 21916 23248
rect 21968 23236 21974 23248
rect 21968 23208 24256 23236
rect 21968 23196 21974 23208
rect 20312 23140 20760 23168
rect 20312 23128 20318 23140
rect 23106 23128 23112 23180
rect 23164 23168 23170 23180
rect 24029 23171 24087 23177
rect 24029 23168 24041 23171
rect 23164 23140 24041 23168
rect 23164 23128 23170 23140
rect 24029 23137 24041 23140
rect 24075 23137 24087 23171
rect 24029 23131 24087 23137
rect 24228 23112 24256 23208
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25774 23168 25780 23180
rect 25271 23140 25780 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23069 19855 23103
rect 19797 23063 19855 23069
rect 19886 23060 19892 23112
rect 19944 23100 19950 23112
rect 20898 23100 20904 23112
rect 19944 23072 20904 23100
rect 19944 23060 19950 23072
rect 20898 23060 20904 23072
rect 20956 23100 20962 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 20956 23072 21189 23100
rect 20956 23060 20962 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 23569 23103 23627 23109
rect 23569 23069 23581 23103
rect 23615 23100 23627 23103
rect 23658 23100 23664 23112
rect 23615 23072 23664 23100
rect 23615 23069 23627 23072
rect 23569 23063 23627 23069
rect 23658 23060 23664 23072
rect 23716 23060 23722 23112
rect 24118 23100 24124 23112
rect 24079 23072 24124 23100
rect 24118 23060 24124 23072
rect 24176 23060 24182 23112
rect 24210 23060 24216 23112
rect 24268 23100 24274 23112
rect 24268 23072 24361 23100
rect 24268 23060 24274 23072
rect 13725 23035 13783 23041
rect 13725 23032 13737 23035
rect 12452 23004 13737 23032
rect 12452 22976 12480 23004
rect 13725 23001 13737 23004
rect 13771 23001 13783 23035
rect 13725 22995 13783 23001
rect 19150 22992 19156 23044
rect 19208 23032 19214 23044
rect 19426 23032 19432 23044
rect 19208 23004 19432 23032
rect 19208 22992 19214 23004
rect 19426 22992 19432 23004
rect 19484 23032 19490 23044
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 19484 23004 20269 23032
rect 19484 22992 19490 23004
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 11204 22936 11253 22964
rect 11204 22924 11210 22936
rect 11241 22933 11253 22936
rect 11287 22964 11299 22967
rect 12434 22964 12440 22976
rect 11287 22936 12440 22964
rect 11287 22933 11299 22936
rect 11241 22927 11299 22933
rect 12434 22924 12440 22936
rect 12492 22924 12498 22976
rect 12802 22964 12808 22976
rect 12763 22936 12808 22964
rect 12802 22924 12808 22936
rect 12860 22924 12866 22976
rect 17865 22967 17923 22973
rect 17865 22933 17877 22967
rect 17911 22964 17923 22967
rect 18046 22964 18052 22976
rect 17911 22936 18052 22964
rect 17911 22933 17923 22936
rect 17865 22927 17923 22933
rect 18046 22924 18052 22936
rect 18104 22924 18110 22976
rect 18785 22967 18843 22973
rect 18785 22933 18797 22967
rect 18831 22964 18843 22967
rect 18966 22964 18972 22976
rect 18831 22936 18972 22964
rect 18831 22933 18843 22936
rect 18785 22927 18843 22933
rect 18966 22924 18972 22936
rect 19024 22924 19030 22976
rect 19242 22964 19248 22976
rect 19203 22936 19248 22964
rect 19242 22924 19248 22936
rect 19300 22924 19306 22976
rect 22462 22924 22468 22976
rect 22520 22964 22526 22976
rect 23109 22967 23167 22973
rect 23109 22964 23121 22967
rect 22520 22936 23121 22964
rect 22520 22924 22526 22936
rect 23109 22933 23121 22936
rect 23155 22964 23167 22967
rect 23198 22964 23204 22976
rect 23155 22936 23204 22964
rect 23155 22933 23167 22936
rect 23109 22927 23167 22933
rect 23198 22924 23204 22936
rect 23256 22924 23262 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 566 22720 572 22772
rect 624 22760 630 22772
rect 5629 22763 5687 22769
rect 5629 22760 5641 22763
rect 624 22732 5641 22760
rect 624 22720 630 22732
rect 5629 22729 5641 22732
rect 5675 22729 5687 22763
rect 5629 22723 5687 22729
rect 7101 22763 7159 22769
rect 7101 22729 7113 22763
rect 7147 22760 7159 22763
rect 7374 22760 7380 22772
rect 7147 22732 7380 22760
rect 7147 22729 7159 22732
rect 7101 22723 7159 22729
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 9674 22720 9680 22772
rect 9732 22760 9738 22772
rect 10042 22760 10048 22772
rect 9732 22732 10048 22760
rect 9732 22720 9738 22732
rect 10042 22720 10048 22732
rect 10100 22720 10106 22772
rect 10318 22760 10324 22772
rect 10279 22732 10324 22760
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 11882 22760 11888 22772
rect 11843 22732 11888 22760
rect 11882 22720 11888 22732
rect 11940 22720 11946 22772
rect 15013 22763 15071 22769
rect 15013 22729 15025 22763
rect 15059 22760 15071 22763
rect 15654 22760 15660 22772
rect 15059 22732 15660 22760
rect 15059 22729 15071 22732
rect 15013 22723 15071 22729
rect 2958 22624 2964 22636
rect 2919 22596 2964 22624
rect 2958 22584 2964 22596
rect 3016 22584 3022 22636
rect 7392 22624 7420 22720
rect 9953 22695 10011 22701
rect 9953 22661 9965 22695
rect 9999 22692 10011 22695
rect 10226 22692 10232 22704
rect 9999 22664 10232 22692
rect 9999 22661 10011 22664
rect 9953 22655 10011 22661
rect 10226 22652 10232 22664
rect 10284 22652 10290 22704
rect 9585 22627 9643 22633
rect 7392 22596 7512 22624
rect 1489 22559 1547 22565
rect 1489 22525 1501 22559
rect 1535 22556 1547 22559
rect 2406 22556 2412 22568
rect 1535 22528 2412 22556
rect 1535 22525 1547 22528
rect 1489 22519 1547 22525
rect 2406 22516 2412 22528
rect 2464 22516 2470 22568
rect 2774 22516 2780 22568
rect 2832 22516 2838 22568
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 5445 22559 5503 22565
rect 5445 22556 5457 22559
rect 5408 22528 5457 22556
rect 5408 22516 5414 22528
rect 5445 22525 5457 22528
rect 5491 22556 5503 22559
rect 5997 22559 6055 22565
rect 5997 22556 6009 22559
rect 5491 22528 6009 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 5997 22525 6009 22528
rect 6043 22525 6055 22559
rect 5997 22519 6055 22525
rect 7282 22516 7288 22568
rect 7340 22556 7346 22568
rect 7377 22559 7435 22565
rect 7377 22556 7389 22559
rect 7340 22528 7389 22556
rect 7340 22516 7346 22528
rect 7377 22525 7389 22528
rect 7423 22525 7435 22559
rect 7484 22556 7512 22596
rect 9585 22593 9597 22627
rect 9631 22624 9643 22627
rect 11422 22624 11428 22636
rect 9631 22596 11428 22624
rect 9631 22593 9643 22596
rect 9585 22587 9643 22593
rect 11422 22584 11428 22596
rect 11480 22624 11486 22636
rect 11900 22624 11928 22720
rect 13998 22652 14004 22704
rect 14056 22692 14062 22704
rect 15028 22692 15056 22723
rect 15654 22720 15660 22732
rect 15712 22720 15718 22772
rect 18233 22763 18291 22769
rect 18233 22729 18245 22763
rect 18279 22760 18291 22763
rect 19150 22760 19156 22772
rect 18279 22732 19156 22760
rect 18279 22729 18291 22732
rect 18233 22723 18291 22729
rect 19150 22720 19156 22732
rect 19208 22720 19214 22772
rect 19337 22763 19395 22769
rect 19337 22729 19349 22763
rect 19383 22760 19395 22763
rect 19610 22760 19616 22772
rect 19383 22732 19616 22760
rect 19383 22729 19395 22732
rect 19337 22723 19395 22729
rect 19610 22720 19616 22732
rect 19668 22720 19674 22772
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 21634 22760 21640 22772
rect 21223 22732 21640 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21634 22720 21640 22732
rect 21692 22760 21698 22772
rect 21729 22763 21787 22769
rect 21729 22760 21741 22763
rect 21692 22732 21741 22760
rect 21692 22720 21698 22732
rect 21729 22729 21741 22732
rect 21775 22729 21787 22763
rect 21729 22723 21787 22729
rect 22646 22720 22652 22772
rect 22704 22760 22710 22772
rect 23106 22760 23112 22772
rect 22704 22732 23112 22760
rect 22704 22720 22710 22732
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 25409 22763 25467 22769
rect 25409 22729 25421 22763
rect 25455 22760 25467 22763
rect 25590 22760 25596 22772
rect 25455 22732 25596 22760
rect 25455 22729 25467 22732
rect 25409 22723 25467 22729
rect 25590 22720 25596 22732
rect 25648 22720 25654 22772
rect 16850 22692 16856 22704
rect 14056 22664 15056 22692
rect 16763 22664 16856 22692
rect 14056 22652 14062 22664
rect 16850 22652 16856 22664
rect 16908 22692 16914 22704
rect 18414 22692 18420 22704
rect 16908 22664 18420 22692
rect 16908 22652 16914 22664
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 12434 22624 12440 22636
rect 11480 22596 11928 22624
rect 12395 22596 12440 22624
rect 11480 22584 11486 22596
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 17586 22584 17592 22636
rect 17644 22624 17650 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17644 22596 17877 22624
rect 17644 22584 17650 22596
rect 17865 22593 17877 22596
rect 17911 22624 17923 22627
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 17911 22596 18705 22624
rect 17911 22593 17923 22596
rect 17865 22587 17923 22593
rect 18693 22593 18705 22596
rect 18739 22624 18751 22627
rect 18782 22624 18788 22636
rect 18739 22596 18788 22624
rect 18739 22593 18751 22596
rect 18693 22587 18751 22593
rect 18782 22584 18788 22596
rect 18840 22584 18846 22636
rect 18877 22627 18935 22633
rect 18877 22593 18889 22627
rect 18923 22624 18935 22627
rect 18966 22624 18972 22636
rect 18923 22596 18972 22624
rect 18923 22593 18935 22596
rect 18877 22587 18935 22593
rect 18966 22584 18972 22596
rect 19024 22584 19030 22636
rect 19518 22584 19524 22636
rect 19576 22624 19582 22636
rect 24305 22627 24363 22633
rect 19576 22596 19932 22624
rect 19576 22584 19582 22596
rect 7633 22559 7691 22565
rect 7633 22556 7645 22559
rect 7484 22528 7645 22556
rect 7377 22519 7435 22525
rect 7633 22525 7645 22528
rect 7679 22525 7691 22559
rect 10594 22556 10600 22568
rect 10555 22528 10600 22556
rect 7633 22519 7691 22525
rect 10594 22516 10600 22528
rect 10652 22516 10658 22568
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11149 22559 11207 22565
rect 11149 22556 11161 22559
rect 11020 22528 11161 22556
rect 11020 22516 11026 22528
rect 11149 22525 11161 22528
rect 11195 22556 11207 22559
rect 12158 22556 12164 22568
rect 11195 22528 12164 22556
rect 11195 22525 11207 22528
rect 11149 22519 11207 22525
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12704 22559 12762 22565
rect 12704 22556 12716 22559
rect 12636 22528 12716 22556
rect 1762 22488 1768 22500
rect 1723 22460 1768 22488
rect 1762 22448 1768 22460
rect 1820 22448 1826 22500
rect 2501 22491 2559 22497
rect 2501 22457 2513 22491
rect 2547 22488 2559 22491
rect 2792 22488 2820 22516
rect 3206 22491 3264 22497
rect 3206 22488 3218 22491
rect 2547 22460 3218 22488
rect 2547 22457 2559 22460
rect 2501 22451 2559 22457
rect 3206 22457 3218 22460
rect 3252 22457 3264 22491
rect 10612 22488 10640 22516
rect 11238 22488 11244 22500
rect 10612 22460 11244 22488
rect 3206 22451 3264 22457
rect 11238 22448 11244 22460
rect 11296 22448 11302 22500
rect 12250 22488 12256 22500
rect 12163 22460 12256 22488
rect 12250 22448 12256 22460
rect 12308 22488 12314 22500
rect 12636 22488 12664 22528
rect 12704 22525 12716 22528
rect 12750 22556 12762 22559
rect 13722 22556 13728 22568
rect 12750 22528 13728 22556
rect 12750 22525 12762 22528
rect 12704 22519 12762 22525
rect 13004 22500 13032 22528
rect 13722 22516 13728 22528
rect 13780 22516 13786 22568
rect 15102 22516 15108 22568
rect 15160 22556 15166 22568
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 15160 22528 15485 22556
rect 15160 22516 15166 22528
rect 15473 22525 15485 22528
rect 15519 22556 15531 22559
rect 16574 22556 16580 22568
rect 15519 22528 16580 22556
rect 15519 22525 15531 22528
rect 15473 22519 15531 22525
rect 16574 22516 16580 22528
rect 16632 22516 16638 22568
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 19484 22528 19625 22556
rect 19484 22516 19490 22528
rect 19613 22525 19625 22528
rect 19659 22525 19671 22559
rect 19794 22556 19800 22568
rect 19755 22528 19800 22556
rect 19613 22519 19671 22525
rect 19794 22516 19800 22528
rect 19852 22516 19858 22568
rect 19904 22556 19932 22596
rect 24305 22593 24317 22627
rect 24351 22624 24363 22627
rect 24351 22596 25176 22624
rect 24351 22593 24363 22596
rect 24305 22587 24363 22593
rect 20070 22565 20076 22568
rect 20053 22559 20076 22565
rect 20053 22556 20065 22559
rect 19904 22528 20065 22556
rect 20053 22525 20065 22528
rect 20128 22556 20134 22568
rect 22281 22559 22339 22565
rect 22281 22556 22293 22559
rect 20128 22528 20201 22556
rect 22112 22528 22293 22556
rect 20053 22519 20076 22525
rect 20070 22516 20076 22519
rect 20128 22516 20134 22528
rect 12308 22460 12664 22488
rect 12308 22448 12314 22460
rect 12986 22448 12992 22500
rect 13044 22448 13050 22500
rect 15746 22497 15752 22500
rect 15381 22491 15439 22497
rect 15381 22457 15393 22491
rect 15427 22488 15439 22491
rect 15740 22488 15752 22497
rect 15427 22460 15752 22488
rect 15427 22457 15439 22460
rect 15381 22451 15439 22457
rect 15740 22451 15752 22460
rect 15746 22448 15752 22451
rect 15804 22448 15810 22500
rect 17402 22448 17408 22500
rect 17460 22488 17466 22500
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 17460 22460 17509 22488
rect 17460 22448 17466 22460
rect 17497 22457 17509 22460
rect 17543 22488 17555 22491
rect 18601 22491 18659 22497
rect 18601 22488 18613 22491
rect 17543 22460 18613 22488
rect 17543 22457 17555 22460
rect 17497 22451 17555 22457
rect 18601 22457 18613 22460
rect 18647 22457 18659 22491
rect 18601 22451 18659 22457
rect 22112 22432 22140 22528
rect 22281 22525 22293 22528
rect 22327 22525 22339 22559
rect 23474 22556 23480 22568
rect 23435 22528 23480 22556
rect 22281 22519 22339 22525
rect 23474 22516 23480 22528
rect 23532 22556 23538 22568
rect 24121 22559 24179 22565
rect 24121 22556 24133 22559
rect 23532 22528 24133 22556
rect 23532 22516 23538 22528
rect 24121 22525 24133 22528
rect 24167 22556 24179 22559
rect 24854 22556 24860 22568
rect 24167 22528 24860 22556
rect 24167 22525 24179 22528
rect 24121 22519 24179 22525
rect 24854 22516 24860 22528
rect 24912 22516 24918 22568
rect 22554 22488 22560 22500
rect 22515 22460 22560 22488
rect 22554 22448 22560 22460
rect 22612 22448 22618 22500
rect 23566 22448 23572 22500
rect 23624 22488 23630 22500
rect 24029 22491 24087 22497
rect 24029 22488 24041 22491
rect 23624 22460 24041 22488
rect 23624 22448 23630 22460
rect 24029 22457 24041 22460
rect 24075 22488 24087 22491
rect 24673 22491 24731 22497
rect 24673 22488 24685 22491
rect 24075 22460 24685 22488
rect 24075 22457 24087 22460
rect 24029 22451 24087 22457
rect 24673 22457 24685 22460
rect 24719 22457 24731 22491
rect 24673 22451 24731 22457
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 2958 22420 2964 22432
rect 2915 22392 2964 22420
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 4246 22380 4252 22432
rect 4304 22420 4310 22432
rect 4341 22423 4399 22429
rect 4341 22420 4353 22423
rect 4304 22392 4353 22420
rect 4304 22380 4310 22392
rect 4341 22389 4353 22392
rect 4387 22420 4399 22423
rect 4893 22423 4951 22429
rect 4893 22420 4905 22423
rect 4387 22392 4905 22420
rect 4387 22389 4399 22392
rect 4341 22383 4399 22389
rect 4893 22389 4905 22392
rect 4939 22389 4951 22423
rect 4893 22383 4951 22389
rect 5353 22423 5411 22429
rect 5353 22389 5365 22423
rect 5399 22420 5411 22423
rect 5534 22420 5540 22432
rect 5399 22392 5540 22420
rect 5399 22389 5411 22392
rect 5353 22383 5411 22389
rect 5534 22380 5540 22392
rect 5592 22380 5598 22432
rect 6638 22420 6644 22432
rect 6599 22392 6644 22420
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 7466 22380 7472 22432
rect 7524 22420 7530 22432
rect 7834 22420 7840 22432
rect 7524 22392 7840 22420
rect 7524 22380 7530 22392
rect 7834 22380 7840 22392
rect 7892 22380 7898 22432
rect 8754 22420 8760 22432
rect 8715 22392 8760 22420
rect 8754 22380 8760 22392
rect 8812 22420 8818 22432
rect 9122 22420 9128 22432
rect 8812 22392 9128 22420
rect 8812 22380 8818 22392
rect 9122 22380 9128 22392
rect 9180 22380 9186 22432
rect 10778 22420 10784 22432
rect 10739 22392 10784 22420
rect 10778 22380 10784 22392
rect 10836 22380 10842 22432
rect 13817 22423 13875 22429
rect 13817 22389 13829 22423
rect 13863 22420 13875 22423
rect 13906 22420 13912 22432
rect 13863 22392 13912 22420
rect 13863 22389 13875 22392
rect 13817 22383 13875 22389
rect 13906 22380 13912 22392
rect 13964 22380 13970 22432
rect 13998 22380 14004 22432
rect 14056 22420 14062 22432
rect 14274 22420 14280 22432
rect 14056 22392 14280 22420
rect 14056 22380 14062 22392
rect 14274 22380 14280 22392
rect 14332 22420 14338 22432
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 14332 22392 14381 22420
rect 14332 22380 14338 22392
rect 14369 22389 14381 22392
rect 14415 22389 14427 22423
rect 14369 22383 14427 22389
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 22152 22392 22197 22420
rect 22152 22380 22158 22392
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 25148 22429 25176 22596
rect 25225 22559 25283 22565
rect 25225 22525 25237 22559
rect 25271 22556 25283 22559
rect 25590 22556 25596 22568
rect 25271 22528 25596 22556
rect 25271 22525 25283 22528
rect 25225 22519 25283 22525
rect 25590 22516 25596 22528
rect 25648 22516 25654 22568
rect 23661 22423 23719 22429
rect 23661 22420 23673 22423
rect 23440 22392 23673 22420
rect 23440 22380 23446 22392
rect 23661 22389 23673 22392
rect 23707 22389 23719 22423
rect 23661 22383 23719 22389
rect 25133 22423 25191 22429
rect 25133 22389 25145 22423
rect 25179 22420 25191 22423
rect 25222 22420 25228 22432
rect 25179 22392 25228 22420
rect 25179 22389 25191 22392
rect 25133 22383 25191 22389
rect 25222 22380 25228 22392
rect 25280 22380 25286 22432
rect 25774 22420 25780 22432
rect 25735 22392 25780 22420
rect 25774 22380 25780 22392
rect 25832 22380 25838 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 2406 22216 2412 22228
rect 2367 22188 2412 22216
rect 2406 22176 2412 22188
rect 2464 22176 2470 22228
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 3142 22216 3148 22228
rect 2823 22188 3148 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 3142 22176 3148 22188
rect 3200 22216 3206 22228
rect 3421 22219 3479 22225
rect 3421 22216 3433 22219
rect 3200 22188 3433 22216
rect 3200 22176 3206 22188
rect 3421 22185 3433 22188
rect 3467 22185 3479 22219
rect 4522 22216 4528 22228
rect 4483 22188 4528 22216
rect 3421 22179 3479 22185
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 5997 22219 6055 22225
rect 5997 22185 6009 22219
rect 6043 22216 6055 22219
rect 6546 22216 6552 22228
rect 6043 22188 6552 22216
rect 6043 22185 6055 22188
rect 5997 22179 6055 22185
rect 6546 22176 6552 22188
rect 6604 22176 6610 22228
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7561 22219 7619 22225
rect 7561 22216 7573 22219
rect 6696 22188 7573 22216
rect 6696 22176 6702 22188
rect 7561 22185 7573 22188
rect 7607 22185 7619 22219
rect 7561 22179 7619 22185
rect 7929 22219 7987 22225
rect 7929 22185 7941 22219
rect 7975 22216 7987 22219
rect 8202 22216 8208 22228
rect 7975 22188 8208 22216
rect 7975 22185 7987 22188
rect 7929 22179 7987 22185
rect 1394 22148 1400 22160
rect 1355 22120 1400 22148
rect 1394 22108 1400 22120
rect 1452 22108 1458 22160
rect 2869 22151 2927 22157
rect 2869 22148 2881 22151
rect 2792 22120 2881 22148
rect 1949 22083 2007 22089
rect 1949 22049 1961 22083
rect 1995 22080 2007 22083
rect 2038 22080 2044 22092
rect 1995 22052 2044 22080
rect 1995 22049 2007 22052
rect 1949 22043 2007 22049
rect 2038 22040 2044 22052
rect 2096 22040 2102 22092
rect 2317 21947 2375 21953
rect 2317 21913 2329 21947
rect 2363 21944 2375 21947
rect 2792 21944 2820 22120
rect 2869 22117 2881 22120
rect 2915 22117 2927 22151
rect 2869 22111 2927 22117
rect 4433 22151 4491 22157
rect 4433 22117 4445 22151
rect 4479 22148 4491 22151
rect 4614 22148 4620 22160
rect 4479 22120 4620 22148
rect 4479 22117 4491 22120
rect 4433 22111 4491 22117
rect 4614 22108 4620 22120
rect 4672 22108 4678 22160
rect 7374 22148 7380 22160
rect 7335 22120 7380 22148
rect 7374 22108 7380 22120
rect 7432 22108 7438 22160
rect 4246 22080 4252 22092
rect 3068 22052 4252 22080
rect 3068 22024 3096 22052
rect 4246 22040 4252 22052
rect 4304 22040 4310 22092
rect 6086 22040 6092 22092
rect 6144 22080 6150 22092
rect 6365 22083 6423 22089
rect 6365 22080 6377 22083
rect 6144 22052 6377 22080
rect 6144 22040 6150 22052
rect 6365 22049 6377 22052
rect 6411 22049 6423 22083
rect 6365 22043 6423 22049
rect 7101 22083 7159 22089
rect 7101 22049 7113 22083
rect 7147 22080 7159 22083
rect 7944 22080 7972 22179
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10413 22219 10471 22225
rect 10413 22216 10425 22219
rect 10192 22188 10425 22216
rect 10192 22176 10198 22188
rect 10413 22185 10425 22188
rect 10459 22185 10471 22219
rect 10413 22179 10471 22185
rect 11149 22219 11207 22225
rect 11149 22185 11161 22219
rect 11195 22216 11207 22219
rect 11422 22216 11428 22228
rect 11195 22188 11428 22216
rect 11195 22185 11207 22188
rect 11149 22179 11207 22185
rect 11422 22176 11428 22188
rect 11480 22176 11486 22228
rect 12342 22216 12348 22228
rect 12303 22188 12348 22216
rect 12342 22176 12348 22188
rect 12400 22176 12406 22228
rect 12618 22216 12624 22228
rect 12452 22188 12624 22216
rect 7147 22052 7972 22080
rect 7147 22049 7159 22052
rect 7101 22043 7159 22049
rect 8018 22040 8024 22092
rect 8076 22080 8082 22092
rect 11146 22080 11152 22092
rect 8076 22052 8121 22080
rect 10060 22052 11152 22080
rect 8076 22040 8082 22052
rect 10060 22024 10088 22052
rect 11146 22040 11152 22052
rect 11204 22040 11210 22092
rect 11885 22083 11943 22089
rect 11885 22049 11897 22083
rect 11931 22080 11943 22083
rect 12452 22080 12480 22188
rect 12618 22176 12624 22188
rect 12676 22216 12682 22228
rect 12713 22219 12771 22225
rect 12713 22216 12725 22219
rect 12676 22188 12725 22216
rect 12676 22176 12682 22188
rect 12713 22185 12725 22188
rect 12759 22185 12771 22219
rect 12713 22179 12771 22185
rect 13817 22219 13875 22225
rect 13817 22185 13829 22219
rect 13863 22216 13875 22219
rect 15102 22216 15108 22228
rect 13863 22188 15108 22216
rect 13863 22185 13875 22188
rect 13817 22179 13875 22185
rect 15102 22176 15108 22188
rect 15160 22216 15166 22228
rect 15378 22216 15384 22228
rect 15160 22188 15384 22216
rect 15160 22176 15166 22188
rect 15378 22176 15384 22188
rect 15436 22176 15442 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 16669 22219 16727 22225
rect 16669 22216 16681 22219
rect 16632 22188 16681 22216
rect 16632 22176 16638 22188
rect 16669 22185 16681 22188
rect 16715 22185 16727 22219
rect 17954 22216 17960 22228
rect 17915 22188 17960 22216
rect 16669 22179 16727 22185
rect 17954 22176 17960 22188
rect 18012 22176 18018 22228
rect 19889 22219 19947 22225
rect 19889 22185 19901 22219
rect 19935 22216 19947 22219
rect 20070 22216 20076 22228
rect 19935 22188 20076 22216
rect 19935 22185 19947 22188
rect 19889 22179 19947 22185
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 20254 22216 20260 22228
rect 20215 22188 20260 22216
rect 20254 22176 20260 22188
rect 20312 22176 20318 22228
rect 24118 22216 24124 22228
rect 24079 22188 24124 22216
rect 24118 22176 24124 22188
rect 24176 22216 24182 22228
rect 24578 22216 24584 22228
rect 24176 22188 24584 22216
rect 24176 22176 24182 22188
rect 24578 22176 24584 22188
rect 24636 22176 24642 22228
rect 12526 22108 12532 22160
rect 12584 22148 12590 22160
rect 22370 22157 22376 22160
rect 13357 22151 13415 22157
rect 13357 22148 13369 22151
rect 12584 22120 13369 22148
rect 12584 22108 12590 22120
rect 13357 22117 13369 22120
rect 13403 22117 13415 22151
rect 22364 22148 22376 22157
rect 22331 22120 22376 22148
rect 13357 22111 13415 22117
rect 22364 22111 22376 22120
rect 22370 22108 22376 22111
rect 22428 22108 22434 22160
rect 24210 22108 24216 22160
rect 24268 22148 24274 22160
rect 24397 22151 24455 22157
rect 24397 22148 24409 22151
rect 24268 22120 24409 22148
rect 24268 22108 24274 22120
rect 24397 22117 24409 22120
rect 24443 22117 24455 22151
rect 24397 22111 24455 22117
rect 11931 22052 12480 22080
rect 13909 22083 13967 22089
rect 11931 22049 11943 22052
rect 11885 22043 11943 22049
rect 13909 22049 13921 22083
rect 13955 22080 13967 22083
rect 13998 22080 14004 22092
rect 13955 22052 14004 22080
rect 13955 22049 13967 22052
rect 13909 22043 13967 22049
rect 13998 22040 14004 22052
rect 14056 22080 14062 22092
rect 14645 22083 14703 22089
rect 14645 22080 14657 22083
rect 14056 22052 14657 22080
rect 14056 22040 14062 22052
rect 14645 22049 14657 22052
rect 14691 22049 14703 22083
rect 14645 22043 14703 22049
rect 14826 22040 14832 22092
rect 14884 22080 14890 22092
rect 15194 22080 15200 22092
rect 14884 22052 15200 22080
rect 14884 22040 14890 22052
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15654 22080 15660 22092
rect 15344 22052 15660 22080
rect 15344 22040 15350 22052
rect 15654 22040 15660 22052
rect 15712 22040 15718 22092
rect 17037 22083 17095 22089
rect 17037 22049 17049 22083
rect 17083 22080 17095 22083
rect 17126 22080 17132 22092
rect 17083 22052 17132 22080
rect 17083 22049 17095 22052
rect 17037 22043 17095 22049
rect 17126 22040 17132 22052
rect 17184 22080 17190 22092
rect 17862 22080 17868 22092
rect 17184 22052 17868 22080
rect 17184 22040 17190 22052
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 19058 22080 19064 22092
rect 18739 22052 19064 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 19058 22040 19064 22052
rect 19116 22040 19122 22092
rect 20990 22080 20996 22092
rect 20951 22052 20996 22080
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 23382 22040 23388 22092
rect 23440 22040 23446 22092
rect 24949 22083 25007 22089
rect 24949 22049 24961 22083
rect 24995 22080 25007 22083
rect 26050 22080 26056 22092
rect 24995 22052 26056 22080
rect 24995 22049 25007 22052
rect 24949 22043 25007 22049
rect 26050 22040 26056 22052
rect 26108 22040 26114 22092
rect 3050 22012 3056 22024
rect 2963 21984 3056 22012
rect 3050 21972 3056 21984
rect 3108 21972 3114 22024
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4065 21947 4123 21953
rect 4065 21944 4077 21947
rect 2363 21916 4077 21944
rect 2363 21913 2375 21916
rect 2317 21907 2375 21913
rect 4065 21913 4077 21916
rect 4111 21913 4123 21947
rect 4065 21907 4123 21913
rect 4430 21904 4436 21956
rect 4488 21944 4494 21956
rect 4632 21944 4660 21975
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 6454 22012 6460 22024
rect 5224 21984 6460 22012
rect 5224 21972 5230 21984
rect 6454 21972 6460 21984
rect 6512 21972 6518 22024
rect 6641 22015 6699 22021
rect 6641 21981 6653 22015
rect 6687 22012 6699 22015
rect 6822 22012 6828 22024
rect 6687 21984 6828 22012
rect 6687 21981 6699 21984
rect 6641 21975 6699 21981
rect 6822 21972 6828 21984
rect 6880 21972 6886 22024
rect 8110 22012 8116 22024
rect 8071 21984 8116 22012
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 9493 22015 9551 22021
rect 9493 21981 9505 22015
rect 9539 22012 9551 22015
rect 9953 22015 10011 22021
rect 9953 22012 9965 22015
rect 9539 21984 9965 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 9953 21981 9965 21984
rect 9999 22012 10011 22015
rect 10042 22012 10048 22024
rect 9999 21984 10048 22012
rect 9999 21981 10011 21984
rect 9953 21975 10011 21981
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10502 22012 10508 22024
rect 10463 21984 10508 22012
rect 10502 21972 10508 21984
rect 10560 21972 10566 22024
rect 10686 22012 10692 22024
rect 10647 21984 10692 22012
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 22012 12311 22015
rect 12434 22012 12440 22024
rect 12299 21984 12440 22012
rect 12299 21981 12311 21984
rect 12253 21975 12311 21981
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 12805 22015 12863 22021
rect 12805 22012 12817 22015
rect 12492 21984 12817 22012
rect 12492 21972 12498 21984
rect 12805 21981 12817 21984
rect 12851 21981 12863 22015
rect 12986 22012 12992 22024
rect 12947 21984 12992 22012
rect 12805 21975 12863 21981
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 14182 22012 14188 22024
rect 14143 21984 14188 22012
rect 14182 21972 14188 21984
rect 14240 21972 14246 22024
rect 15749 22015 15807 22021
rect 15749 22012 15761 22015
rect 14660 21984 15761 22012
rect 14660 21956 14688 21984
rect 15749 21981 15761 21984
rect 15795 21981 15807 22015
rect 15930 22012 15936 22024
rect 15891 21984 15936 22012
rect 15749 21975 15807 21981
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 17310 22012 17316 22024
rect 17271 21984 17316 22012
rect 17310 21972 17316 21984
rect 17368 21972 17374 22024
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 18785 22015 18843 22021
rect 18785 22012 18797 22015
rect 17736 21984 18797 22012
rect 17736 21972 17742 21984
rect 18785 21981 18797 21984
rect 18831 21981 18843 22015
rect 18966 22012 18972 22024
rect 18927 21984 18972 22012
rect 18785 21975 18843 21981
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 22097 22015 22155 22021
rect 22097 22012 22109 22015
rect 21560 21984 22109 22012
rect 8941 21947 8999 21953
rect 8941 21944 8953 21947
rect 4488 21916 4660 21944
rect 7300 21916 8953 21944
rect 4488 21904 4494 21916
rect 7300 21888 7328 21916
rect 8941 21913 8953 21916
rect 8987 21913 8999 21947
rect 8941 21907 8999 21913
rect 14642 21904 14648 21956
rect 14700 21904 14706 21956
rect 15194 21904 15200 21956
rect 15252 21944 15258 21956
rect 15289 21947 15347 21953
rect 15289 21944 15301 21947
rect 15252 21916 15301 21944
rect 15252 21904 15258 21916
rect 15289 21913 15301 21916
rect 15335 21913 15347 21947
rect 18322 21944 18328 21956
rect 18283 21916 18328 21944
rect 15289 21907 15347 21913
rect 18322 21904 18328 21916
rect 18380 21904 18386 21956
rect 21177 21947 21235 21953
rect 21177 21913 21189 21947
rect 21223 21944 21235 21947
rect 21266 21944 21272 21956
rect 21223 21916 21272 21944
rect 21223 21913 21235 21916
rect 21177 21907 21235 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 3786 21876 3792 21888
rect 3292 21848 3792 21876
rect 3292 21836 3298 21848
rect 3786 21836 3792 21848
rect 3844 21876 3850 21888
rect 5077 21879 5135 21885
rect 5077 21876 5089 21879
rect 3844 21848 5089 21876
rect 3844 21836 3850 21848
rect 5077 21845 5089 21848
rect 5123 21876 5135 21879
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 5123 21848 5457 21876
rect 5123 21845 5135 21848
rect 5077 21839 5135 21845
rect 5445 21845 5457 21848
rect 5491 21876 5503 21879
rect 5534 21876 5540 21888
rect 5491 21848 5540 21876
rect 5491 21845 5503 21848
rect 5445 21839 5503 21845
rect 5534 21836 5540 21848
rect 5592 21876 5598 21888
rect 5813 21879 5871 21885
rect 5813 21876 5825 21879
rect 5592 21848 5825 21876
rect 5592 21836 5598 21848
rect 5813 21845 5825 21848
rect 5859 21876 5871 21879
rect 7282 21876 7288 21888
rect 5859 21848 7288 21876
rect 5859 21845 5871 21848
rect 5813 21839 5871 21845
rect 7282 21836 7288 21848
rect 7340 21836 7346 21888
rect 8662 21876 8668 21888
rect 8623 21848 8668 21876
rect 8662 21836 8668 21848
rect 8720 21836 8726 21888
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 11238 21876 11244 21888
rect 10091 21848 11244 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 11238 21836 11244 21848
rect 11296 21876 11302 21888
rect 11425 21879 11483 21885
rect 11425 21876 11437 21879
rect 11296 21848 11437 21876
rect 11296 21836 11302 21848
rect 11425 21845 11437 21848
rect 11471 21845 11483 21879
rect 11425 21839 11483 21845
rect 16114 21836 16120 21888
rect 16172 21876 16178 21888
rect 16301 21879 16359 21885
rect 16301 21876 16313 21879
rect 16172 21848 16313 21876
rect 16172 21836 16178 21848
rect 16301 21845 16313 21848
rect 16347 21845 16359 21879
rect 19426 21876 19432 21888
rect 19387 21848 19432 21876
rect 16301 21839 16359 21845
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 20254 21836 20260 21888
rect 20312 21876 20318 21888
rect 20533 21879 20591 21885
rect 20533 21876 20545 21879
rect 20312 21848 20545 21876
rect 20312 21836 20318 21848
rect 20533 21845 20545 21848
rect 20579 21876 20591 21879
rect 20898 21876 20904 21888
rect 20579 21848 20904 21876
rect 20579 21845 20591 21848
rect 20533 21839 20591 21845
rect 20898 21836 20904 21848
rect 20956 21876 20962 21888
rect 21560 21885 21588 21984
rect 22097 21981 22109 21984
rect 22143 21981 22155 22015
rect 22097 21975 22155 21981
rect 21545 21879 21603 21885
rect 21545 21876 21557 21879
rect 20956 21848 21557 21876
rect 20956 21836 20962 21848
rect 21545 21845 21557 21848
rect 21591 21845 21603 21879
rect 21545 21839 21603 21845
rect 22005 21879 22063 21885
rect 22005 21845 22017 21879
rect 22051 21876 22063 21879
rect 22278 21876 22284 21888
rect 22051 21848 22284 21876
rect 22051 21845 22063 21848
rect 22005 21839 22063 21845
rect 22278 21836 22284 21848
rect 22336 21876 22342 21888
rect 23400 21876 23428 22040
rect 25038 22012 25044 22024
rect 24999 21984 25044 22012
rect 25038 21972 25044 21984
rect 25096 21972 25102 22024
rect 25222 22012 25228 22024
rect 25183 21984 25228 22012
rect 25222 21972 25228 21984
rect 25280 21972 25286 22024
rect 25590 22012 25596 22024
rect 25551 21984 25596 22012
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 22336 21848 23428 21876
rect 22336 21836 22342 21848
rect 23474 21836 23480 21888
rect 23532 21876 23538 21888
rect 23532 21848 23577 21876
rect 23532 21836 23538 21848
rect 23750 21836 23756 21888
rect 23808 21876 23814 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23808 21848 24593 21876
rect 23808 21836 23814 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 2593 21675 2651 21681
rect 2593 21641 2605 21675
rect 2639 21672 2651 21675
rect 3050 21672 3056 21684
rect 2639 21644 3056 21672
rect 2639 21641 2651 21644
rect 2593 21635 2651 21641
rect 3050 21632 3056 21644
rect 3108 21632 3114 21684
rect 4522 21632 4528 21684
rect 4580 21672 4586 21684
rect 4985 21675 5043 21681
rect 4985 21672 4997 21675
rect 4580 21644 4997 21672
rect 4580 21632 4586 21644
rect 4985 21641 4997 21644
rect 5031 21641 5043 21675
rect 5350 21672 5356 21684
rect 5311 21644 5356 21672
rect 4985 21635 5043 21641
rect 5350 21632 5356 21644
rect 5408 21632 5414 21684
rect 6549 21675 6607 21681
rect 6549 21641 6561 21675
rect 6595 21672 6607 21675
rect 6822 21672 6828 21684
rect 6595 21644 6828 21672
rect 6595 21641 6607 21644
rect 6549 21635 6607 21641
rect 6822 21632 6828 21644
rect 6880 21672 6886 21684
rect 7653 21675 7711 21681
rect 7653 21672 7665 21675
rect 6880 21644 7665 21672
rect 6880 21632 6886 21644
rect 7653 21641 7665 21644
rect 7699 21672 7711 21675
rect 8110 21672 8116 21684
rect 7699 21644 8116 21672
rect 7699 21641 7711 21644
rect 7653 21635 7711 21641
rect 8110 21632 8116 21644
rect 8168 21632 8174 21684
rect 9122 21672 9128 21684
rect 9035 21644 9128 21672
rect 9122 21632 9128 21644
rect 9180 21672 9186 21684
rect 9582 21672 9588 21684
rect 9180 21644 9588 21672
rect 9180 21632 9186 21644
rect 9582 21632 9588 21644
rect 9640 21632 9646 21684
rect 10134 21672 10140 21684
rect 10095 21644 10140 21672
rect 10134 21632 10140 21644
rect 10192 21632 10198 21684
rect 10502 21672 10508 21684
rect 10463 21644 10508 21672
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 12250 21672 12256 21684
rect 12211 21644 12256 21672
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 13998 21672 14004 21684
rect 12492 21644 12537 21672
rect 13959 21644 14004 21672
rect 12492 21632 12498 21644
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 14182 21632 14188 21684
rect 14240 21672 14246 21684
rect 14366 21672 14372 21684
rect 14240 21644 14372 21672
rect 14240 21632 14246 21644
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 14458 21632 14464 21684
rect 14516 21632 14522 21684
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 15013 21675 15071 21681
rect 15013 21672 15025 21675
rect 14700 21644 15025 21672
rect 14700 21632 14706 21644
rect 15013 21641 15025 21644
rect 15059 21641 15071 21675
rect 15013 21635 15071 21641
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 16206 21672 16212 21684
rect 15988 21644 16212 21672
rect 15988 21632 15994 21644
rect 16206 21632 16212 21644
rect 16264 21672 16270 21684
rect 16945 21675 17003 21681
rect 16945 21672 16957 21675
rect 16264 21644 16957 21672
rect 16264 21632 16270 21644
rect 16945 21641 16957 21644
rect 16991 21641 17003 21675
rect 16945 21635 17003 21641
rect 17497 21675 17555 21681
rect 17497 21641 17509 21675
rect 17543 21672 17555 21675
rect 18966 21672 18972 21684
rect 17543 21644 18972 21672
rect 17543 21641 17555 21644
rect 17497 21635 17555 21641
rect 18966 21632 18972 21644
rect 19024 21632 19030 21684
rect 19150 21632 19156 21684
rect 19208 21672 19214 21684
rect 20165 21675 20223 21681
rect 20165 21672 20177 21675
rect 19208 21644 20177 21672
rect 19208 21632 19214 21644
rect 20165 21641 20177 21644
rect 20211 21641 20223 21675
rect 22002 21672 22008 21684
rect 21963 21644 22008 21672
rect 20165 21635 20223 21641
rect 22002 21632 22008 21644
rect 22060 21632 22066 21684
rect 25222 21632 25228 21684
rect 25280 21672 25286 21684
rect 25961 21675 26019 21681
rect 25961 21672 25973 21675
rect 25280 21644 25973 21672
rect 25280 21632 25286 21644
rect 25961 21641 25973 21644
rect 26007 21641 26019 21675
rect 25961 21635 26019 21641
rect 2314 21604 2320 21616
rect 2056 21576 2320 21604
rect 2056 21545 2084 21576
rect 2314 21564 2320 21576
rect 2372 21604 2378 21616
rect 2372 21576 3004 21604
rect 2372 21564 2378 21576
rect 2976 21545 3004 21576
rect 12802 21564 12808 21616
rect 12860 21604 12866 21616
rect 14476 21604 14504 21632
rect 12860 21576 13032 21604
rect 14476 21576 14688 21604
rect 12860 21564 12866 21576
rect 13004 21548 13032 21576
rect 14660 21548 14688 21576
rect 17678 21564 17684 21616
rect 17736 21604 17742 21616
rect 17773 21607 17831 21613
rect 17773 21604 17785 21607
rect 17736 21576 17785 21604
rect 17736 21564 17742 21576
rect 17773 21573 17785 21576
rect 17819 21604 17831 21607
rect 18138 21604 18144 21616
rect 17819 21576 18144 21604
rect 17819 21573 17831 21576
rect 17773 21567 17831 21573
rect 18138 21564 18144 21576
rect 18196 21564 18202 21616
rect 21913 21607 21971 21613
rect 21913 21573 21925 21607
rect 21959 21604 21971 21607
rect 22370 21604 22376 21616
rect 21959 21576 22376 21604
rect 21959 21573 21971 21576
rect 21913 21567 21971 21573
rect 22370 21564 22376 21576
rect 22428 21564 22434 21616
rect 23109 21607 23167 21613
rect 23109 21604 23121 21607
rect 22480 21576 23121 21604
rect 2041 21539 2099 21545
rect 2041 21505 2053 21539
rect 2087 21505 2099 21539
rect 2041 21499 2099 21505
rect 2961 21539 3019 21545
rect 2961 21505 2973 21539
rect 3007 21536 3019 21539
rect 3007 21508 3188 21536
rect 3007 21505 3019 21508
rect 2961 21499 3019 21505
rect 3050 21468 3056 21480
rect 3011 21440 3056 21468
rect 3050 21428 3056 21440
rect 3108 21428 3114 21480
rect 3160 21468 3188 21508
rect 7282 21496 7288 21548
rect 7340 21536 7346 21548
rect 7745 21539 7803 21545
rect 7745 21536 7757 21539
rect 7340 21508 7757 21536
rect 7340 21496 7346 21508
rect 7745 21505 7757 21508
rect 7791 21505 7803 21539
rect 11238 21536 11244 21548
rect 11199 21508 11244 21536
rect 7745 21499 7803 21505
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 11425 21539 11483 21545
rect 11425 21505 11437 21539
rect 11471 21536 11483 21539
rect 11882 21536 11888 21548
rect 11471 21508 11888 21536
rect 11471 21505 11483 21508
rect 11425 21499 11483 21505
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 12894 21536 12900 21548
rect 12855 21508 12900 21536
rect 12894 21496 12900 21508
rect 12952 21496 12958 21548
rect 12986 21496 12992 21548
rect 13044 21536 13050 21548
rect 13044 21508 13089 21536
rect 13044 21496 13050 21508
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14056 21508 14565 21536
rect 14056 21496 14062 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 14642 21496 14648 21548
rect 14700 21496 14706 21548
rect 16114 21536 16120 21548
rect 16075 21508 16120 21536
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 22480 21545 22508 21576
rect 23109 21573 23121 21576
rect 23155 21604 23167 21607
rect 23155 21576 23428 21604
rect 23155 21573 23167 21576
rect 23109 21567 23167 21573
rect 22465 21539 22523 21545
rect 22465 21505 22477 21539
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21536 22707 21539
rect 22695 21508 23336 21536
rect 22695 21505 22707 21508
rect 22649 21499 22707 21505
rect 3320 21471 3378 21477
rect 3320 21468 3332 21471
rect 3160 21440 3332 21468
rect 3320 21437 3332 21440
rect 3366 21468 3378 21471
rect 3602 21468 3608 21480
rect 3366 21440 3608 21468
rect 3366 21437 3378 21440
rect 3320 21431 3378 21437
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 5350 21428 5356 21480
rect 5408 21468 5414 21480
rect 5537 21471 5595 21477
rect 5537 21468 5549 21471
rect 5408 21440 5549 21468
rect 5408 21428 5414 21440
rect 5537 21437 5549 21440
rect 5583 21437 5595 21471
rect 5537 21431 5595 21437
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12768 21440 12817 21468
rect 12768 21428 12774 21440
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 13449 21471 13507 21477
rect 13449 21468 13461 21471
rect 12851 21440 13461 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 13449 21437 13461 21440
rect 13495 21437 13507 21471
rect 16025 21471 16083 21477
rect 16025 21468 16037 21471
rect 13449 21431 13507 21437
rect 15396 21440 16037 21468
rect 1949 21403 2007 21409
rect 1949 21369 1961 21403
rect 1995 21400 2007 21403
rect 2038 21400 2044 21412
rect 1995 21372 2044 21400
rect 1995 21369 2007 21372
rect 1949 21363 2007 21369
rect 2038 21360 2044 21372
rect 2096 21360 2102 21412
rect 7285 21403 7343 21409
rect 7285 21369 7297 21403
rect 7331 21400 7343 21403
rect 8012 21403 8070 21409
rect 8012 21400 8024 21403
rect 7331 21372 8024 21400
rect 7331 21369 7343 21372
rect 7285 21363 7343 21369
rect 8012 21369 8024 21372
rect 8058 21400 8070 21403
rect 8110 21400 8116 21412
rect 8058 21372 8116 21400
rect 8058 21369 8070 21372
rect 8012 21363 8070 21369
rect 8110 21360 8116 21372
rect 8168 21360 8174 21412
rect 9769 21403 9827 21409
rect 9769 21369 9781 21403
rect 9815 21400 9827 21403
rect 10686 21400 10692 21412
rect 9815 21372 10692 21400
rect 9815 21369 9827 21372
rect 9769 21363 9827 21369
rect 10686 21360 10692 21372
rect 10744 21360 10750 21412
rect 11146 21400 11152 21412
rect 11059 21372 11152 21400
rect 11146 21360 11152 21372
rect 11204 21400 11210 21412
rect 12342 21400 12348 21412
rect 11204 21372 12348 21400
rect 11204 21360 11210 21372
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 14090 21360 14096 21412
rect 14148 21400 14154 21412
rect 14461 21403 14519 21409
rect 14461 21400 14473 21403
rect 14148 21372 14473 21400
rect 14148 21360 14154 21372
rect 14461 21369 14473 21372
rect 14507 21369 14519 21403
rect 14461 21363 14519 21369
rect 15396 21344 15424 21440
rect 16025 21437 16037 21440
rect 16071 21437 16083 21471
rect 16025 21431 16083 21437
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18322 21468 18328 21480
rect 18104 21440 18328 21468
rect 18104 21428 18110 21440
rect 18322 21428 18328 21440
rect 18380 21468 18386 21480
rect 18785 21471 18843 21477
rect 18785 21468 18797 21471
rect 18380 21440 18797 21468
rect 18380 21428 18386 21440
rect 18785 21437 18797 21440
rect 18831 21437 18843 21471
rect 18785 21431 18843 21437
rect 19052 21471 19110 21477
rect 19052 21437 19064 21471
rect 19098 21468 19110 21471
rect 19426 21468 19432 21480
rect 19098 21440 19432 21468
rect 19098 21437 19110 21440
rect 19052 21431 19110 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 22278 21428 22284 21480
rect 22336 21468 22342 21480
rect 22373 21471 22431 21477
rect 22373 21468 22385 21471
rect 22336 21440 22385 21468
rect 22336 21428 22342 21440
rect 22373 21437 22385 21440
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 15930 21400 15936 21412
rect 15891 21372 15936 21400
rect 15930 21360 15936 21372
rect 15988 21400 15994 21412
rect 16577 21403 16635 21409
rect 16577 21400 16589 21403
rect 15988 21372 16589 21400
rect 15988 21360 15994 21372
rect 16577 21369 16589 21372
rect 16623 21369 16635 21403
rect 16577 21363 16635 21369
rect 21545 21403 21603 21409
rect 21545 21369 21557 21403
rect 21591 21400 21603 21403
rect 22664 21400 22692 21499
rect 21591 21372 22692 21400
rect 21591 21369 21603 21372
rect 21545 21363 21603 21369
rect 1486 21332 1492 21344
rect 1447 21304 1492 21332
rect 1486 21292 1492 21304
rect 1544 21292 1550 21344
rect 1857 21335 1915 21341
rect 1857 21301 1869 21335
rect 1903 21332 1915 21335
rect 2130 21332 2136 21344
rect 1903 21304 2136 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 2130 21292 2136 21304
rect 2188 21292 2194 21344
rect 4430 21332 4436 21344
rect 4391 21304 4436 21332
rect 4430 21292 4436 21304
rect 4488 21292 4494 21344
rect 5718 21332 5724 21344
rect 5679 21304 5724 21332
rect 5718 21292 5724 21304
rect 5776 21292 5782 21344
rect 6086 21332 6092 21344
rect 6047 21304 6092 21332
rect 6086 21292 6092 21304
rect 6144 21292 6150 21344
rect 10778 21332 10784 21344
rect 10739 21304 10784 21332
rect 10778 21292 10784 21304
rect 10836 21292 10842 21344
rect 11882 21332 11888 21344
rect 11843 21304 11888 21332
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 13909 21335 13967 21341
rect 13909 21301 13921 21335
rect 13955 21332 13967 21335
rect 13998 21332 14004 21344
rect 13955 21304 14004 21332
rect 13955 21301 13967 21304
rect 13909 21295 13967 21301
rect 13998 21292 14004 21304
rect 14056 21292 14062 21344
rect 14366 21332 14372 21344
rect 14327 21304 14372 21332
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 15378 21332 15384 21344
rect 15339 21304 15384 21332
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15528 21304 15577 21332
rect 15528 21292 15534 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 18414 21332 18420 21344
rect 18327 21304 18420 21332
rect 15565 21295 15623 21301
rect 18414 21292 18420 21304
rect 18472 21332 18478 21344
rect 19058 21332 19064 21344
rect 18472 21304 19064 21332
rect 18472 21292 18478 21304
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 20990 21292 20996 21344
rect 21048 21332 21054 21344
rect 21085 21335 21143 21341
rect 21085 21332 21097 21335
rect 21048 21304 21097 21332
rect 21048 21292 21054 21304
rect 21085 21301 21097 21304
rect 21131 21332 21143 21335
rect 21174 21332 21180 21344
rect 21131 21304 21180 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 23308 21332 23336 21508
rect 23400 21468 23428 21576
rect 23658 21536 23664 21548
rect 23619 21508 23664 21536
rect 23658 21496 23664 21508
rect 23716 21496 23722 21548
rect 23750 21468 23756 21480
rect 23400 21440 23756 21468
rect 23750 21428 23756 21440
rect 23808 21428 23814 21480
rect 23928 21471 23986 21477
rect 23928 21437 23940 21471
rect 23974 21468 23986 21471
rect 25222 21468 25228 21480
rect 23974 21440 25228 21468
rect 23974 21437 23986 21440
rect 23928 21431 23986 21437
rect 23474 21400 23480 21412
rect 23387 21372 23480 21400
rect 23474 21360 23480 21372
rect 23532 21400 23538 21412
rect 23943 21400 23971 21431
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 23532 21372 23971 21400
rect 23532 21360 23538 21372
rect 23750 21332 23756 21344
rect 23308 21304 23756 21332
rect 23750 21292 23756 21304
rect 23808 21332 23814 21344
rect 25041 21335 25099 21341
rect 25041 21332 25053 21335
rect 23808 21304 25053 21332
rect 23808 21292 23814 21304
rect 25041 21301 25053 21304
rect 25087 21301 25099 21335
rect 25041 21295 25099 21301
rect 25685 21335 25743 21341
rect 25685 21301 25697 21335
rect 25731 21332 25743 21335
rect 26050 21332 26056 21344
rect 25731 21304 26056 21332
rect 25731 21301 25743 21304
rect 25685 21295 25743 21301
rect 26050 21292 26056 21304
rect 26108 21292 26114 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1394 21128 1400 21140
rect 1355 21100 1400 21128
rect 1394 21088 1400 21100
rect 1452 21088 1458 21140
rect 2314 21128 2320 21140
rect 2275 21100 2320 21128
rect 2314 21088 2320 21100
rect 2372 21088 2378 21140
rect 2409 21131 2467 21137
rect 2409 21097 2421 21131
rect 2455 21128 2467 21131
rect 3142 21128 3148 21140
rect 2455 21100 3148 21128
rect 2455 21097 2467 21100
rect 2409 21091 2467 21097
rect 3142 21088 3148 21100
rect 3200 21088 3206 21140
rect 4614 21128 4620 21140
rect 4575 21100 4620 21128
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 6273 21131 6331 21137
rect 6273 21097 6285 21131
rect 6319 21097 6331 21131
rect 6273 21091 6331 21097
rect 3602 21020 3608 21072
rect 3660 21060 3666 21072
rect 6288 21060 6316 21091
rect 6454 21088 6460 21140
rect 6512 21128 6518 21140
rect 6825 21131 6883 21137
rect 6825 21128 6837 21131
rect 6512 21100 6837 21128
rect 6512 21088 6518 21100
rect 6825 21097 6837 21100
rect 6871 21097 6883 21131
rect 7742 21128 7748 21140
rect 7703 21100 7748 21128
rect 6825 21091 6883 21097
rect 7742 21088 7748 21100
rect 7800 21088 7806 21140
rect 7834 21088 7840 21140
rect 7892 21128 7898 21140
rect 7892 21100 7937 21128
rect 7892 21088 7898 21100
rect 8018 21088 8024 21140
rect 8076 21128 8082 21140
rect 8389 21131 8447 21137
rect 8389 21128 8401 21131
rect 8076 21100 8401 21128
rect 8076 21088 8082 21100
rect 8389 21097 8401 21100
rect 8435 21097 8447 21131
rect 8389 21091 8447 21097
rect 10505 21131 10563 21137
rect 10505 21097 10517 21131
rect 10551 21128 10563 21131
rect 11146 21128 11152 21140
rect 10551 21100 11152 21128
rect 10551 21097 10563 21100
rect 10505 21091 10563 21097
rect 11146 21088 11152 21100
rect 11204 21088 11210 21140
rect 11882 21088 11888 21140
rect 11940 21128 11946 21140
rect 11977 21131 12035 21137
rect 11977 21128 11989 21131
rect 11940 21100 11989 21128
rect 11940 21088 11946 21100
rect 11977 21097 11989 21100
rect 12023 21097 12035 21131
rect 12894 21128 12900 21140
rect 12855 21100 12900 21128
rect 11977 21091 12035 21097
rect 12894 21088 12900 21100
rect 12952 21088 12958 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 14090 21128 14096 21140
rect 14051 21100 14096 21128
rect 14090 21088 14096 21100
rect 14148 21088 14154 21140
rect 15105 21131 15163 21137
rect 15105 21097 15117 21131
rect 15151 21128 15163 21131
rect 15286 21128 15292 21140
rect 15151 21100 15292 21128
rect 15151 21097 15163 21100
rect 15105 21091 15163 21097
rect 15286 21088 15292 21100
rect 15344 21088 15350 21140
rect 15565 21131 15623 21137
rect 15565 21097 15577 21131
rect 15611 21128 15623 21131
rect 15654 21128 15660 21140
rect 15611 21100 15660 21128
rect 15611 21097 15623 21100
rect 15565 21091 15623 21097
rect 15654 21088 15660 21100
rect 15712 21088 15718 21140
rect 17034 21128 17040 21140
rect 16995 21100 17040 21128
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 17126 21088 17132 21140
rect 17184 21128 17190 21140
rect 17589 21131 17647 21137
rect 17589 21128 17601 21131
rect 17184 21100 17601 21128
rect 17184 21088 17190 21100
rect 17589 21097 17601 21100
rect 17635 21097 17647 21131
rect 17589 21091 17647 21097
rect 18598 21088 18604 21140
rect 18656 21128 18662 21140
rect 18966 21128 18972 21140
rect 18656 21100 18972 21128
rect 18656 21088 18662 21100
rect 18966 21088 18972 21100
rect 19024 21128 19030 21140
rect 19153 21131 19211 21137
rect 19153 21128 19165 21131
rect 19024 21100 19165 21128
rect 19024 21088 19030 21100
rect 19153 21097 19165 21100
rect 19199 21097 19211 21131
rect 19153 21091 19211 21097
rect 19334 21088 19340 21140
rect 19392 21128 19398 21140
rect 19889 21131 19947 21137
rect 19889 21128 19901 21131
rect 19392 21100 19901 21128
rect 19392 21088 19398 21100
rect 19889 21097 19901 21100
rect 19935 21097 19947 21131
rect 20714 21128 20720 21140
rect 20675 21100 20720 21128
rect 19889 21091 19947 21097
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 20901 21131 20959 21137
rect 20901 21097 20913 21131
rect 20947 21097 20959 21131
rect 20901 21091 20959 21097
rect 22465 21131 22523 21137
rect 22465 21097 22477 21131
rect 22511 21128 22523 21131
rect 23382 21128 23388 21140
rect 22511 21100 23388 21128
rect 22511 21097 22523 21100
rect 22465 21091 22523 21097
rect 3660 21032 6316 21060
rect 12621 21063 12679 21069
rect 3660 21020 3666 21032
rect 12621 21029 12633 21063
rect 12667 21060 12679 21063
rect 12986 21060 12992 21072
rect 12667 21032 12992 21060
rect 12667 21029 12679 21032
rect 12621 21023 12679 21029
rect 12986 21020 12992 21032
rect 13044 21020 13050 21072
rect 2682 20952 2688 21004
rect 2740 20992 2746 21004
rect 5166 21001 5172 21004
rect 2777 20995 2835 21001
rect 2777 20992 2789 20995
rect 2740 20964 2789 20992
rect 2740 20952 2746 20964
rect 2777 20961 2789 20964
rect 2823 20992 2835 20995
rect 3421 20995 3479 21001
rect 3421 20992 3433 20995
rect 2823 20964 3433 20992
rect 2823 20961 2835 20964
rect 2777 20955 2835 20961
rect 3421 20961 3433 20964
rect 3467 20961 3479 20995
rect 5160 20992 5172 21001
rect 5127 20964 5172 20992
rect 3421 20955 3479 20961
rect 5160 20955 5172 20964
rect 5166 20952 5172 20955
rect 5224 20952 5230 21004
rect 10686 20952 10692 21004
rect 10744 20992 10750 21004
rect 10864 20995 10922 21001
rect 10864 20992 10876 20995
rect 10744 20964 10876 20992
rect 10744 20952 10750 20964
rect 10864 20961 10876 20964
rect 10910 20992 10922 20995
rect 11146 20992 11152 21004
rect 10910 20964 11152 20992
rect 10910 20961 10922 20964
rect 10864 20955 10922 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 12802 20952 12808 21004
rect 12860 20992 12866 21004
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 12860 20964 13461 20992
rect 12860 20952 12866 20964
rect 13449 20961 13461 20964
rect 13495 20961 13507 20995
rect 13449 20955 13507 20961
rect 13541 20995 13599 21001
rect 13541 20961 13553 20995
rect 13587 20992 13599 20995
rect 13722 20992 13728 21004
rect 13587 20964 13728 20992
rect 13587 20961 13599 20964
rect 13541 20955 13599 20961
rect 13722 20952 13728 20964
rect 13780 20952 13786 21004
rect 15304 20992 15332 21088
rect 18049 21063 18107 21069
rect 18049 21029 18061 21063
rect 18095 21060 18107 21063
rect 18509 21063 18567 21069
rect 18509 21060 18521 21063
rect 18095 21032 18521 21060
rect 18095 21029 18107 21032
rect 18049 21023 18107 21029
rect 18509 21029 18521 21032
rect 18555 21060 18567 21063
rect 20916 21060 20944 21091
rect 23382 21088 23388 21100
rect 23440 21088 23446 21140
rect 23658 21128 23664 21140
rect 23492 21100 23664 21128
rect 18555 21032 20944 21060
rect 23017 21063 23075 21069
rect 18555 21029 18567 21032
rect 18509 21023 18567 21029
rect 23017 21029 23029 21063
rect 23063 21060 23075 21063
rect 23106 21060 23112 21072
rect 23063 21032 23112 21060
rect 23063 21029 23075 21032
rect 23017 21023 23075 21029
rect 23106 21020 23112 21032
rect 23164 21060 23170 21072
rect 23293 21063 23351 21069
rect 23293 21060 23305 21063
rect 23164 21032 23305 21060
rect 23164 21020 23170 21032
rect 23293 21029 23305 21032
rect 23339 21060 23351 21063
rect 23492 21060 23520 21100
rect 23658 21088 23664 21100
rect 23716 21088 23722 21140
rect 25038 21088 25044 21140
rect 25096 21128 25102 21140
rect 25409 21131 25467 21137
rect 25409 21128 25421 21131
rect 25096 21100 25421 21128
rect 25096 21088 25102 21100
rect 25409 21097 25421 21100
rect 25455 21097 25467 21131
rect 25409 21091 25467 21097
rect 23750 21069 23756 21072
rect 23744 21060 23756 21069
rect 23339 21032 23520 21060
rect 23711 21032 23756 21060
rect 23339 21029 23351 21032
rect 23293 21023 23351 21029
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15304 20964 15669 20992
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15924 20995 15982 21001
rect 15924 20961 15936 20995
rect 15970 20992 15982 20995
rect 16482 20992 16488 21004
rect 15970 20964 16488 20992
rect 15970 20961 15982 20964
rect 15924 20955 15982 20961
rect 16482 20952 16488 20964
rect 16540 20952 16546 21004
rect 18414 20952 18420 21004
rect 18472 20992 18478 21004
rect 18601 20995 18659 21001
rect 18601 20992 18613 20995
rect 18472 20964 18613 20992
rect 18472 20952 18478 20964
rect 18601 20961 18613 20964
rect 18647 20961 18659 20995
rect 18601 20955 18659 20961
rect 19705 20995 19763 21001
rect 19705 20961 19717 20995
rect 19751 20992 19763 20995
rect 20162 20992 20168 21004
rect 19751 20964 20168 20992
rect 19751 20961 19763 20964
rect 19705 20955 19763 20961
rect 20162 20952 20168 20964
rect 20220 20952 20226 21004
rect 20714 20952 20720 21004
rect 20772 20992 20778 21004
rect 23492 21001 23520 21032
rect 23744 21023 23756 21032
rect 23750 21020 23756 21023
rect 23808 21020 23814 21072
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 20772 20964 21281 20992
rect 20772 20952 20778 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 21269 20955 21327 20961
rect 23477 20995 23535 21001
rect 23477 20961 23489 20995
rect 23523 20992 23535 20995
rect 23523 20964 23557 20992
rect 23523 20961 23535 20964
rect 23477 20955 23535 20961
rect 2590 20884 2596 20936
rect 2648 20924 2654 20936
rect 2869 20927 2927 20933
rect 2869 20924 2881 20927
rect 2648 20896 2881 20924
rect 2648 20884 2654 20896
rect 2869 20893 2881 20896
rect 2915 20893 2927 20927
rect 2869 20887 2927 20893
rect 2961 20927 3019 20933
rect 2961 20893 2973 20927
rect 3007 20924 3019 20927
rect 4249 20927 4307 20933
rect 4249 20924 4261 20927
rect 3007 20896 4261 20924
rect 3007 20893 3019 20896
rect 2961 20887 3019 20893
rect 4249 20893 4261 20896
rect 4295 20924 4307 20927
rect 4430 20924 4436 20936
rect 4295 20896 4436 20924
rect 4295 20893 4307 20896
rect 4249 20887 4307 20893
rect 2774 20816 2780 20868
rect 2832 20856 2838 20868
rect 2976 20856 3004 20887
rect 4430 20884 4436 20896
rect 4488 20884 4494 20936
rect 4893 20927 4951 20933
rect 4893 20893 4905 20927
rect 4939 20893 4951 20927
rect 4893 20887 4951 20893
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7926 20924 7932 20936
rect 7331 20896 7932 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 4908 20856 4936 20887
rect 7926 20884 7932 20896
rect 7984 20884 7990 20936
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10597 20927 10655 20933
rect 10597 20924 10609 20927
rect 10192 20896 10609 20924
rect 10192 20884 10198 20896
rect 10597 20893 10609 20896
rect 10643 20893 10655 20927
rect 10597 20887 10655 20893
rect 11974 20884 11980 20936
rect 12032 20924 12038 20936
rect 13633 20927 13691 20933
rect 13633 20924 13645 20927
rect 12032 20896 13645 20924
rect 12032 20884 12038 20896
rect 13633 20893 13645 20896
rect 13679 20924 13691 20927
rect 14274 20924 14280 20936
rect 13679 20896 14280 20924
rect 13679 20893 13691 20896
rect 13633 20887 13691 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 18690 20884 18696 20936
rect 18748 20924 18754 20936
rect 18748 20896 18793 20924
rect 18748 20884 18754 20896
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21358 20924 21364 20936
rect 21140 20896 21364 20924
rect 21140 20884 21146 20896
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 2832 20828 3004 20856
rect 4264 20828 4936 20856
rect 8849 20859 8907 20865
rect 2832 20816 2838 20828
rect 4264 20800 4292 20828
rect 8849 20825 8861 20859
rect 8895 20856 8907 20859
rect 9490 20856 9496 20868
rect 8895 20828 9496 20856
rect 8895 20825 8907 20828
rect 8849 20819 8907 20825
rect 9490 20816 9496 20828
rect 9548 20816 9554 20868
rect 11698 20816 11704 20868
rect 11756 20856 11762 20868
rect 14826 20856 14832 20868
rect 11756 20828 14832 20856
rect 11756 20816 11762 20828
rect 14826 20816 14832 20828
rect 14884 20816 14890 20868
rect 18322 20816 18328 20868
rect 18380 20856 18386 20868
rect 19521 20859 19579 20865
rect 19521 20856 19533 20859
rect 18380 20828 19533 20856
rect 18380 20816 18386 20828
rect 19521 20825 19533 20828
rect 19567 20856 19579 20859
rect 20254 20856 20260 20868
rect 19567 20828 20260 20856
rect 19567 20825 19579 20828
rect 19521 20819 19579 20825
rect 20254 20816 20260 20828
rect 20312 20856 20318 20868
rect 20806 20856 20812 20868
rect 20312 20828 20812 20856
rect 20312 20816 20318 20828
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 20898 20816 20904 20868
rect 20956 20856 20962 20868
rect 21468 20856 21496 20887
rect 23106 20856 23112 20868
rect 20956 20828 21496 20856
rect 21560 20828 23112 20856
rect 20956 20816 20962 20828
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 2130 20788 2136 20800
rect 1995 20760 2136 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 2130 20748 2136 20760
rect 2188 20748 2194 20800
rect 3050 20748 3056 20800
rect 3108 20788 3114 20800
rect 3786 20788 3792 20800
rect 3108 20760 3792 20788
rect 3108 20748 3114 20760
rect 3786 20748 3792 20760
rect 3844 20788 3850 20800
rect 3881 20791 3939 20797
rect 3881 20788 3893 20791
rect 3844 20760 3893 20788
rect 3844 20748 3850 20760
rect 3881 20757 3893 20760
rect 3927 20788 3939 20791
rect 4246 20788 4252 20800
rect 3927 20760 4252 20788
rect 3927 20757 3939 20760
rect 3881 20751 3939 20757
rect 4246 20748 4252 20760
rect 4304 20748 4310 20800
rect 7282 20748 7288 20800
rect 7340 20788 7346 20800
rect 7377 20791 7435 20797
rect 7377 20788 7389 20791
rect 7340 20760 7389 20788
rect 7340 20748 7346 20760
rect 7377 20757 7389 20760
rect 7423 20757 7435 20791
rect 7377 20751 7435 20757
rect 9030 20748 9036 20800
rect 9088 20788 9094 20800
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 9088 20760 9137 20788
rect 9088 20748 9094 20760
rect 9125 20757 9137 20760
rect 9171 20788 9183 20791
rect 9861 20791 9919 20797
rect 9861 20788 9873 20791
rect 9171 20760 9873 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9861 20757 9873 20760
rect 9907 20757 9919 20791
rect 14458 20788 14464 20800
rect 14419 20760 14464 20788
rect 9861 20751 9919 20757
rect 14458 20748 14464 20760
rect 14516 20748 14522 20800
rect 14844 20788 14872 20816
rect 16298 20788 16304 20800
rect 14844 20760 16304 20788
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 19242 20788 19248 20800
rect 18187 20760 19248 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 20824 20788 20852 20816
rect 21560 20788 21588 20828
rect 23106 20816 23112 20828
rect 23164 20816 23170 20868
rect 24578 20816 24584 20868
rect 24636 20816 24642 20868
rect 20824 20760 21588 20788
rect 22097 20791 22155 20797
rect 22097 20757 22109 20791
rect 22143 20788 22155 20791
rect 22278 20788 22284 20800
rect 22143 20760 22284 20788
rect 22143 20757 22155 20760
rect 22097 20751 22155 20757
rect 22278 20748 22284 20760
rect 22336 20748 22342 20800
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 24596 20788 24624 20816
rect 24854 20788 24860 20800
rect 23532 20760 24624 20788
rect 24815 20760 24860 20788
rect 23532 20748 23538 20760
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2682 20584 2688 20596
rect 2639 20556 2688 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 7653 20587 7711 20593
rect 7653 20553 7665 20587
rect 7699 20584 7711 20587
rect 7742 20584 7748 20596
rect 7699 20556 7748 20584
rect 7699 20553 7711 20556
rect 7653 20547 7711 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 7834 20544 7840 20596
rect 7892 20584 7898 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 7892 20556 7941 20584
rect 7892 20544 7898 20556
rect 7929 20553 7941 20556
rect 7975 20553 7987 20587
rect 10778 20584 10784 20596
rect 10739 20556 10784 20584
rect 7929 20547 7987 20553
rect 10778 20544 10784 20556
rect 10836 20544 10842 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11885 20587 11943 20593
rect 11885 20584 11897 20587
rect 11204 20556 11897 20584
rect 11204 20544 11210 20556
rect 11885 20553 11897 20556
rect 11931 20584 11943 20587
rect 14274 20584 14280 20596
rect 11931 20556 12756 20584
rect 14235 20556 14280 20584
rect 11931 20553 11943 20556
rect 11885 20547 11943 20553
rect 4246 20476 4252 20528
rect 4304 20516 4310 20528
rect 6457 20519 6515 20525
rect 6457 20516 6469 20519
rect 4304 20488 6469 20516
rect 4304 20476 4310 20488
rect 6457 20485 6469 20488
rect 6503 20516 6515 20519
rect 10321 20519 10379 20525
rect 6503 20488 8156 20516
rect 6503 20485 6515 20488
rect 6457 20479 6515 20485
rect 8128 20460 8156 20488
rect 10321 20485 10333 20519
rect 10367 20516 10379 20519
rect 11164 20516 11192 20544
rect 10367 20488 11192 20516
rect 10367 20485 10379 20488
rect 10321 20479 10379 20485
rect 11238 20476 11244 20528
rect 11296 20516 11302 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 11296 20488 12449 20516
rect 11296 20476 11302 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12437 20479 12495 20485
rect 12728 20460 12756 20556
rect 14274 20544 14280 20556
rect 14332 20544 14338 20596
rect 14642 20544 14648 20596
rect 14700 20584 14706 20596
rect 15654 20584 15660 20596
rect 14700 20556 15660 20584
rect 14700 20544 14706 20556
rect 15654 20544 15660 20556
rect 15712 20584 15718 20596
rect 16025 20587 16083 20593
rect 16025 20584 16037 20587
rect 15712 20556 16037 20584
rect 15712 20544 15718 20556
rect 16025 20553 16037 20556
rect 16071 20553 16083 20587
rect 16666 20584 16672 20596
rect 16579 20556 16672 20584
rect 16025 20547 16083 20553
rect 16666 20544 16672 20556
rect 16724 20584 16730 20596
rect 18325 20587 18383 20593
rect 18325 20584 18337 20587
rect 16724 20556 18337 20584
rect 16724 20544 16730 20556
rect 18325 20553 18337 20556
rect 18371 20584 18383 20587
rect 18690 20584 18696 20596
rect 18371 20556 18696 20584
rect 18371 20553 18383 20556
rect 18325 20547 18383 20553
rect 18690 20544 18696 20556
rect 18748 20544 18754 20596
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 20073 20587 20131 20593
rect 20073 20584 20085 20587
rect 19484 20556 20085 20584
rect 19484 20544 19490 20556
rect 20073 20553 20085 20556
rect 20119 20553 20131 20587
rect 20073 20547 20131 20553
rect 23477 20587 23535 20593
rect 23477 20553 23489 20587
rect 23523 20584 23535 20587
rect 23750 20584 23756 20596
rect 23523 20556 23756 20584
rect 23523 20553 23535 20556
rect 23477 20547 23535 20553
rect 23750 20544 23756 20556
rect 23808 20544 23814 20596
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 13449 20519 13507 20525
rect 13449 20516 13461 20519
rect 12860 20488 13461 20516
rect 12860 20476 12866 20488
rect 13449 20485 13461 20488
rect 13495 20485 13507 20519
rect 17494 20516 17500 20528
rect 17455 20488 17500 20516
rect 13449 20479 13507 20485
rect 17494 20476 17500 20488
rect 17552 20476 17558 20528
rect 23661 20519 23719 20525
rect 23661 20485 23673 20519
rect 23707 20485 23719 20519
rect 23661 20479 23719 20485
rect 3237 20451 3295 20457
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3602 20448 3608 20460
rect 3283 20420 3608 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 5077 20451 5135 20457
rect 5077 20448 5089 20451
rect 4387 20420 5089 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 5077 20417 5089 20420
rect 5123 20448 5135 20451
rect 5166 20448 5172 20460
rect 5123 20420 5172 20448
rect 5123 20417 5135 20420
rect 5077 20411 5135 20417
rect 5166 20408 5172 20420
rect 5224 20448 5230 20460
rect 5534 20448 5540 20460
rect 5224 20420 5540 20448
rect 5224 20408 5230 20420
rect 5534 20408 5540 20420
rect 5592 20408 5598 20460
rect 7098 20448 7104 20460
rect 7059 20420 7104 20448
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 8110 20448 8116 20460
rect 8023 20420 8116 20448
rect 8110 20408 8116 20420
rect 8168 20408 8174 20460
rect 11422 20448 11428 20460
rect 11335 20420 11428 20448
rect 11422 20408 11428 20420
rect 11480 20448 11486 20460
rect 11882 20448 11888 20460
rect 11480 20420 11888 20448
rect 11480 20408 11486 20420
rect 11882 20408 11888 20420
rect 11940 20408 11946 20460
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 13081 20451 13139 20457
rect 13081 20448 13093 20451
rect 12768 20420 13093 20448
rect 12768 20408 12774 20420
rect 13081 20417 13093 20420
rect 13127 20448 13139 20451
rect 13906 20448 13912 20460
rect 13127 20420 13912 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 21545 20451 21603 20457
rect 21545 20417 21557 20451
rect 21591 20448 21603 20451
rect 22557 20451 22615 20457
rect 22557 20448 22569 20451
rect 21591 20420 22569 20448
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 22557 20417 22569 20420
rect 22603 20448 22615 20451
rect 23566 20448 23572 20460
rect 22603 20420 23572 20448
rect 22603 20417 22615 20420
rect 22557 20411 22615 20417
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 3053 20383 3111 20389
rect 3053 20380 3065 20383
rect 1443 20352 2084 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 2056 20256 2084 20352
rect 2424 20352 3065 20380
rect 2314 20272 2320 20324
rect 2372 20312 2378 20324
rect 2424 20321 2452 20352
rect 3053 20349 3065 20352
rect 3099 20349 3111 20383
rect 4798 20380 4804 20392
rect 4711 20352 4804 20380
rect 3053 20343 3111 20349
rect 4798 20340 4804 20352
rect 4856 20380 4862 20392
rect 6181 20383 6239 20389
rect 6181 20380 6193 20383
rect 4856 20352 6193 20380
rect 4856 20340 4862 20352
rect 6181 20349 6193 20352
rect 6227 20349 6239 20383
rect 6638 20380 6644 20392
rect 6599 20352 6644 20380
rect 6181 20343 6239 20349
rect 6638 20340 6644 20352
rect 6696 20340 6702 20392
rect 8386 20389 8392 20392
rect 8380 20380 8392 20389
rect 8299 20352 8392 20380
rect 8380 20343 8392 20352
rect 8444 20380 8450 20392
rect 9122 20380 9128 20392
rect 8444 20352 9128 20380
rect 8386 20340 8392 20343
rect 8444 20340 8450 20352
rect 9122 20340 9128 20352
rect 9180 20340 9186 20392
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 15286 20380 15292 20392
rect 14691 20352 15292 20380
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 15286 20340 15292 20352
rect 15344 20340 15350 20392
rect 18966 20389 18972 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 17604 20352 17877 20380
rect 2409 20315 2467 20321
rect 2409 20312 2421 20315
rect 2372 20284 2421 20312
rect 2372 20272 2378 20284
rect 2409 20281 2421 20284
rect 2455 20281 2467 20315
rect 2409 20275 2467 20281
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20312 4951 20315
rect 11149 20315 11207 20321
rect 11149 20312 11161 20315
rect 4939 20284 5948 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 2038 20244 2044 20256
rect 1999 20216 2044 20244
rect 2038 20204 2044 20216
rect 2096 20204 2102 20256
rect 2958 20244 2964 20256
rect 2871 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20244 3022 20256
rect 3605 20247 3663 20253
rect 3605 20244 3617 20247
rect 3016 20216 3617 20244
rect 3016 20204 3022 20216
rect 3605 20213 3617 20216
rect 3651 20213 3663 20247
rect 4430 20244 4436 20256
rect 4391 20216 4436 20244
rect 3605 20207 3663 20213
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 5534 20244 5540 20256
rect 5495 20216 5540 20244
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 5920 20253 5948 20284
rect 10612 20284 11161 20312
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 5994 20244 6000 20256
rect 5951 20216 6000 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 9493 20247 9551 20253
rect 9493 20244 9505 20247
rect 9456 20216 9505 20244
rect 9456 20204 9462 20216
rect 9493 20213 9505 20216
rect 9539 20213 9551 20247
rect 9493 20207 9551 20213
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 10612 20253 10640 20284
rect 11149 20281 11161 20284
rect 11195 20281 11207 20315
rect 12805 20315 12863 20321
rect 12805 20312 12817 20315
rect 11149 20275 11207 20281
rect 12452 20284 12817 20312
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 9824 20216 10609 20244
rect 9824 20204 9830 20216
rect 10597 20213 10609 20216
rect 10643 20213 10655 20247
rect 11238 20244 11244 20256
rect 11199 20216 11244 20244
rect 10597 20207 10655 20213
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 12161 20247 12219 20253
rect 12161 20244 12173 20247
rect 11388 20216 12173 20244
rect 11388 20204 11394 20216
rect 12161 20213 12173 20216
rect 12207 20244 12219 20247
rect 12452 20244 12480 20284
rect 12805 20281 12817 20284
rect 12851 20312 12863 20315
rect 12986 20312 12992 20324
rect 12851 20284 12992 20312
rect 12851 20281 12863 20284
rect 12805 20275 12863 20281
rect 12986 20272 12992 20284
rect 13044 20272 13050 20324
rect 14918 20321 14924 20324
rect 14912 20312 14924 20321
rect 14831 20284 14924 20312
rect 14912 20275 14924 20284
rect 14976 20312 14982 20324
rect 16206 20312 16212 20324
rect 14976 20284 16212 20312
rect 14918 20272 14924 20275
rect 14976 20272 14982 20284
rect 16206 20272 16212 20284
rect 16264 20272 16270 20324
rect 17604 20256 17632 20352
rect 17865 20349 17877 20352
rect 17911 20349 17923 20383
rect 18693 20383 18751 20389
rect 18693 20380 18705 20383
rect 17865 20343 17923 20349
rect 18340 20352 18705 20380
rect 18340 20256 18368 20352
rect 18693 20349 18705 20352
rect 18739 20349 18751 20383
rect 18960 20380 18972 20389
rect 18927 20352 18972 20380
rect 18693 20343 18751 20349
rect 18960 20343 18972 20352
rect 18966 20340 18972 20343
rect 19024 20340 19030 20392
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21821 20383 21879 20389
rect 21821 20380 21833 20383
rect 20772 20352 21833 20380
rect 20772 20340 20778 20352
rect 21821 20349 21833 20352
rect 21867 20380 21879 20383
rect 23676 20380 23704 20479
rect 24210 20448 24216 20460
rect 24171 20420 24216 20448
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 21867 20352 22232 20380
rect 23676 20352 25237 20380
rect 21867 20349 21879 20352
rect 21821 20343 21879 20349
rect 12894 20244 12900 20256
rect 12207 20216 12480 20244
rect 12855 20216 12900 20244
rect 12207 20213 12219 20216
rect 12161 20207 12219 20213
rect 12894 20204 12900 20216
rect 12952 20204 12958 20256
rect 13906 20244 13912 20256
rect 13867 20216 13912 20244
rect 13906 20204 13912 20216
rect 13964 20204 13970 20256
rect 17221 20247 17279 20253
rect 17221 20213 17233 20247
rect 17267 20244 17279 20247
rect 17586 20244 17592 20256
rect 17267 20216 17592 20244
rect 17267 20213 17279 20216
rect 17221 20207 17279 20213
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 17681 20247 17739 20253
rect 17681 20213 17693 20247
rect 17727 20244 17739 20247
rect 18322 20244 18328 20256
rect 17727 20216 18328 20244
rect 17727 20213 17739 20216
rect 17681 20207 17739 20213
rect 18322 20204 18328 20216
rect 18380 20204 18386 20256
rect 20898 20244 20904 20256
rect 20859 20216 20904 20244
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 20990 20204 20996 20256
rect 21048 20244 21054 20256
rect 21266 20244 21272 20256
rect 21048 20216 21272 20244
rect 21048 20204 21054 20216
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 22002 20244 22008 20256
rect 21963 20216 22008 20244
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22204 20244 22232 20352
rect 25225 20349 25237 20352
rect 25271 20380 25283 20383
rect 25961 20383 26019 20389
rect 25961 20380 25973 20383
rect 25271 20352 25973 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25961 20349 25973 20352
rect 26007 20349 26019 20383
rect 25961 20343 26019 20349
rect 22278 20272 22284 20324
rect 22336 20312 22342 20324
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 22336 20284 22477 20312
rect 22336 20272 22342 20284
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 23750 20272 23756 20324
rect 23808 20312 23814 20324
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23808 20284 24041 20312
rect 23808 20272 23814 20284
rect 24029 20281 24041 20284
rect 24075 20312 24087 20315
rect 25041 20315 25099 20321
rect 25041 20312 25053 20315
rect 24075 20284 25053 20312
rect 24075 20281 24087 20284
rect 24029 20275 24087 20281
rect 25041 20281 25053 20284
rect 25087 20281 25099 20315
rect 25041 20275 25099 20281
rect 25130 20272 25136 20324
rect 25188 20312 25194 20324
rect 25501 20315 25559 20321
rect 25501 20312 25513 20315
rect 25188 20284 25513 20312
rect 25188 20272 25194 20284
rect 25501 20281 25513 20284
rect 25547 20281 25559 20315
rect 25501 20275 25559 20281
rect 22370 20244 22376 20256
rect 22204 20216 22376 20244
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 24118 20244 24124 20256
rect 24079 20216 24124 20244
rect 24118 20204 24124 20216
rect 24176 20244 24182 20256
rect 24673 20247 24731 20253
rect 24673 20244 24685 20247
rect 24176 20216 24685 20244
rect 24176 20204 24182 20216
rect 24673 20213 24685 20216
rect 24719 20213 24731 20247
rect 24673 20207 24731 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1397 20043 1455 20049
rect 1397 20009 1409 20043
rect 1443 20040 1455 20043
rect 2958 20040 2964 20052
rect 1443 20012 2964 20040
rect 1443 20009 1455 20012
rect 1397 20003 1455 20009
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 3513 20043 3571 20049
rect 3513 20009 3525 20043
rect 3559 20040 3571 20043
rect 3602 20040 3608 20052
rect 3559 20012 3608 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 2317 19975 2375 19981
rect 2317 19941 2329 19975
rect 2363 19972 2375 19975
rect 2682 19972 2688 19984
rect 2363 19944 2688 19972
rect 2363 19941 2375 19944
rect 2317 19935 2375 19941
rect 2682 19932 2688 19944
rect 2740 19932 2746 19984
rect 2774 19864 2780 19916
rect 2832 19904 2838 19916
rect 2832 19876 2877 19904
rect 2832 19864 2838 19876
rect 3528 19848 3556 20003
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 8386 20040 8392 20052
rect 8347 20012 8392 20040
rect 8386 20000 8392 20012
rect 8444 20000 8450 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 11238 20040 11244 20052
rect 10183 20012 11244 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11974 20040 11980 20052
rect 11935 20012 11980 20040
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12621 20043 12679 20049
rect 12621 20009 12633 20043
rect 12667 20040 12679 20043
rect 12894 20040 12900 20052
rect 12667 20012 12900 20040
rect 12667 20009 12679 20012
rect 12621 20003 12679 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13630 20040 13636 20052
rect 13587 20012 13636 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 14737 20043 14795 20049
rect 14737 20009 14749 20043
rect 14783 20040 14795 20043
rect 14918 20040 14924 20052
rect 14783 20012 14924 20040
rect 14783 20009 14795 20012
rect 14737 20003 14795 20009
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 16666 20040 16672 20052
rect 16627 20012 16672 20040
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 18966 20000 18972 20052
rect 19024 20040 19030 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19024 20012 19625 20040
rect 19024 20000 19030 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 20717 20043 20775 20049
rect 20717 20009 20729 20043
rect 20763 20040 20775 20043
rect 21358 20040 21364 20052
rect 20763 20012 21364 20040
rect 20763 20009 20775 20012
rect 20717 20003 20775 20009
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 22373 20043 22431 20049
rect 22373 20009 22385 20043
rect 22419 20040 22431 20043
rect 22462 20040 22468 20052
rect 22419 20012 22468 20040
rect 22419 20009 22431 20012
rect 22373 20003 22431 20009
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 23106 20040 23112 20052
rect 23067 20012 23112 20040
rect 23106 20000 23112 20012
rect 23164 20040 23170 20052
rect 23477 20043 23535 20049
rect 23477 20040 23489 20043
rect 23164 20012 23489 20040
rect 23164 20000 23170 20012
rect 23477 20009 23489 20012
rect 23523 20009 23535 20043
rect 23477 20003 23535 20009
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 9030 19972 9036 19984
rect 8168 19944 9036 19972
rect 8168 19932 8174 19944
rect 9030 19932 9036 19944
rect 9088 19932 9094 19984
rect 10505 19975 10563 19981
rect 10505 19941 10517 19975
rect 10551 19972 10563 19975
rect 10864 19975 10922 19981
rect 10864 19972 10876 19975
rect 10551 19944 10876 19972
rect 10551 19941 10563 19944
rect 10505 19935 10563 19941
rect 10864 19941 10876 19944
rect 10910 19972 10922 19975
rect 11422 19972 11428 19984
rect 10910 19944 11428 19972
rect 10910 19941 10922 19944
rect 10864 19935 10922 19941
rect 11422 19932 11428 19944
rect 11480 19932 11486 19984
rect 15556 19975 15614 19981
rect 15556 19941 15568 19975
rect 15602 19972 15614 19975
rect 15654 19972 15660 19984
rect 15602 19944 15660 19972
rect 15602 19941 15614 19944
rect 15556 19935 15614 19941
rect 15654 19932 15660 19944
rect 15712 19932 15718 19984
rect 18500 19975 18558 19981
rect 18500 19941 18512 19975
rect 18546 19972 18558 19975
rect 19150 19972 19156 19984
rect 18546 19944 19156 19972
rect 18546 19941 18558 19944
rect 18500 19935 18558 19941
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 5074 19913 5080 19916
rect 5068 19904 5080 19913
rect 5035 19876 5080 19904
rect 5068 19867 5080 19876
rect 5074 19864 5080 19867
rect 5132 19864 5138 19916
rect 7650 19904 7656 19916
rect 7563 19876 7656 19904
rect 7650 19864 7656 19876
rect 7708 19904 7714 19916
rect 7834 19904 7840 19916
rect 7708 19876 7840 19904
rect 7708 19864 7714 19876
rect 7834 19864 7840 19876
rect 7892 19864 7898 19916
rect 9490 19904 9496 19916
rect 9451 19876 9496 19904
rect 9490 19864 9496 19876
rect 9548 19864 9554 19916
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13262 19904 13268 19916
rect 13044 19876 13268 19904
rect 13044 19864 13050 19876
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 13722 19904 13728 19916
rect 13495 19876 13728 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 13722 19864 13728 19876
rect 13780 19864 13786 19916
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 15378 19904 15384 19916
rect 15335 19876 15384 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15378 19864 15384 19876
rect 15436 19864 15442 19916
rect 17586 19864 17592 19916
rect 17644 19904 17650 19916
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17644 19876 17969 19904
rect 17644 19864 17650 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 18233 19907 18291 19913
rect 18233 19873 18245 19907
rect 18279 19904 18291 19907
rect 18322 19904 18328 19916
rect 18279 19876 18328 19904
rect 18279 19873 18291 19876
rect 18233 19867 18291 19873
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 21266 19913 21272 19916
rect 20993 19907 21051 19913
rect 20993 19904 21005 19907
rect 20864 19876 21005 19904
rect 20864 19864 20870 19876
rect 20993 19873 21005 19876
rect 21039 19873 21051 19907
rect 21260 19904 21272 19913
rect 21227 19876 21272 19904
rect 20993 19867 21051 19873
rect 21260 19867 21272 19876
rect 21266 19864 21272 19867
rect 21324 19864 21330 19916
rect 23492 19904 23520 20003
rect 24302 20000 24308 20052
rect 24360 20040 24366 20052
rect 25133 20043 25191 20049
rect 25133 20040 25145 20043
rect 24360 20012 25145 20040
rect 24360 20000 24366 20012
rect 25133 20009 25145 20012
rect 25179 20009 25191 20043
rect 25133 20003 25191 20009
rect 24020 19975 24078 19981
rect 24020 19941 24032 19975
rect 24066 19972 24078 19975
rect 24210 19972 24216 19984
rect 24066 19944 24216 19972
rect 24066 19941 24078 19944
rect 24020 19935 24078 19941
rect 24210 19932 24216 19944
rect 24268 19972 24274 19984
rect 24854 19972 24860 19984
rect 24268 19944 24860 19972
rect 24268 19932 24274 19944
rect 24854 19932 24860 19944
rect 24912 19932 24918 19984
rect 23753 19907 23811 19913
rect 23753 19904 23765 19907
rect 23492 19876 23765 19904
rect 23753 19873 23765 19876
rect 23799 19873 23811 19907
rect 23753 19867 23811 19873
rect 2866 19836 2872 19848
rect 2827 19808 2872 19836
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19836 3111 19839
rect 3510 19836 3516 19848
rect 3099 19808 3516 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 4246 19796 4252 19848
rect 4304 19836 4310 19848
rect 4801 19839 4859 19845
rect 4801 19836 4813 19839
rect 4304 19808 4813 19836
rect 4304 19796 4310 19808
rect 4801 19805 4813 19808
rect 4847 19805 4859 19839
rect 7742 19836 7748 19848
rect 7703 19808 7748 19836
rect 4801 19799 4859 19805
rect 7742 19796 7748 19808
rect 7800 19796 7806 19848
rect 7926 19836 7932 19848
rect 7887 19808 7932 19836
rect 7926 19796 7932 19808
rect 7984 19796 7990 19848
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 9030 19836 9036 19848
rect 8803 19808 9036 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 10134 19836 10140 19848
rect 9324 19808 10140 19836
rect 1949 19771 2007 19777
rect 1949 19737 1961 19771
rect 1995 19768 2007 19771
rect 2409 19771 2467 19777
rect 2409 19768 2421 19771
rect 1995 19740 2421 19768
rect 1995 19737 2007 19740
rect 1949 19731 2007 19737
rect 2409 19737 2421 19740
rect 2455 19768 2467 19771
rect 2590 19768 2596 19780
rect 2455 19740 2596 19768
rect 2455 19737 2467 19740
rect 2409 19731 2467 19737
rect 2590 19728 2596 19740
rect 2648 19728 2654 19780
rect 3602 19660 3608 19712
rect 3660 19700 3666 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3660 19672 3801 19700
rect 3660 19660 3666 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 4338 19700 4344 19712
rect 4299 19672 4344 19700
rect 3789 19663 3847 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 4706 19700 4712 19712
rect 4667 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 6181 19703 6239 19709
rect 6181 19700 6193 19703
rect 5500 19672 6193 19700
rect 5500 19660 5506 19672
rect 6181 19669 6193 19672
rect 6227 19700 6239 19703
rect 6822 19700 6828 19712
rect 6227 19672 6828 19700
rect 6227 19669 6239 19672
rect 6181 19663 6239 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7190 19660 7196 19712
rect 7248 19700 7254 19712
rect 7285 19703 7343 19709
rect 7285 19700 7297 19703
rect 7248 19672 7297 19700
rect 7248 19660 7254 19672
rect 7285 19669 7297 19672
rect 7331 19669 7343 19703
rect 7285 19663 7343 19669
rect 8570 19660 8576 19712
rect 8628 19700 8634 19712
rect 9324 19709 9352 19808
rect 10134 19796 10140 19808
rect 10192 19836 10198 19848
rect 10597 19839 10655 19845
rect 10597 19836 10609 19839
rect 10192 19808 10609 19836
rect 10192 19796 10198 19808
rect 10597 19805 10609 19808
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 12989 19771 13047 19777
rect 12989 19737 13001 19771
rect 13035 19768 13047 19771
rect 13262 19768 13268 19780
rect 13035 19740 13268 19768
rect 13035 19737 13047 19740
rect 12989 19731 13047 19737
rect 13262 19728 13268 19740
rect 13320 19768 13326 19780
rect 13648 19768 13676 19799
rect 13320 19740 13676 19768
rect 13320 19728 13326 19740
rect 14550 19728 14556 19780
rect 14608 19768 14614 19780
rect 15013 19771 15071 19777
rect 15013 19768 15025 19771
rect 14608 19740 15025 19768
rect 14608 19728 14614 19740
rect 15013 19737 15025 19740
rect 15059 19737 15071 19771
rect 15013 19731 15071 19737
rect 17313 19771 17371 19777
rect 17313 19737 17325 19771
rect 17359 19768 17371 19771
rect 17773 19771 17831 19777
rect 17773 19768 17785 19771
rect 17359 19740 17785 19768
rect 17359 19737 17371 19740
rect 17313 19731 17371 19737
rect 17773 19737 17785 19740
rect 17819 19768 17831 19771
rect 17862 19768 17868 19780
rect 17819 19740 17868 19768
rect 17819 19737 17831 19740
rect 17773 19731 17831 19737
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 8628 19672 9321 19700
rect 8628 19660 8634 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 13078 19700 13084 19712
rect 13039 19672 13084 19700
rect 9309 19663 9367 19669
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 14185 19703 14243 19709
rect 14185 19669 14197 19703
rect 14231 19700 14243 19703
rect 14458 19700 14464 19712
rect 14231 19672 14464 19700
rect 14231 19669 14243 19672
rect 14185 19663 14243 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 17586 19700 17592 19712
rect 17547 19672 17592 19700
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2130 19456 2136 19508
rect 2188 19496 2194 19508
rect 2590 19496 2596 19508
rect 2188 19468 2596 19496
rect 2188 19456 2194 19468
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 3510 19456 3516 19508
rect 3568 19496 3574 19508
rect 3697 19499 3755 19505
rect 3697 19496 3709 19499
rect 3568 19468 3709 19496
rect 3568 19456 3574 19468
rect 3697 19465 3709 19468
rect 3743 19465 3755 19499
rect 3697 19459 3755 19465
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 5629 19499 5687 19505
rect 5629 19496 5641 19499
rect 5592 19468 5641 19496
rect 5592 19456 5598 19468
rect 5629 19465 5641 19468
rect 5675 19465 5687 19499
rect 5629 19459 5687 19465
rect 5994 19456 6000 19508
rect 6052 19496 6058 19508
rect 6825 19499 6883 19505
rect 6825 19496 6837 19499
rect 6052 19468 6837 19496
rect 6052 19456 6058 19468
rect 6825 19465 6837 19468
rect 6871 19465 6883 19499
rect 6825 19459 6883 19465
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11422 19496 11428 19508
rect 11379 19468 11428 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 11422 19456 11428 19468
rect 11480 19456 11486 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 13541 19499 13599 19505
rect 12492 19468 12537 19496
rect 12492 19456 12498 19468
rect 13541 19465 13553 19499
rect 13587 19496 13599 19499
rect 13630 19496 13636 19508
rect 13587 19468 13636 19496
rect 13587 19465 13599 19468
rect 13541 19459 13599 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 16850 19496 16856 19508
rect 15712 19468 16856 19496
rect 15712 19456 15718 19468
rect 16850 19456 16856 19468
rect 16908 19496 16914 19508
rect 16945 19499 17003 19505
rect 16945 19496 16957 19499
rect 16908 19468 16957 19496
rect 16908 19456 16914 19468
rect 16945 19465 16957 19468
rect 16991 19465 17003 19499
rect 19150 19496 19156 19508
rect 19111 19468 19156 19496
rect 16945 19459 17003 19465
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 19334 19456 19340 19508
rect 19392 19496 19398 19508
rect 23750 19496 23756 19508
rect 19392 19468 23612 19496
rect 23711 19468 23756 19496
rect 19392 19456 19398 19468
rect 2501 19431 2559 19437
rect 2501 19397 2513 19431
rect 2547 19428 2559 19431
rect 2866 19428 2872 19440
rect 2547 19400 2872 19428
rect 2547 19397 2559 19400
rect 2501 19391 2559 19397
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 6641 19431 6699 19437
rect 6641 19397 6653 19431
rect 6687 19428 6699 19431
rect 7926 19428 7932 19440
rect 6687 19400 7932 19428
rect 6687 19397 6699 19400
rect 6641 19391 6699 19397
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3510 19360 3516 19372
rect 3375 19332 3516 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 6656 19360 6684 19391
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 10229 19431 10287 19437
rect 10229 19397 10241 19431
rect 10275 19428 10287 19431
rect 10778 19428 10784 19440
rect 10275 19400 10784 19428
rect 10275 19397 10287 19400
rect 10229 19391 10287 19397
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 12618 19388 12624 19440
rect 12676 19428 12682 19440
rect 15746 19428 15752 19440
rect 12676 19400 15752 19428
rect 12676 19388 12682 19400
rect 15746 19388 15752 19400
rect 15804 19388 15810 19440
rect 23584 19428 23612 19468
rect 23750 19456 23756 19468
rect 23808 19456 23814 19508
rect 25774 19428 25780 19440
rect 23584 19400 25780 19428
rect 25774 19388 25780 19400
rect 25832 19388 25838 19440
rect 6196 19332 6684 19360
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 4246 19292 4252 19304
rect 4207 19264 4252 19292
rect 4246 19252 4252 19264
rect 4304 19252 4310 19304
rect 5074 19292 5080 19304
rect 4356 19264 5080 19292
rect 1670 19224 1676 19236
rect 1631 19196 1676 19224
rect 1670 19184 1676 19196
rect 1728 19184 1734 19236
rect 3145 19227 3203 19233
rect 3145 19193 3157 19227
rect 3191 19224 3203 19227
rect 3878 19224 3884 19236
rect 3191 19196 3884 19224
rect 3191 19193 3203 19196
rect 3145 19187 3203 19193
rect 3878 19184 3884 19196
rect 3936 19184 3942 19236
rect 4154 19224 4160 19236
rect 4067 19196 4160 19224
rect 4154 19184 4160 19196
rect 4212 19224 4218 19236
rect 4356 19224 4384 19264
rect 5074 19252 5080 19264
rect 5132 19292 5138 19304
rect 6196 19292 6224 19332
rect 6822 19320 6828 19372
rect 6880 19360 6886 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 6880 19332 7389 19360
rect 6880 19320 6886 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 9214 19360 9220 19372
rect 9175 19332 9220 19360
rect 7377 19323 7435 19329
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 9769 19363 9827 19369
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 10873 19363 10931 19369
rect 10873 19360 10885 19363
rect 9815 19332 10885 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 10873 19329 10885 19332
rect 10919 19360 10931 19363
rect 11146 19360 11152 19372
rect 10919 19332 11152 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12710 19360 12716 19372
rect 11931 19332 12716 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12710 19320 12716 19332
rect 12768 19360 12774 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12768 19332 13001 19360
rect 12768 19320 12774 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13998 19320 14004 19372
rect 14056 19360 14062 19372
rect 14553 19363 14611 19369
rect 14553 19360 14565 19363
rect 14056 19332 14565 19360
rect 14056 19320 14062 19332
rect 14553 19329 14565 19332
rect 14599 19329 14611 19363
rect 14553 19323 14611 19329
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 16577 19363 16635 19369
rect 16577 19360 16589 19363
rect 16264 19332 16589 19360
rect 16264 19320 16270 19332
rect 16577 19329 16589 19332
rect 16623 19360 16635 19363
rect 16850 19360 16856 19372
rect 16623 19332 16856 19360
rect 16623 19329 16635 19332
rect 16577 19323 16635 19329
rect 16850 19320 16856 19332
rect 16908 19320 16914 19372
rect 18598 19360 18604 19372
rect 18559 19332 18604 19360
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 20806 19360 20812 19372
rect 20767 19332 20812 19360
rect 20806 19320 20812 19332
rect 20864 19320 20870 19372
rect 24302 19360 24308 19372
rect 24263 19332 24308 19360
rect 24302 19320 24308 19332
rect 24360 19360 24366 19372
rect 24765 19363 24823 19369
rect 24765 19360 24777 19363
rect 24360 19332 24777 19360
rect 24360 19320 24366 19332
rect 24765 19329 24777 19332
rect 24811 19329 24823 19363
rect 24765 19323 24823 19329
rect 5132 19264 6224 19292
rect 6273 19295 6331 19301
rect 5132 19252 5138 19264
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 7282 19292 7288 19304
rect 6319 19264 7288 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 9858 19252 9864 19304
rect 9916 19292 9922 19304
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 9916 19264 10609 19292
rect 9916 19252 9922 19264
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 12897 19295 12955 19301
rect 12897 19292 12909 19295
rect 10597 19255 10655 19261
rect 12176 19264 12909 19292
rect 4522 19233 4528 19236
rect 4516 19224 4528 19233
rect 4212 19196 4384 19224
rect 4483 19196 4528 19224
rect 4212 19184 4218 19196
rect 4516 19187 4528 19196
rect 4522 19184 4528 19187
rect 4580 19184 4586 19236
rect 8573 19227 8631 19233
rect 8573 19193 8585 19227
rect 8619 19224 8631 19227
rect 8938 19224 8944 19236
rect 8619 19196 8944 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 8938 19184 8944 19196
rect 8996 19224 9002 19236
rect 9125 19227 9183 19233
rect 9125 19224 9137 19227
rect 8996 19196 9137 19224
rect 8996 19184 9002 19196
rect 9125 19193 9137 19196
rect 9171 19193 9183 19227
rect 10042 19224 10048 19236
rect 10003 19196 10048 19224
rect 9125 19187 9183 19193
rect 10042 19184 10048 19196
rect 10100 19184 10106 19236
rect 2685 19159 2743 19165
rect 2685 19125 2697 19159
rect 2731 19156 2743 19159
rect 2866 19156 2872 19168
rect 2731 19128 2872 19156
rect 2731 19125 2743 19128
rect 2685 19119 2743 19125
rect 2866 19116 2872 19128
rect 2924 19116 2930 19168
rect 3053 19159 3111 19165
rect 3053 19125 3065 19159
rect 3099 19156 3111 19159
rect 3602 19156 3608 19168
rect 3099 19128 3608 19156
rect 3099 19125 3111 19128
rect 3053 19119 3111 19125
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19116 7254 19168
rect 7834 19156 7840 19168
rect 7795 19128 7840 19156
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 8662 19156 8668 19168
rect 8623 19128 8668 19156
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 9030 19156 9036 19168
rect 8991 19128 9036 19156
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 10060 19156 10088 19184
rect 10689 19159 10747 19165
rect 10689 19156 10701 19159
rect 10060 19128 10701 19156
rect 10689 19125 10701 19128
rect 10735 19125 10747 19159
rect 10689 19119 10747 19125
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12176 19165 12204 19264
rect 12897 19261 12909 19264
rect 12943 19292 12955 19295
rect 13354 19292 13360 19304
rect 12943 19264 13360 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 13354 19252 13360 19264
rect 13412 19252 13418 19304
rect 15013 19295 15071 19301
rect 15013 19292 15025 19295
rect 13832 19264 15025 19292
rect 13832 19168 13860 19264
rect 15013 19261 15025 19264
rect 15059 19261 15071 19295
rect 15013 19255 15071 19261
rect 15473 19295 15531 19301
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 16022 19292 16028 19304
rect 15519 19264 16028 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 14366 19224 14372 19236
rect 14327 19196 14372 19224
rect 14366 19184 14372 19196
rect 14424 19184 14430 19236
rect 15028 19224 15056 19255
rect 16022 19252 16028 19264
rect 16080 19252 16086 19304
rect 18414 19292 18420 19304
rect 17420 19264 18420 19292
rect 15933 19227 15991 19233
rect 15933 19224 15945 19227
rect 15028 19196 15945 19224
rect 15933 19193 15945 19196
rect 15979 19193 15991 19227
rect 15933 19187 15991 19193
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 12032 19128 12173 19156
rect 12032 19116 12038 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 12161 19119 12219 19125
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12492 19128 12817 19156
rect 12492 19116 12498 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 12805 19119 12863 19125
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14001 19159 14059 19165
rect 14001 19125 14013 19159
rect 14047 19156 14059 19159
rect 14090 19156 14096 19168
rect 14047 19128 14096 19156
rect 14047 19125 14059 19128
rect 14001 19119 14059 19125
rect 14090 19116 14096 19128
rect 14148 19116 14154 19168
rect 14458 19156 14464 19168
rect 14419 19128 14464 19156
rect 14458 19116 14464 19128
rect 14516 19116 14522 19168
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 14792 19128 15577 19156
rect 14792 19116 14798 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 17126 19116 17132 19168
rect 17184 19156 17190 19168
rect 17420 19165 17448 19264
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19536 19264 19625 19292
rect 18506 19224 18512 19236
rect 17788 19196 18512 19224
rect 17788 19168 17816 19196
rect 18506 19184 18512 19196
rect 18564 19184 18570 19236
rect 19536 19168 19564 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 24780 19292 24808 19323
rect 25133 19295 25191 19301
rect 25133 19292 25145 19295
rect 24780 19264 25145 19292
rect 19613 19255 19671 19261
rect 25133 19261 25145 19264
rect 25179 19261 25191 19295
rect 25314 19292 25320 19304
rect 25275 19264 25320 19292
rect 25133 19255 25191 19261
rect 25314 19252 25320 19264
rect 25372 19292 25378 19304
rect 26053 19295 26111 19301
rect 26053 19292 26065 19295
rect 25372 19264 26065 19292
rect 25372 19252 25378 19264
rect 26053 19261 26065 19264
rect 26099 19261 26111 19295
rect 26053 19255 26111 19261
rect 19702 19184 19708 19236
rect 19760 19184 19766 19236
rect 20349 19227 20407 19233
rect 20349 19193 20361 19227
rect 20395 19224 20407 19227
rect 21054 19227 21112 19233
rect 21054 19224 21066 19227
rect 20395 19196 21066 19224
rect 20395 19193 20407 19196
rect 20349 19187 20407 19193
rect 21054 19193 21066 19196
rect 21100 19224 21112 19227
rect 21542 19224 21548 19236
rect 21100 19196 21548 19224
rect 21100 19193 21112 19196
rect 21054 19187 21112 19193
rect 21542 19184 21548 19196
rect 21600 19184 21606 19236
rect 22462 19184 22468 19236
rect 22520 19224 22526 19236
rect 23109 19227 23167 19233
rect 23109 19224 23121 19227
rect 22520 19196 23121 19224
rect 22520 19184 22526 19196
rect 23109 19193 23121 19196
rect 23155 19224 23167 19227
rect 24121 19227 24179 19233
rect 24121 19224 24133 19227
rect 23155 19196 24133 19224
rect 23155 19193 23167 19196
rect 23109 19187 23167 19193
rect 24121 19193 24133 19196
rect 24167 19193 24179 19227
rect 25590 19224 25596 19236
rect 25551 19196 25596 19224
rect 24121 19187 24179 19193
rect 25590 19184 25596 19196
rect 25648 19184 25654 19236
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 17184 19128 17417 19156
rect 17184 19116 17190 19128
rect 17405 19125 17417 19128
rect 17451 19125 17463 19159
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17405 19119 17463 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18046 19156 18052 19168
rect 18007 19128 18052 19156
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 19518 19156 19524 19168
rect 19479 19128 19524 19156
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 19720 19156 19748 19184
rect 19797 19159 19855 19165
rect 19797 19156 19809 19159
rect 19720 19128 19809 19156
rect 19797 19125 19809 19128
rect 19843 19125 19855 19159
rect 19797 19119 19855 19125
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 21266 19156 21272 19168
rect 20763 19128 21272 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 21266 19116 21272 19128
rect 21324 19156 21330 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21324 19128 22201 19156
rect 21324 19116 21330 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 22189 19119 22247 19125
rect 23477 19159 23535 19165
rect 23477 19125 23489 19159
rect 23523 19156 23535 19159
rect 24213 19159 24271 19165
rect 24213 19156 24225 19159
rect 23523 19128 24225 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 24213 19125 24225 19128
rect 24259 19156 24271 19159
rect 25774 19156 25780 19168
rect 24259 19128 25780 19156
rect 24259 19125 24271 19128
rect 24213 19119 24271 19125
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 2498 18952 2504 18964
rect 2459 18924 2504 18952
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 3053 18955 3111 18961
rect 3053 18952 3065 18955
rect 2832 18924 3065 18952
rect 2832 18912 2838 18924
rect 3053 18921 3065 18924
rect 3099 18952 3111 18955
rect 3326 18952 3332 18964
rect 3099 18924 3332 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 3326 18912 3332 18924
rect 3384 18912 3390 18964
rect 4706 18912 4712 18964
rect 4764 18952 4770 18964
rect 5074 18952 5080 18964
rect 4764 18924 5080 18952
rect 4764 18912 4770 18924
rect 5074 18912 5080 18924
rect 5132 18952 5138 18964
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 5132 18924 5273 18952
rect 5132 18912 5138 18924
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 5261 18915 5319 18921
rect 6270 18912 6276 18964
rect 6328 18952 6334 18964
rect 6457 18955 6515 18961
rect 6457 18952 6469 18955
rect 6328 18924 6469 18952
rect 6328 18912 6334 18924
rect 6457 18921 6469 18924
rect 6503 18921 6515 18955
rect 6457 18915 6515 18921
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 6825 18955 6883 18961
rect 6825 18952 6837 18955
rect 6788 18924 6837 18952
rect 6788 18912 6794 18924
rect 6825 18921 6837 18924
rect 6871 18921 6883 18955
rect 6825 18915 6883 18921
rect 7561 18955 7619 18961
rect 7561 18921 7573 18955
rect 7607 18952 7619 18955
rect 7742 18952 7748 18964
rect 7607 18924 7748 18952
rect 7607 18921 7619 18924
rect 7561 18915 7619 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 9125 18955 9183 18961
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9214 18952 9220 18964
rect 9171 18924 9220 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 10229 18955 10287 18961
rect 10229 18952 10241 18955
rect 9916 18924 10241 18952
rect 9916 18912 9922 18924
rect 10229 18921 10241 18924
rect 10275 18921 10287 18955
rect 10229 18915 10287 18921
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13078 18952 13084 18964
rect 12860 18924 13084 18952
rect 12860 18912 12866 18924
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 14366 18952 14372 18964
rect 14327 18924 14372 18952
rect 14366 18912 14372 18924
rect 14424 18912 14430 18964
rect 15010 18952 15016 18964
rect 14971 18924 15016 18952
rect 15010 18912 15016 18924
rect 15068 18952 15074 18964
rect 15749 18955 15807 18961
rect 15749 18952 15761 18955
rect 15068 18924 15761 18952
rect 15068 18912 15074 18924
rect 15749 18921 15761 18924
rect 15795 18921 15807 18955
rect 15749 18915 15807 18921
rect 18138 18912 18144 18964
rect 18196 18952 18202 18964
rect 18233 18955 18291 18961
rect 18233 18952 18245 18955
rect 18196 18924 18245 18952
rect 18196 18912 18202 18924
rect 18233 18921 18245 18924
rect 18279 18921 18291 18955
rect 18233 18915 18291 18921
rect 20806 18912 20812 18964
rect 20864 18952 20870 18964
rect 21913 18955 21971 18961
rect 21913 18952 21925 18955
rect 20864 18924 21925 18952
rect 20864 18912 20870 18924
rect 21913 18921 21925 18924
rect 21959 18952 21971 18955
rect 22189 18955 22247 18961
rect 22189 18952 22201 18955
rect 21959 18924 22201 18952
rect 21959 18921 21971 18924
rect 21913 18915 21971 18921
rect 22189 18921 22201 18924
rect 22235 18921 22247 18955
rect 22462 18952 22468 18964
rect 22423 18924 22468 18952
rect 22189 18915 22247 18921
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 23477 18955 23535 18961
rect 23477 18921 23489 18955
rect 23523 18952 23535 18955
rect 24118 18952 24124 18964
rect 23523 18924 24124 18952
rect 23523 18921 23535 18924
rect 23477 18915 23535 18921
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 25225 18955 25283 18961
rect 25225 18952 25237 18955
rect 24912 18924 25237 18952
rect 24912 18912 24918 18924
rect 25225 18921 25237 18924
rect 25271 18921 25283 18955
rect 25225 18915 25283 18921
rect 4338 18844 4344 18896
rect 4396 18884 4402 18896
rect 5166 18884 5172 18896
rect 4396 18856 5172 18884
rect 4396 18844 4402 18856
rect 5166 18844 5172 18856
rect 5224 18844 5230 18896
rect 5997 18887 6055 18893
rect 5997 18853 6009 18887
rect 6043 18884 6055 18887
rect 7190 18884 7196 18896
rect 6043 18856 7196 18884
rect 6043 18853 6055 18856
rect 5997 18847 6055 18853
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 8018 18844 8024 18896
rect 8076 18884 8082 18896
rect 8481 18887 8539 18893
rect 8481 18884 8493 18887
rect 8076 18856 8493 18884
rect 8076 18844 8082 18856
rect 8481 18853 8493 18856
rect 8527 18884 8539 18887
rect 8754 18884 8760 18896
rect 8527 18856 8760 18884
rect 8527 18853 8539 18856
rect 8481 18847 8539 18853
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 10502 18844 10508 18896
rect 10560 18884 10566 18896
rect 10680 18887 10738 18893
rect 10680 18884 10692 18887
rect 10560 18856 10692 18884
rect 10560 18844 10566 18856
rect 10680 18853 10692 18856
rect 10726 18884 10738 18887
rect 10962 18884 10968 18896
rect 10726 18856 10968 18884
rect 10726 18853 10738 18856
rect 10680 18847 10738 18853
rect 10962 18844 10968 18856
rect 11020 18844 11026 18896
rect 15654 18884 15660 18896
rect 15615 18856 15660 18884
rect 15654 18844 15660 18856
rect 15712 18884 15718 18896
rect 16301 18887 16359 18893
rect 16301 18884 16313 18887
rect 15712 18856 16313 18884
rect 15712 18844 15718 18856
rect 16301 18853 16313 18856
rect 16347 18853 16359 18887
rect 16301 18847 16359 18853
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 19242 18884 19248 18896
rect 18012 18856 19248 18884
rect 18012 18844 18018 18856
rect 19242 18844 19248 18856
rect 19300 18844 19306 18896
rect 23566 18844 23572 18896
rect 23624 18884 23630 18896
rect 23750 18884 23756 18896
rect 23624 18856 23756 18884
rect 23624 18844 23630 18856
rect 23750 18844 23756 18856
rect 23808 18884 23814 18896
rect 24489 18887 24547 18893
rect 24489 18884 24501 18887
rect 23808 18856 24501 18884
rect 23808 18844 23814 18856
rect 24489 18853 24501 18856
rect 24535 18853 24547 18887
rect 24489 18847 24547 18853
rect 1762 18776 1768 18828
rect 1820 18816 1826 18828
rect 2409 18819 2467 18825
rect 2409 18816 2421 18819
rect 1820 18788 2421 18816
rect 1820 18776 1826 18788
rect 2409 18785 2421 18788
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 6365 18819 6423 18825
rect 6365 18785 6377 18819
rect 6411 18816 6423 18819
rect 6730 18816 6736 18828
rect 6411 18788 6736 18816
rect 6411 18785 6423 18788
rect 6365 18779 6423 18785
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 8110 18776 8116 18828
rect 8168 18816 8174 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 8168 18788 8401 18816
rect 8168 18776 8174 18788
rect 8389 18785 8401 18788
rect 8435 18816 8447 18819
rect 11790 18816 11796 18828
rect 8435 18788 11796 18816
rect 8435 18785 8447 18788
rect 8389 18779 8447 18785
rect 11790 18776 11796 18788
rect 11848 18776 11854 18828
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 12492 18788 13277 18816
rect 12492 18776 12498 18788
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 17494 18776 17500 18828
rect 17552 18816 17558 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 17552 18788 18153 18816
rect 17552 18776 17558 18788
rect 18141 18785 18153 18788
rect 18187 18816 18199 18819
rect 19150 18816 19156 18828
rect 18187 18788 19156 18816
rect 18187 18785 18199 18788
rect 18141 18779 18199 18785
rect 19150 18776 19156 18788
rect 19208 18776 19214 18828
rect 19334 18816 19340 18828
rect 19295 18788 19340 18816
rect 19334 18776 19340 18788
rect 19392 18816 19398 18828
rect 20073 18819 20131 18825
rect 20073 18816 20085 18819
rect 19392 18788 20085 18816
rect 19392 18776 19398 18788
rect 20073 18785 20085 18788
rect 20119 18785 20131 18819
rect 20714 18816 20720 18828
rect 20627 18788 20720 18816
rect 20073 18779 20131 18785
rect 20714 18776 20720 18788
rect 20772 18816 20778 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 20772 18788 21281 18816
rect 20772 18776 20778 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18816 21419 18819
rect 21542 18816 21548 18828
rect 21407 18788 21548 18816
rect 21407 18785 21419 18788
rect 21361 18779 21419 18785
rect 21542 18776 21548 18788
rect 21600 18776 21606 18828
rect 23845 18819 23903 18825
rect 23845 18785 23857 18819
rect 23891 18816 23903 18819
rect 24118 18816 24124 18828
rect 23891 18788 24124 18816
rect 23891 18785 23903 18788
rect 23845 18779 23903 18785
rect 24118 18776 24124 18788
rect 24176 18776 24182 18828
rect 25041 18819 25099 18825
rect 25041 18785 25053 18819
rect 25087 18816 25099 18819
rect 25130 18816 25136 18828
rect 25087 18788 25136 18816
rect 25087 18785 25099 18788
rect 25041 18779 25099 18785
rect 25130 18776 25136 18788
rect 25188 18776 25194 18828
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18748 2743 18751
rect 4341 18751 4399 18757
rect 2731 18720 3556 18748
rect 2731 18717 2743 18720
rect 2685 18711 2743 18717
rect 1946 18680 1952 18692
rect 1907 18652 1952 18680
rect 1946 18640 1952 18652
rect 2004 18640 2010 18692
rect 3528 18624 3556 18720
rect 4341 18717 4353 18751
rect 4387 18748 4399 18751
rect 4522 18748 4528 18760
rect 4387 18720 4528 18748
rect 4387 18717 4399 18720
rect 4341 18711 4399 18717
rect 4522 18708 4528 18720
rect 4580 18748 4586 18760
rect 4709 18751 4767 18757
rect 4709 18748 4721 18751
rect 4580 18720 4721 18748
rect 4580 18708 4586 18720
rect 4709 18717 4721 18720
rect 4755 18748 4767 18751
rect 5442 18748 5448 18760
rect 4755 18720 5448 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 5442 18708 5448 18720
rect 5500 18708 5506 18760
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6840 18720 6929 18748
rect 6840 18692 6868 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 8294 18748 8300 18760
rect 7147 18720 8300 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 4798 18680 4804 18692
rect 4759 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 6822 18640 6828 18692
rect 6880 18640 6886 18692
rect 2038 18612 2044 18624
rect 1999 18584 2044 18612
rect 2038 18572 2044 18584
rect 2096 18572 2102 18624
rect 3510 18612 3516 18624
rect 3471 18584 3516 18612
rect 3510 18572 3516 18584
rect 3568 18572 3574 18624
rect 3878 18612 3884 18624
rect 3839 18584 3884 18612
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 7116 18612 7144 18711
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 10410 18748 10416 18760
rect 8573 18711 8631 18717
rect 9324 18720 10416 18748
rect 7929 18683 7987 18689
rect 7929 18649 7941 18683
rect 7975 18680 7987 18683
rect 8588 18680 8616 18711
rect 8662 18680 8668 18692
rect 7975 18652 8668 18680
rect 7975 18649 7987 18652
rect 7929 18643 7987 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 6604 18584 7144 18612
rect 8021 18615 8079 18621
rect 6604 18572 6610 18584
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 8294 18612 8300 18624
rect 8067 18584 8300 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9324 18612 9352 18720
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 12584 18720 13369 18748
rect 12584 18708 12590 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 12400 18652 13032 18680
rect 12400 18640 12406 18652
rect 9490 18612 9496 18624
rect 8628 18584 9352 18612
rect 9451 18584 9496 18612
rect 8628 18572 8634 18584
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 9858 18612 9864 18624
rect 9819 18584 9864 18612
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11793 18615 11851 18621
rect 11793 18612 11805 18615
rect 11112 18584 11805 18612
rect 11112 18572 11118 18584
rect 11793 18581 11805 18584
rect 11839 18581 11851 18615
rect 11793 18575 11851 18581
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12492 18584 12537 18612
rect 12492 18572 12498 18584
rect 12710 18572 12716 18624
rect 12768 18612 12774 18624
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 12768 18584 12909 18612
rect 12768 18572 12774 18584
rect 12897 18581 12909 18584
rect 12943 18581 12955 18615
rect 13004 18612 13032 18652
rect 13262 18640 13268 18692
rect 13320 18680 13326 18692
rect 13464 18680 13492 18711
rect 14734 18708 14740 18760
rect 14792 18748 14798 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 14792 18720 15853 18748
rect 14792 18708 14798 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18748 18475 18751
rect 18598 18748 18604 18760
rect 18463 18720 18604 18748
rect 18463 18717 18475 18720
rect 18417 18711 18475 18717
rect 18598 18708 18604 18720
rect 18656 18748 18662 18760
rect 18656 18720 18920 18748
rect 18656 18708 18662 18720
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 13320 18652 13492 18680
rect 13556 18652 16773 18680
rect 13320 18640 13326 18652
rect 13556 18612 13584 18652
rect 16761 18649 16773 18652
rect 16807 18680 16819 18683
rect 17129 18683 17187 18689
rect 17129 18680 17141 18683
rect 16807 18652 17141 18680
rect 16807 18649 16819 18652
rect 16761 18643 16819 18649
rect 17129 18649 17141 18652
rect 17175 18680 17187 18683
rect 18506 18680 18512 18692
rect 17175 18652 18512 18680
rect 17175 18649 17187 18652
rect 17129 18643 17187 18649
rect 18506 18640 18512 18652
rect 18564 18640 18570 18692
rect 13998 18612 14004 18624
rect 13004 18584 13584 18612
rect 13959 18584 14004 18612
rect 12897 18575 12955 18581
rect 13998 18572 14004 18584
rect 14056 18572 14062 18624
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 15289 18615 15347 18621
rect 15289 18612 15301 18615
rect 14148 18584 15301 18612
rect 14148 18572 14154 18584
rect 15289 18581 15301 18584
rect 15335 18581 15347 18615
rect 15289 18575 15347 18581
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 17727 18584 17785 18612
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 17773 18581 17785 18584
rect 17819 18612 17831 18615
rect 18414 18612 18420 18624
rect 17819 18584 18420 18612
rect 17819 18581 17831 18584
rect 17773 18575 17831 18581
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18892 18621 18920 18720
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19484 18720 19533 18748
rect 19484 18708 19490 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 21450 18748 21456 18760
rect 21411 18720 21456 18748
rect 19521 18711 19579 18717
rect 21450 18708 21456 18720
rect 21508 18708 21514 18760
rect 23106 18708 23112 18760
rect 23164 18748 23170 18760
rect 23937 18751 23995 18757
rect 23937 18748 23949 18751
rect 23164 18720 23949 18748
rect 23164 18708 23170 18720
rect 23937 18717 23949 18720
rect 23983 18717 23995 18751
rect 23937 18711 23995 18717
rect 24029 18751 24087 18757
rect 24029 18717 24041 18751
rect 24075 18748 24087 18751
rect 24302 18748 24308 18760
rect 24075 18720 24308 18748
rect 24075 18717 24087 18720
rect 24029 18711 24087 18717
rect 23566 18640 23572 18692
rect 23624 18680 23630 18692
rect 24044 18680 24072 18711
rect 24302 18708 24308 18720
rect 24360 18708 24366 18760
rect 23624 18652 24072 18680
rect 23624 18640 23630 18652
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 18966 18612 18972 18624
rect 18923 18584 18972 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 19242 18612 19248 18624
rect 19203 18584 19248 18612
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 20901 18615 20959 18621
rect 20901 18581 20913 18615
rect 20947 18612 20959 18615
rect 21358 18612 21364 18624
rect 20947 18584 21364 18612
rect 20947 18581 20959 18584
rect 20901 18575 20959 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 22189 18615 22247 18621
rect 22189 18581 22201 18615
rect 22235 18612 22247 18615
rect 22373 18615 22431 18621
rect 22373 18612 22385 18615
rect 22235 18584 22385 18612
rect 22235 18581 22247 18584
rect 22189 18575 22247 18581
rect 22373 18581 22385 18584
rect 22419 18612 22431 18615
rect 23290 18612 23296 18624
rect 22419 18584 23296 18612
rect 22419 18581 22431 18584
rect 22373 18575 22431 18581
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24210 18612 24216 18624
rect 23900 18584 24216 18612
rect 23900 18572 23906 18584
rect 24210 18572 24216 18584
rect 24268 18572 24274 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1762 18408 1768 18420
rect 1723 18380 1768 18408
rect 1762 18368 1768 18380
rect 1820 18368 1826 18420
rect 2133 18411 2191 18417
rect 2133 18377 2145 18411
rect 2179 18408 2191 18411
rect 2498 18408 2504 18420
rect 2179 18380 2504 18408
rect 2179 18377 2191 18380
rect 2133 18371 2191 18377
rect 2498 18368 2504 18380
rect 2556 18368 2562 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4249 18411 4307 18417
rect 4249 18408 4261 18411
rect 4212 18380 4261 18408
rect 4212 18368 4218 18380
rect 4249 18377 4261 18380
rect 4295 18377 4307 18411
rect 5166 18408 5172 18420
rect 5127 18380 5172 18408
rect 4249 18371 4307 18377
rect 4264 18272 4292 18371
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 6546 18408 6552 18420
rect 6507 18380 6552 18408
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 8110 18408 8116 18420
rect 8071 18380 8116 18408
rect 8110 18368 8116 18380
rect 8168 18368 8174 18420
rect 9214 18368 9220 18420
rect 9272 18408 9278 18420
rect 9861 18411 9919 18417
rect 9861 18408 9873 18411
rect 9272 18380 9873 18408
rect 9272 18368 9278 18380
rect 9861 18377 9873 18380
rect 9907 18377 9919 18411
rect 10502 18408 10508 18420
rect 10463 18380 10508 18408
rect 9861 18371 9919 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 12158 18368 12164 18420
rect 12216 18408 12222 18420
rect 12526 18408 12532 18420
rect 12216 18380 12532 18408
rect 12216 18368 12222 18380
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 15838 18408 15844 18420
rect 12636 18380 15844 18408
rect 10410 18300 10416 18352
rect 10468 18340 10474 18352
rect 11238 18340 11244 18352
rect 10468 18312 11244 18340
rect 10468 18300 10474 18312
rect 11238 18300 11244 18312
rect 11296 18300 11302 18352
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 12636 18340 12664 18380
rect 15838 18368 15844 18380
rect 15896 18368 15902 18420
rect 16850 18408 16856 18420
rect 16811 18380 16856 18408
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 17494 18408 17500 18420
rect 17455 18380 17500 18408
rect 17494 18368 17500 18380
rect 17552 18368 17558 18420
rect 17865 18411 17923 18417
rect 17865 18377 17877 18411
rect 17911 18408 17923 18411
rect 18138 18408 18144 18420
rect 17911 18380 18144 18408
rect 17911 18377 17923 18380
rect 17865 18371 17923 18377
rect 18138 18368 18144 18380
rect 18196 18408 18202 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 18196 18380 19809 18408
rect 18196 18368 18202 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 19981 18411 20039 18417
rect 19981 18377 19993 18411
rect 20027 18408 20039 18411
rect 20714 18408 20720 18420
rect 20027 18380 20720 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 11664 18312 12664 18340
rect 11664 18300 11670 18312
rect 4614 18272 4620 18284
rect 4264 18244 4620 18272
rect 4614 18232 4620 18244
rect 4672 18272 4678 18284
rect 5442 18272 5448 18284
rect 4672 18244 5448 18272
rect 4672 18232 4678 18244
rect 5442 18232 5448 18244
rect 5500 18272 5506 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5500 18244 5733 18272
rect 5500 18232 5506 18244
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 5721 18235 5779 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 11882 18272 11888 18284
rect 11256 18244 11888 18272
rect 2130 18164 2136 18216
rect 2188 18204 2194 18216
rect 2317 18207 2375 18213
rect 2317 18204 2329 18207
rect 2188 18176 2329 18204
rect 2188 18164 2194 18176
rect 2317 18173 2329 18176
rect 2363 18173 2375 18207
rect 2317 18167 2375 18173
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 8570 18204 8576 18216
rect 8527 18176 8576 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 8570 18164 8576 18176
rect 8628 18164 8634 18216
rect 11256 18213 11284 18244
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 18046 18232 18052 18284
rect 18104 18272 18110 18284
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 18104 18244 18521 18272
rect 18104 18232 18110 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 18509 18235 18567 18241
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18204 12311 18207
rect 12434 18204 12440 18216
rect 12299 18176 12440 18204
rect 12299 18173 12311 18176
rect 12253 18167 12311 18173
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 12802 18204 12808 18216
rect 12492 18176 12808 18204
rect 12492 18164 12498 18176
rect 12802 18164 12808 18176
rect 12860 18164 12866 18216
rect 12989 18207 13047 18213
rect 12989 18173 13001 18207
rect 13035 18204 13047 18207
rect 15378 18204 15384 18216
rect 13035 18176 15384 18204
rect 13035 18173 13047 18176
rect 12989 18167 13047 18173
rect 15378 18164 15384 18176
rect 15436 18204 15442 18216
rect 15473 18207 15531 18213
rect 15473 18204 15485 18207
rect 15436 18176 15485 18204
rect 15436 18164 15442 18176
rect 15473 18173 15485 18176
rect 15519 18173 15531 18207
rect 18414 18204 18420 18216
rect 18375 18176 18420 18204
rect 15473 18167 15531 18173
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 19812 18204 19840 18371
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 20990 18408 20996 18420
rect 20951 18380 20996 18408
rect 20990 18368 20996 18380
rect 21048 18368 21054 18420
rect 21450 18368 21456 18420
rect 21508 18408 21514 18420
rect 21818 18408 21824 18420
rect 21508 18380 21824 18408
rect 21508 18368 21514 18380
rect 21818 18368 21824 18380
rect 21876 18408 21882 18420
rect 22557 18411 22615 18417
rect 22557 18408 22569 18411
rect 21876 18380 22569 18408
rect 21876 18368 21882 18380
rect 22557 18377 22569 18380
rect 22603 18377 22615 18411
rect 23106 18408 23112 18420
rect 23067 18380 23112 18408
rect 22557 18371 22615 18377
rect 23106 18368 23112 18380
rect 23164 18408 23170 18420
rect 23382 18408 23388 18420
rect 23164 18380 23388 18408
rect 23164 18368 23170 18380
rect 23382 18368 23388 18380
rect 23440 18368 23446 18420
rect 25038 18408 25044 18420
rect 24999 18380 25044 18408
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 25130 18368 25136 18420
rect 25188 18408 25194 18420
rect 25590 18408 25596 18420
rect 25188 18380 25596 18408
rect 25188 18368 25194 18380
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 20530 18272 20536 18284
rect 20491 18244 20536 18272
rect 20530 18232 20536 18244
rect 20588 18272 20594 18284
rect 22097 18275 22155 18281
rect 22097 18272 22109 18275
rect 20588 18244 22109 18272
rect 20588 18232 20594 18244
rect 22097 18241 22109 18244
rect 22143 18241 22155 18275
rect 22097 18235 22155 18241
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 19812 18176 20453 18204
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 21913 18207 21971 18213
rect 21913 18204 21925 18207
rect 21048 18176 21925 18204
rect 21048 18164 21054 18176
rect 21913 18173 21925 18176
rect 21959 18173 21971 18207
rect 21913 18167 21971 18173
rect 23290 18164 23296 18216
rect 23348 18204 23354 18216
rect 23661 18207 23719 18213
rect 23661 18204 23673 18207
rect 23348 18176 23673 18204
rect 23348 18164 23354 18176
rect 23661 18173 23673 18176
rect 23707 18173 23719 18207
rect 23661 18167 23719 18173
rect 23750 18164 23756 18216
rect 23808 18204 23814 18216
rect 23917 18207 23975 18213
rect 23917 18204 23929 18207
rect 23808 18176 23929 18204
rect 23808 18164 23814 18176
rect 23917 18173 23929 18176
rect 23963 18204 23975 18207
rect 24762 18204 24768 18216
rect 23963 18176 24768 18204
rect 23963 18173 23975 18176
rect 23917 18167 23975 18173
rect 24762 18164 24768 18176
rect 24820 18164 24826 18216
rect 1946 18096 1952 18148
rect 2004 18136 2010 18148
rect 2562 18139 2620 18145
rect 2562 18136 2574 18139
rect 2004 18108 2574 18136
rect 2004 18096 2010 18108
rect 2562 18105 2574 18108
rect 2608 18105 2620 18139
rect 4709 18139 4767 18145
rect 2562 18099 2620 18105
rect 2700 18108 4660 18136
rect 1762 18028 1768 18080
rect 1820 18068 1826 18080
rect 2700 18068 2728 18108
rect 1820 18040 2728 18068
rect 3697 18071 3755 18077
rect 1820 18028 1826 18040
rect 3697 18037 3709 18071
rect 3743 18068 3755 18071
rect 4062 18068 4068 18080
rect 3743 18040 4068 18068
rect 3743 18037 3755 18040
rect 3697 18031 3755 18037
rect 4062 18028 4068 18040
rect 4120 18028 4126 18080
rect 4632 18068 4660 18108
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 5537 18139 5595 18145
rect 5537 18136 5549 18139
rect 4755 18108 5549 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 5537 18105 5549 18108
rect 5583 18136 5595 18139
rect 5718 18136 5724 18148
rect 5583 18108 5724 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 7193 18139 7251 18145
rect 7193 18105 7205 18139
rect 7239 18136 7251 18139
rect 7650 18136 7656 18148
rect 7239 18108 7656 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 7650 18096 7656 18108
rect 7708 18096 7714 18148
rect 8662 18096 8668 18148
rect 8720 18145 8726 18148
rect 8720 18139 8784 18145
rect 8720 18105 8738 18139
rect 8772 18136 8784 18139
rect 9122 18136 9128 18148
rect 8772 18108 9128 18136
rect 8772 18105 8784 18108
rect 8720 18099 8784 18105
rect 8720 18096 8726 18099
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 13256 18139 13314 18145
rect 13256 18105 13268 18139
rect 13302 18136 13314 18139
rect 13722 18136 13728 18148
rect 13302 18108 13728 18136
rect 13302 18105 13314 18108
rect 13256 18099 13314 18105
rect 13722 18096 13728 18108
rect 13780 18136 13786 18148
rect 14734 18136 14740 18148
rect 13780 18108 14740 18136
rect 13780 18096 13786 18108
rect 14734 18096 14740 18108
rect 14792 18136 14798 18148
rect 14921 18139 14979 18145
rect 14921 18136 14933 18139
rect 14792 18108 14933 18136
rect 14792 18096 14798 18108
rect 14921 18105 14933 18108
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 15740 18139 15798 18145
rect 15740 18105 15752 18139
rect 15786 18136 15798 18139
rect 21453 18139 21511 18145
rect 15786 18108 15820 18136
rect 15786 18105 15798 18108
rect 15740 18099 15798 18105
rect 21453 18105 21465 18139
rect 21499 18136 21511 18139
rect 22005 18139 22063 18145
rect 22005 18136 22017 18139
rect 21499 18108 22017 18136
rect 21499 18105 21511 18108
rect 21453 18099 21511 18105
rect 22005 18105 22017 18108
rect 22051 18105 22063 18139
rect 22005 18099 22063 18105
rect 4982 18068 4988 18080
rect 4632 18040 4988 18068
rect 4982 18028 4988 18040
rect 5040 18068 5046 18080
rect 5629 18071 5687 18077
rect 5629 18068 5641 18071
rect 5040 18040 5641 18068
rect 5040 18028 5046 18040
rect 5629 18037 5641 18040
rect 5675 18037 5687 18071
rect 6822 18068 6828 18080
rect 6783 18040 6828 18068
rect 5629 18031 5687 18037
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 7558 18068 7564 18080
rect 7331 18040 7564 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7558 18028 7564 18040
rect 7616 18028 7622 18080
rect 10778 18068 10784 18080
rect 10739 18040 10784 18068
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11422 18068 11428 18080
rect 11383 18040 11428 18068
rect 11422 18028 11428 18040
rect 11480 18028 11486 18080
rect 12526 18028 12532 18080
rect 12584 18068 12590 18080
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 12584 18040 12817 18068
rect 12584 18028 12590 18040
rect 12805 18037 12817 18040
rect 12851 18037 12863 18071
rect 12805 18031 12863 18037
rect 14090 18028 14096 18080
rect 14148 18068 14154 18080
rect 14369 18071 14427 18077
rect 14369 18068 14381 18071
rect 14148 18040 14381 18068
rect 14148 18028 14154 18040
rect 14369 18037 14381 18040
rect 14415 18068 14427 18071
rect 15102 18068 15108 18080
rect 14415 18040 15108 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 15102 18028 15108 18040
rect 15160 18028 15166 18080
rect 15381 18071 15439 18077
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15755 18068 15783 18099
rect 15838 18068 15844 18080
rect 15427 18040 15844 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15838 18028 15844 18040
rect 15896 18068 15902 18080
rect 16482 18068 16488 18080
rect 15896 18040 16488 18068
rect 15896 18028 15902 18040
rect 16482 18028 16488 18040
rect 16540 18028 16546 18080
rect 18046 18068 18052 18080
rect 18007 18040 18052 18068
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18966 18028 18972 18080
rect 19024 18068 19030 18080
rect 19061 18071 19119 18077
rect 19061 18068 19073 18071
rect 19024 18040 19073 18068
rect 19024 18028 19030 18040
rect 19061 18037 19073 18040
rect 19107 18037 19119 18071
rect 19061 18031 19119 18037
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 19208 18040 19533 18068
rect 19208 18028 19214 18040
rect 19521 18037 19533 18040
rect 19567 18068 19579 18071
rect 20349 18071 20407 18077
rect 20349 18068 20361 18071
rect 19567 18040 20361 18068
rect 19567 18037 19579 18040
rect 19521 18031 19579 18037
rect 20349 18037 20361 18040
rect 20395 18068 20407 18071
rect 20438 18068 20444 18080
rect 20395 18040 20444 18068
rect 20395 18037 20407 18040
rect 20349 18031 20407 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 21542 18068 21548 18080
rect 21503 18040 21548 18068
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 22020 18068 22048 18099
rect 22278 18068 22284 18080
rect 22020 18040 22284 18068
rect 22278 18028 22284 18040
rect 22336 18028 22342 18080
rect 23477 18071 23535 18077
rect 23477 18037 23489 18071
rect 23523 18068 23535 18071
rect 23750 18068 23756 18080
rect 23523 18040 23756 18068
rect 23523 18037 23535 18040
rect 23477 18031 23535 18037
rect 23750 18028 23756 18040
rect 23808 18068 23814 18080
rect 24118 18068 24124 18080
rect 23808 18040 24124 18068
rect 23808 18028 23814 18040
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1394 17824 1400 17876
rect 1452 17864 1458 17876
rect 1581 17867 1639 17873
rect 1581 17864 1593 17867
rect 1452 17836 1593 17864
rect 1452 17824 1458 17836
rect 1581 17833 1593 17836
rect 1627 17864 1639 17867
rect 1857 17867 1915 17873
rect 1857 17864 1869 17867
rect 1627 17836 1869 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1857 17833 1869 17836
rect 1903 17833 1915 17867
rect 1857 17827 1915 17833
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 3237 17867 3295 17873
rect 3237 17864 3249 17867
rect 2096 17836 3249 17864
rect 2096 17824 2102 17836
rect 3237 17833 3249 17836
rect 3283 17833 3295 17867
rect 5442 17864 5448 17876
rect 5403 17836 5448 17864
rect 3237 17827 3295 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 5592 17836 6745 17864
rect 5592 17824 5598 17836
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 8018 17864 8024 17876
rect 7979 17836 8024 17864
rect 6733 17827 6791 17833
rect 8018 17824 8024 17836
rect 8076 17824 8082 17876
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 8352 17836 8493 17864
rect 8352 17824 8358 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 10134 17864 10140 17876
rect 10047 17836 10140 17864
rect 8481 17827 8539 17833
rect 10134 17824 10140 17836
rect 10192 17864 10198 17876
rect 10870 17864 10876 17876
rect 10192 17836 10876 17864
rect 10192 17824 10198 17836
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11698 17824 11704 17876
rect 11756 17864 11762 17876
rect 12621 17867 12679 17873
rect 12621 17864 12633 17867
rect 11756 17836 12633 17864
rect 11756 17824 11762 17836
rect 12621 17833 12633 17836
rect 12667 17864 12679 17867
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 12667 17836 13553 17864
rect 12667 17833 12679 17836
rect 12621 17827 12679 17833
rect 13541 17833 13553 17836
rect 13587 17864 13599 17867
rect 13722 17864 13728 17876
rect 13587 17836 13728 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14734 17864 14740 17876
rect 14200 17836 14740 17864
rect 9122 17796 9128 17808
rect 9083 17768 9128 17796
rect 9122 17756 9128 17768
rect 9180 17796 9186 17808
rect 9401 17799 9459 17805
rect 9401 17796 9413 17799
rect 9180 17768 9413 17796
rect 9180 17756 9186 17768
rect 9401 17765 9413 17768
rect 9447 17765 9459 17799
rect 9401 17759 9459 17765
rect 2222 17728 2228 17740
rect 2183 17700 2228 17728
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17728 2375 17731
rect 2774 17728 2780 17740
rect 2363 17700 2780 17728
rect 2363 17697 2375 17700
rect 2317 17691 2375 17697
rect 2774 17688 2780 17700
rect 2832 17728 2838 17740
rect 3605 17731 3663 17737
rect 3605 17728 3617 17731
rect 2832 17700 3617 17728
rect 2832 17688 2838 17700
rect 3605 17697 3617 17700
rect 3651 17697 3663 17731
rect 3605 17691 3663 17697
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4321 17731 4379 17737
rect 4321 17728 4333 17731
rect 4212 17700 4333 17728
rect 4212 17688 4218 17700
rect 4321 17697 4333 17700
rect 4367 17697 4379 17731
rect 6546 17728 6552 17740
rect 6507 17700 6552 17728
rect 4321 17691 4379 17697
rect 6546 17688 6552 17700
rect 6604 17688 6610 17740
rect 8386 17728 8392 17740
rect 8347 17700 8392 17728
rect 8386 17688 8392 17700
rect 8444 17688 8450 17740
rect 2406 17660 2412 17672
rect 2367 17632 2412 17660
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 6457 17663 6515 17669
rect 4120 17632 4165 17660
rect 4120 17620 4126 17632
rect 6457 17629 6469 17663
rect 6503 17660 6515 17663
rect 6730 17660 6736 17672
rect 6503 17632 6736 17660
rect 6503 17629 6515 17632
rect 6457 17623 6515 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 8628 17632 8677 17660
rect 8628 17620 8634 17632
rect 8665 17629 8677 17632
rect 8711 17660 8723 17663
rect 9214 17660 9220 17672
rect 8711 17632 9220 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 9416 17660 9444 17759
rect 11146 17756 11152 17808
rect 11204 17796 11210 17808
rect 11508 17799 11566 17805
rect 11508 17796 11520 17799
rect 11204 17768 11520 17796
rect 11204 17756 11210 17768
rect 11508 17765 11520 17768
rect 11554 17796 11566 17799
rect 11882 17796 11888 17808
rect 11554 17768 11888 17796
rect 11554 17765 11566 17768
rect 11508 17759 11566 17765
rect 11882 17756 11888 17768
rect 11940 17796 11946 17808
rect 13173 17799 13231 17805
rect 13173 17796 13185 17799
rect 11940 17768 13185 17796
rect 11940 17756 11946 17768
rect 13173 17765 13185 17768
rect 13219 17796 13231 17799
rect 13262 17796 13268 17808
rect 13219 17768 13268 17796
rect 13219 17765 13231 17768
rect 13173 17759 13231 17765
rect 13262 17756 13268 17768
rect 13320 17756 13326 17808
rect 14200 17805 14228 17836
rect 14734 17824 14740 17836
rect 14792 17824 14798 17876
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 16669 17867 16727 17873
rect 16669 17864 16681 17867
rect 16632 17836 16681 17864
rect 16632 17824 16638 17836
rect 16669 17833 16681 17836
rect 16715 17833 16727 17867
rect 16669 17827 16727 17833
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18046 17864 18052 17876
rect 17359 17836 18052 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18046 17824 18052 17836
rect 18104 17864 18110 17876
rect 18233 17867 18291 17873
rect 18233 17864 18245 17867
rect 18104 17836 18245 17864
rect 18104 17824 18110 17836
rect 18233 17833 18245 17836
rect 18279 17833 18291 17867
rect 18233 17827 18291 17833
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 18785 17867 18843 17873
rect 18785 17864 18797 17867
rect 18748 17836 18797 17864
rect 18748 17824 18754 17836
rect 18785 17833 18797 17836
rect 18831 17833 18843 17867
rect 18785 17827 18843 17833
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 21542 17864 21548 17876
rect 20763 17836 21548 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 21542 17824 21548 17836
rect 21600 17824 21606 17876
rect 22646 17864 22652 17876
rect 22607 17836 22652 17864
rect 22646 17824 22652 17836
rect 22704 17824 22710 17876
rect 23566 17864 23572 17876
rect 23527 17836 23572 17864
rect 23566 17824 23572 17836
rect 23624 17824 23630 17876
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25041 17867 25099 17873
rect 25041 17864 25053 17867
rect 24912 17836 25053 17864
rect 24912 17824 24918 17836
rect 25041 17833 25053 17836
rect 25087 17833 25099 17867
rect 25041 17827 25099 17833
rect 14185 17799 14243 17805
rect 14185 17765 14197 17799
rect 14231 17765 14243 17799
rect 14185 17759 14243 17765
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15534 17799 15592 17805
rect 15534 17796 15546 17799
rect 15252 17768 15546 17796
rect 15252 17756 15258 17768
rect 15534 17765 15546 17768
rect 15580 17796 15592 17799
rect 15930 17796 15936 17808
rect 15580 17768 15936 17796
rect 15580 17765 15592 17768
rect 15534 17759 15592 17765
rect 15930 17756 15936 17768
rect 15988 17756 15994 17808
rect 17681 17799 17739 17805
rect 17681 17765 17693 17799
rect 17727 17796 17739 17799
rect 17862 17796 17868 17808
rect 17727 17768 17868 17796
rect 17727 17765 17739 17768
rect 17681 17759 17739 17765
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 18506 17756 18512 17808
rect 18564 17796 18570 17808
rect 19153 17799 19211 17805
rect 19153 17796 19165 17799
rect 18564 17768 19165 17796
rect 18564 17756 18570 17768
rect 19153 17765 19165 17768
rect 19199 17765 19211 17799
rect 19153 17759 19211 17765
rect 19518 17756 19524 17808
rect 19576 17796 19582 17808
rect 19613 17799 19671 17805
rect 19613 17796 19625 17799
rect 19576 17768 19625 17796
rect 19576 17756 19582 17768
rect 19613 17765 19625 17768
rect 19659 17765 19671 17799
rect 21358 17796 21364 17808
rect 21319 17768 21364 17796
rect 19613 17759 19671 17765
rect 21358 17756 21364 17768
rect 21416 17756 21422 17808
rect 23842 17756 23848 17808
rect 23900 17805 23906 17808
rect 23900 17799 23964 17805
rect 23900 17765 23918 17799
rect 23952 17765 23964 17799
rect 23900 17759 23964 17765
rect 23900 17756 23906 17759
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 10008 17700 10057 17728
rect 10008 17688 10014 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 11238 17728 11244 17740
rect 11151 17700 11244 17728
rect 10045 17691 10103 17697
rect 11238 17688 11244 17700
rect 11296 17728 11302 17740
rect 12342 17728 12348 17740
rect 11296 17700 12348 17728
rect 11296 17688 11302 17700
rect 12342 17688 12348 17700
rect 12400 17688 12406 17740
rect 13909 17731 13967 17737
rect 13909 17697 13921 17731
rect 13955 17728 13967 17731
rect 14550 17728 14556 17740
rect 13955 17700 14556 17728
rect 13955 17697 13967 17700
rect 13909 17691 13967 17697
rect 14550 17688 14556 17700
rect 14608 17728 14614 17740
rect 15102 17728 15108 17740
rect 14608 17700 15108 17728
rect 14608 17688 14614 17700
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 15289 17731 15347 17737
rect 15289 17697 15301 17731
rect 15335 17728 15347 17731
rect 15378 17728 15384 17740
rect 15335 17700 15384 17728
rect 15335 17697 15347 17700
rect 15289 17691 15347 17697
rect 15378 17688 15384 17700
rect 15436 17728 15442 17740
rect 17034 17728 17040 17740
rect 15436 17700 17040 17728
rect 15436 17688 15442 17700
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 18046 17688 18052 17740
rect 18104 17728 18110 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 18104 17700 18153 17728
rect 18104 17688 18110 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 19337 17731 19395 17737
rect 19337 17697 19349 17731
rect 19383 17728 19395 17731
rect 19426 17728 19432 17740
rect 19383 17700 19432 17728
rect 19383 17697 19395 17700
rect 19337 17691 19395 17697
rect 19426 17688 19432 17700
rect 19484 17728 19490 17740
rect 19484 17700 20944 17728
rect 19484 17688 19490 17700
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 9416 17632 10333 17660
rect 10321 17629 10333 17632
rect 10367 17660 10379 17663
rect 10962 17660 10968 17672
rect 10367 17632 10968 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 18322 17660 18328 17672
rect 18283 17632 18328 17660
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 6089 17595 6147 17601
rect 6089 17561 6101 17595
rect 6135 17592 6147 17595
rect 7650 17592 7656 17604
rect 6135 17564 7656 17592
rect 6135 17561 6147 17564
rect 6089 17555 6147 17561
rect 7650 17552 7656 17564
rect 7708 17552 7714 17604
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 9677 17595 9735 17601
rect 9677 17592 9689 17595
rect 8444 17564 9689 17592
rect 8444 17552 8450 17564
rect 9677 17561 9689 17564
rect 9723 17561 9735 17595
rect 9677 17555 9735 17561
rect 13814 17552 13820 17604
rect 13872 17592 13878 17604
rect 14550 17592 14556 17604
rect 13872 17564 14556 17592
rect 13872 17552 13878 17564
rect 14550 17552 14556 17564
rect 14608 17552 14614 17604
rect 14918 17592 14924 17604
rect 14879 17564 14924 17592
rect 14918 17552 14924 17564
rect 14976 17552 14982 17604
rect 17770 17592 17776 17604
rect 17731 17564 17776 17592
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 20916 17601 20944 17700
rect 21082 17688 21088 17740
rect 21140 17728 21146 17740
rect 21269 17731 21327 17737
rect 21269 17728 21281 17731
rect 21140 17700 21281 17728
rect 21140 17688 21146 17700
rect 21269 17697 21281 17700
rect 21315 17697 21327 17731
rect 21269 17691 21327 17697
rect 22465 17731 22523 17737
rect 22465 17697 22477 17731
rect 22511 17728 22523 17731
rect 22922 17728 22928 17740
rect 22511 17700 22928 17728
rect 22511 17697 22523 17700
rect 22465 17691 22523 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 20990 17620 20996 17672
rect 21048 17660 21054 17672
rect 21453 17663 21511 17669
rect 21453 17660 21465 17663
rect 21048 17632 21465 17660
rect 21048 17620 21054 17632
rect 21453 17629 21465 17632
rect 21499 17629 21511 17663
rect 21453 17623 21511 17629
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23532 17632 23673 17660
rect 23532 17620 23538 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 20901 17595 20959 17601
rect 20901 17561 20913 17595
rect 20947 17561 20959 17595
rect 20901 17555 20959 17561
rect 2958 17524 2964 17536
rect 2871 17496 2964 17524
rect 2958 17484 2964 17496
rect 3016 17524 3022 17536
rect 3510 17524 3516 17536
rect 3016 17496 3516 17524
rect 3016 17484 3022 17496
rect 3510 17484 3516 17496
rect 3568 17484 3574 17536
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 6788 17496 7113 17524
rect 6788 17484 6794 17496
rect 7101 17493 7113 17496
rect 7147 17524 7159 17527
rect 7374 17524 7380 17536
rect 7147 17496 7380 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 7558 17524 7564 17536
rect 7519 17496 7564 17524
rect 7558 17484 7564 17496
rect 7616 17484 7622 17536
rect 7926 17524 7932 17536
rect 7887 17496 7932 17524
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 9490 17524 9496 17536
rect 9272 17496 9496 17524
rect 9272 17484 9278 17496
rect 9490 17484 9496 17496
rect 9548 17484 9554 17536
rect 10870 17524 10876 17536
rect 10831 17496 10876 17524
rect 10870 17484 10876 17496
rect 10928 17484 10934 17536
rect 20165 17527 20223 17533
rect 20165 17493 20177 17527
rect 20211 17524 20223 17527
rect 20530 17524 20536 17536
rect 20211 17496 20536 17524
rect 20211 17493 20223 17496
rect 20165 17487 20223 17493
rect 20530 17484 20536 17496
rect 20588 17524 20594 17536
rect 21913 17527 21971 17533
rect 21913 17524 21925 17527
rect 20588 17496 21925 17524
rect 20588 17484 20594 17496
rect 21913 17493 21925 17496
rect 21959 17493 21971 17527
rect 21913 17487 21971 17493
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2406 17320 2412 17332
rect 1995 17292 2412 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2406 17280 2412 17292
rect 2464 17320 2470 17332
rect 4154 17320 4160 17332
rect 2464 17292 4160 17320
rect 2464 17280 2470 17292
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 4614 17320 4620 17332
rect 4575 17292 4620 17320
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 4890 17320 4896 17332
rect 4851 17292 4896 17320
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 5074 17320 5080 17332
rect 5035 17292 5080 17320
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 6086 17320 6092 17332
rect 6047 17292 6092 17320
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6178 17280 6184 17332
rect 6236 17320 6242 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6236 17292 6561 17320
rect 6236 17280 6242 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5629 17187 5687 17193
rect 5629 17184 5641 17187
rect 5500 17156 5641 17184
rect 5500 17144 5506 17156
rect 5629 17153 5641 17156
rect 5675 17153 5687 17187
rect 5629 17147 5687 17153
rect 2130 17116 2136 17128
rect 2043 17088 2136 17116
rect 2130 17076 2136 17088
rect 2188 17116 2194 17128
rect 4062 17116 4068 17128
rect 2188 17088 4068 17116
rect 2188 17076 2194 17088
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4890 17076 4896 17128
rect 4948 17116 4954 17128
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 4948 17088 5549 17116
rect 4948 17076 4954 17088
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 6564 17116 6592 17283
rect 9490 17280 9496 17332
rect 9548 17320 9554 17332
rect 9674 17320 9680 17332
rect 9548 17292 9680 17320
rect 9548 17280 9554 17292
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 10134 17280 10140 17332
rect 10192 17320 10198 17332
rect 10229 17323 10287 17329
rect 10229 17320 10241 17323
rect 10192 17292 10241 17320
rect 10192 17280 10198 17292
rect 10229 17289 10241 17292
rect 10275 17289 10287 17323
rect 10229 17283 10287 17289
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 13170 17320 13176 17332
rect 11204 17292 13176 17320
rect 11204 17280 11210 17292
rect 13170 17280 13176 17292
rect 13228 17280 13234 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 13872 17292 14933 17320
rect 13872 17280 13878 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 15930 17320 15936 17332
rect 15891 17292 15936 17320
rect 14921 17283 14979 17289
rect 15930 17280 15936 17292
rect 15988 17280 15994 17332
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17320 17923 17323
rect 18322 17320 18328 17332
rect 17911 17292 18328 17320
rect 17911 17289 17923 17292
rect 17865 17283 17923 17289
rect 18322 17280 18328 17292
rect 18380 17280 18386 17332
rect 19981 17323 20039 17329
rect 19981 17289 19993 17323
rect 20027 17320 20039 17323
rect 21082 17320 21088 17332
rect 20027 17292 21088 17320
rect 20027 17289 20039 17292
rect 19981 17283 20039 17289
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 21358 17280 21364 17332
rect 21416 17320 21422 17332
rect 22373 17323 22431 17329
rect 22373 17320 22385 17323
rect 21416 17292 22385 17320
rect 21416 17280 21422 17292
rect 22373 17289 22385 17292
rect 22419 17289 22431 17323
rect 22373 17283 22431 17289
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 23155 17292 23489 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 23477 17289 23489 17292
rect 23523 17320 23535 17323
rect 23842 17320 23848 17332
rect 23523 17292 23848 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23842 17280 23848 17292
rect 23900 17320 23906 17332
rect 23900 17292 24348 17320
rect 23900 17280 23906 17292
rect 7006 17252 7012 17264
rect 6967 17224 7012 17252
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 14642 17212 14648 17264
rect 14700 17252 14706 17264
rect 14737 17255 14795 17261
rect 14737 17252 14749 17255
rect 14700 17224 14749 17252
rect 14700 17212 14706 17224
rect 14737 17221 14749 17224
rect 14783 17221 14795 17255
rect 21818 17252 21824 17264
rect 21779 17224 21824 17252
rect 14737 17215 14795 17221
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7791 17156 8125 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 8113 17153 8125 17156
rect 8159 17184 8171 17187
rect 8159 17156 8432 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6564 17088 6837 17116
rect 5537 17079 5595 17085
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17085 8355 17119
rect 8404 17116 8432 17156
rect 10870 17144 10876 17196
rect 10928 17184 10934 17196
rect 11054 17184 11060 17196
rect 10928 17156 11060 17184
rect 10928 17144 10934 17156
rect 11054 17144 11060 17156
rect 11112 17184 11118 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11112 17156 11345 17184
rect 11112 17144 11118 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12400 17156 12449 17184
rect 12400 17144 12406 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 8570 17125 8576 17128
rect 8564 17116 8576 17125
rect 8404 17088 8576 17116
rect 8297 17079 8355 17085
rect 8564 17079 8576 17088
rect 2400 17051 2458 17057
rect 2400 17017 2412 17051
rect 2446 17048 2458 17051
rect 2498 17048 2504 17060
rect 2446 17020 2504 17048
rect 2446 17017 2458 17020
rect 2400 17011 2458 17017
rect 2498 17008 2504 17020
rect 2556 17008 2562 17060
rect 8110 17008 8116 17060
rect 8168 17048 8174 17060
rect 8312 17048 8340 17079
rect 8570 17076 8576 17079
rect 8628 17076 8634 17128
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10778 17116 10784 17128
rect 9732 17088 10784 17116
rect 9732 17076 9738 17088
rect 10778 17076 10784 17088
rect 10836 17116 10842 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 10836 17088 11253 17116
rect 10836 17076 10842 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 14752 17116 14780 17215
rect 21818 17212 21824 17224
rect 21876 17212 21882 17264
rect 23661 17255 23719 17261
rect 23661 17221 23673 17255
rect 23707 17221 23719 17255
rect 23661 17215 23719 17221
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15473 17187 15531 17193
rect 15473 17184 15485 17187
rect 14884 17156 15485 17184
rect 14884 17144 14890 17156
rect 15473 17153 15485 17156
rect 15519 17153 15531 17187
rect 15473 17147 15531 17153
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17184 17555 17187
rect 18690 17184 18696 17196
rect 17543 17156 18696 17184
rect 17543 17153 17555 17156
rect 17497 17147 17555 17153
rect 18690 17144 18696 17156
rect 18748 17144 18754 17196
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 14752 17088 15301 17116
rect 11241 17079 11299 17085
rect 15289 17085 15301 17088
rect 15335 17085 15347 17119
rect 16485 17119 16543 17125
rect 16485 17116 16497 17119
rect 15289 17079 15347 17085
rect 16316 17088 16497 17116
rect 9858 17048 9864 17060
rect 8168 17020 9864 17048
rect 8168 17008 8174 17020
rect 9858 17008 9864 17020
rect 9916 17008 9922 17060
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 11422 17048 11428 17060
rect 10928 17020 11428 17048
rect 10928 17008 10934 17020
rect 11422 17008 11428 17020
rect 11480 17048 11486 17060
rect 12253 17051 12311 17057
rect 12253 17048 12265 17051
rect 11480 17020 12265 17048
rect 11480 17008 11486 17020
rect 12253 17017 12265 17020
rect 12299 17048 12311 17051
rect 12618 17048 12624 17060
rect 12299 17020 12624 17048
rect 12299 17017 12311 17020
rect 12253 17011 12311 17017
rect 12618 17008 12624 17020
rect 12676 17057 12682 17060
rect 12676 17051 12740 17057
rect 12676 17017 12694 17051
rect 12728 17017 12740 17051
rect 12676 17011 12740 17017
rect 12676 17008 12682 17011
rect 14918 17008 14924 17060
rect 14976 17048 14982 17060
rect 15381 17051 15439 17057
rect 15381 17048 15393 17051
rect 14976 17020 15393 17048
rect 14976 17008 14982 17020
rect 15381 17017 15393 17020
rect 15427 17017 15439 17051
rect 15381 17011 15439 17017
rect 16316 16992 16344 17088
rect 16485 17085 16497 17088
rect 16531 17085 16543 17119
rect 20438 17116 20444 17128
rect 20399 17088 20444 17116
rect 16485 17079 16543 17085
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 23676 17116 23704 17215
rect 24320 17196 24348 17292
rect 24302 17184 24308 17196
rect 24263 17156 24308 17184
rect 24302 17144 24308 17156
rect 24360 17144 24366 17196
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 23676 17088 25237 17116
rect 25225 17085 25237 17088
rect 25271 17116 25283 17119
rect 25961 17119 26019 17125
rect 25961 17116 25973 17119
rect 25271 17088 25973 17116
rect 25271 17085 25283 17088
rect 25225 17079 25283 17085
rect 25961 17085 25973 17088
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 16761 17051 16819 17057
rect 16761 17017 16773 17051
rect 16807 17048 16819 17051
rect 17126 17048 17132 17060
rect 16807 17020 17132 17048
rect 16807 17017 16819 17020
rect 16761 17011 16819 17017
rect 17126 17008 17132 17020
rect 17184 17008 17190 17060
rect 18230 17008 18236 17060
rect 18288 17048 18294 17060
rect 18417 17051 18475 17057
rect 18417 17048 18429 17051
rect 18288 17020 18429 17048
rect 18288 17008 18294 17020
rect 18417 17017 18429 17020
rect 18463 17048 18475 17051
rect 19429 17051 19487 17057
rect 19429 17048 19441 17051
rect 18463 17020 19441 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 19429 17017 19441 17020
rect 19475 17017 19487 17051
rect 19429 17011 19487 17017
rect 20530 17008 20536 17060
rect 20588 17048 20594 17060
rect 20686 17051 20744 17057
rect 20686 17048 20698 17051
rect 20588 17020 20698 17048
rect 20588 17008 20594 17020
rect 20686 17017 20698 17020
rect 20732 17017 20744 17051
rect 20686 17011 20744 17017
rect 23750 17008 23756 17060
rect 23808 17048 23814 17060
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 23808 17020 24041 17048
rect 23808 17008 23814 17020
rect 24029 17017 24041 17020
rect 24075 17048 24087 17051
rect 25041 17051 25099 17057
rect 25041 17048 25053 17051
rect 24075 17020 25053 17048
rect 24075 17017 24087 17020
rect 24029 17011 24087 17017
rect 25041 17017 25053 17020
rect 25087 17017 25099 17051
rect 25041 17011 25099 17017
rect 25130 17008 25136 17060
rect 25188 17048 25194 17060
rect 25501 17051 25559 17057
rect 25501 17048 25513 17051
rect 25188 17020 25513 17048
rect 25188 17008 25194 17020
rect 25501 17017 25513 17020
rect 25547 17017 25559 17051
rect 25501 17011 25559 17017
rect 3510 16980 3516 16992
rect 3471 16952 3516 16980
rect 3510 16940 3516 16952
rect 3568 16940 3574 16992
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 5445 16983 5503 16989
rect 5445 16980 5457 16983
rect 5224 16952 5457 16980
rect 5224 16940 5230 16952
rect 5445 16949 5457 16952
rect 5491 16949 5503 16983
rect 5445 16943 5503 16949
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10192 16952 10609 16980
rect 10192 16940 10198 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 10597 16943 10655 16949
rect 10781 16983 10839 16989
rect 10781 16949 10793 16983
rect 10827 16980 10839 16983
rect 10962 16980 10968 16992
rect 10827 16952 10968 16980
rect 10827 16949 10839 16952
rect 10781 16943 10839 16949
rect 10962 16940 10968 16952
rect 11020 16940 11026 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11882 16980 11888 16992
rect 11843 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16980 11946 16992
rect 13817 16983 13875 16989
rect 13817 16980 13829 16983
rect 11940 16952 13829 16980
rect 11940 16940 11946 16952
rect 13817 16949 13829 16952
rect 13863 16949 13875 16983
rect 14366 16980 14372 16992
rect 14327 16952 14372 16980
rect 13817 16943 13875 16949
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 16298 16980 16304 16992
rect 16259 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 18506 16980 18512 16992
rect 18467 16952 18512 16980
rect 18506 16940 18512 16952
rect 18564 16980 18570 16992
rect 19061 16983 19119 16989
rect 19061 16980 19073 16983
rect 18564 16952 19073 16980
rect 18564 16940 18570 16952
rect 19061 16949 19073 16952
rect 19107 16949 19119 16983
rect 19061 16943 19119 16949
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20898 16980 20904 16992
rect 20395 16952 20904 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 24118 16980 24124 16992
rect 24079 16952 24124 16980
rect 24118 16940 24124 16952
rect 24176 16980 24182 16992
rect 24673 16983 24731 16989
rect 24673 16980 24685 16983
rect 24176 16952 24685 16980
rect 24176 16940 24182 16952
rect 24673 16949 24685 16952
rect 24719 16949 24731 16983
rect 24673 16943 24731 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1857 16779 1915 16785
rect 1857 16745 1869 16779
rect 1903 16776 1915 16779
rect 2222 16776 2228 16788
rect 1903 16748 2228 16776
rect 1903 16745 1915 16748
rect 1857 16739 1915 16745
rect 2222 16736 2228 16748
rect 2280 16736 2286 16788
rect 2958 16776 2964 16788
rect 2792 16748 2964 16776
rect 2038 16668 2044 16720
rect 2096 16708 2102 16720
rect 2317 16711 2375 16717
rect 2317 16708 2329 16711
rect 2096 16680 2329 16708
rect 2096 16668 2102 16680
rect 2317 16677 2329 16680
rect 2363 16677 2375 16711
rect 2317 16671 2375 16677
rect 2498 16668 2504 16720
rect 2556 16708 2562 16720
rect 2792 16708 2820 16748
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 3510 16776 3516 16788
rect 3375 16748 3516 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 5166 16776 5172 16788
rect 4580 16748 5172 16776
rect 4580 16736 4586 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6730 16776 6736 16788
rect 6691 16748 6736 16776
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 8021 16779 8079 16785
rect 8021 16776 8033 16779
rect 6972 16748 8033 16776
rect 6972 16736 6978 16748
rect 8021 16745 8033 16748
rect 8067 16745 8079 16779
rect 8021 16739 8079 16745
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9033 16779 9091 16785
rect 9033 16776 9045 16779
rect 8352 16748 9045 16776
rect 8352 16736 8358 16748
rect 9033 16745 9045 16748
rect 9079 16745 9091 16779
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9033 16739 9091 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10134 16776 10140 16788
rect 10095 16748 10140 16776
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10870 16776 10876 16788
rect 10831 16748 10876 16776
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 14918 16776 14924 16788
rect 14879 16748 14924 16776
rect 14918 16736 14924 16748
rect 14976 16736 14982 16788
rect 15289 16779 15347 16785
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 16298 16776 16304 16788
rect 15335 16748 16304 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18969 16779 19027 16785
rect 18969 16776 18981 16779
rect 18104 16748 18981 16776
rect 18104 16736 18110 16748
rect 18969 16745 18981 16748
rect 19015 16745 19027 16779
rect 19426 16776 19432 16788
rect 19387 16748 19432 16776
rect 18969 16739 19027 16745
rect 19426 16736 19432 16748
rect 19484 16736 19490 16788
rect 19705 16779 19763 16785
rect 19705 16745 19717 16779
rect 19751 16776 19763 16779
rect 19978 16776 19984 16788
rect 19751 16748 19984 16776
rect 19751 16745 19763 16748
rect 19705 16739 19763 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 20898 16736 20904 16788
rect 20956 16776 20962 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 20956 16748 22293 16776
rect 20956 16736 20962 16748
rect 22281 16745 22293 16748
rect 22327 16745 22339 16779
rect 22922 16776 22928 16788
rect 22883 16748 22928 16776
rect 22281 16739 22339 16745
rect 22922 16736 22928 16748
rect 22980 16736 22986 16788
rect 23290 16776 23296 16788
rect 23251 16748 23296 16776
rect 23290 16736 23296 16748
rect 23348 16736 23354 16788
rect 24302 16736 24308 16788
rect 24360 16776 24366 16788
rect 25133 16779 25191 16785
rect 25133 16776 25145 16779
rect 24360 16748 25145 16776
rect 24360 16736 24366 16748
rect 25133 16745 25145 16748
rect 25179 16745 25191 16779
rect 25133 16739 25191 16745
rect 2556 16680 2820 16708
rect 2556 16668 2562 16680
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 1854 16640 1860 16652
rect 1811 16612 1860 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 2004 16612 2237 16640
rect 2004 16600 2010 16612
rect 2225 16609 2237 16612
rect 2271 16609 2283 16643
rect 2792 16640 2820 16680
rect 2866 16668 2872 16720
rect 2924 16708 2930 16720
rect 3605 16711 3663 16717
rect 3605 16708 3617 16711
rect 2924 16680 3617 16708
rect 2924 16668 2930 16680
rect 3605 16677 3617 16680
rect 3651 16677 3663 16711
rect 3605 16671 3663 16677
rect 4341 16711 4399 16717
rect 4341 16677 4353 16711
rect 4387 16708 4399 16711
rect 6546 16708 6552 16720
rect 4387 16680 6552 16708
rect 4387 16677 4399 16680
rect 4341 16671 4399 16677
rect 6546 16668 6552 16680
rect 6604 16708 6610 16720
rect 7285 16711 7343 16717
rect 7285 16708 7297 16711
rect 6604 16680 7297 16708
rect 6604 16668 6610 16680
rect 7285 16677 7297 16680
rect 7331 16677 7343 16711
rect 7285 16671 7343 16677
rect 8481 16711 8539 16717
rect 8481 16677 8493 16711
rect 8527 16708 8539 16711
rect 8570 16708 8576 16720
rect 8527 16680 8576 16708
rect 8527 16677 8539 16680
rect 8481 16671 8539 16677
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 9950 16708 9956 16720
rect 9539 16680 9956 16708
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 9950 16668 9956 16680
rect 10008 16708 10014 16720
rect 10686 16708 10692 16720
rect 10008 16680 10692 16708
rect 10008 16668 10014 16680
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 14185 16711 14243 16717
rect 14185 16677 14197 16711
rect 14231 16708 14243 16711
rect 14826 16708 14832 16720
rect 14231 16680 14832 16708
rect 14231 16677 14243 16680
rect 14185 16671 14243 16677
rect 14826 16668 14832 16680
rect 14884 16668 14890 16720
rect 15470 16668 15476 16720
rect 15528 16708 15534 16720
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 15528 16680 15761 16708
rect 15528 16668 15534 16680
rect 15749 16677 15761 16680
rect 15795 16708 15807 16711
rect 16761 16711 16819 16717
rect 16761 16708 16773 16711
rect 15795 16680 16773 16708
rect 15795 16677 15807 16680
rect 15749 16671 15807 16677
rect 16761 16677 16773 16680
rect 16807 16677 16819 16711
rect 16761 16671 16819 16677
rect 17304 16711 17362 16717
rect 17304 16677 17316 16711
rect 17350 16708 17362 16711
rect 17494 16708 17500 16720
rect 17350 16680 17500 16708
rect 17350 16677 17362 16680
rect 17304 16671 17362 16677
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21168 16711 21226 16717
rect 21168 16708 21180 16711
rect 20772 16680 21180 16708
rect 20772 16668 20778 16680
rect 21168 16677 21180 16680
rect 21214 16708 21226 16711
rect 21818 16708 21824 16720
rect 21214 16680 21824 16708
rect 21214 16677 21226 16680
rect 21168 16671 21226 16677
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2792 16612 2973 16640
rect 2225 16603 2283 16609
rect 2961 16609 2973 16612
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5620 16643 5678 16649
rect 5620 16609 5632 16643
rect 5666 16640 5678 16643
rect 6178 16640 6184 16652
rect 5666 16612 6184 16640
rect 5666 16609 5678 16612
rect 5620 16603 5678 16609
rect 1872 16572 1900 16600
rect 2409 16575 2467 16581
rect 2409 16572 2421 16575
rect 1872 16544 2421 16572
rect 2409 16541 2421 16544
rect 2455 16572 2467 16575
rect 3510 16572 3516 16584
rect 2455 16544 3516 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 4080 16572 4108 16603
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 8312 16612 8401 16640
rect 4430 16572 4436 16584
rect 4080 16544 4436 16572
rect 4430 16532 4436 16544
rect 4488 16532 4494 16584
rect 5350 16572 5356 16584
rect 5311 16544 5356 16572
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 7742 16532 7748 16584
rect 7800 16572 7806 16584
rect 8312 16572 8340 16612
rect 8389 16609 8401 16612
rect 8435 16640 8447 16643
rect 9306 16640 9312 16652
rect 8435 16612 9312 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 9306 16600 9312 16612
rect 9364 16640 9370 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9364 16612 10057 16640
rect 9364 16600 9370 16612
rect 10045 16609 10057 16612
rect 10091 16640 10103 16643
rect 10502 16640 10508 16652
rect 10091 16612 10508 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10502 16600 10508 16612
rect 10560 16600 10566 16652
rect 11238 16640 11244 16652
rect 11199 16612 11244 16640
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11508 16643 11566 16649
rect 11508 16609 11520 16643
rect 11554 16640 11566 16643
rect 11790 16640 11796 16652
rect 11554 16612 11796 16640
rect 11554 16609 11566 16612
rect 11508 16603 11566 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12802 16640 12808 16652
rect 12676 16612 12808 16640
rect 12676 16600 12682 16612
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16640 13507 16643
rect 13909 16643 13967 16649
rect 13495 16612 13860 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 7800 16544 8340 16572
rect 8665 16575 8723 16581
rect 7800 16532 7806 16544
rect 8665 16541 8677 16575
rect 8711 16572 8723 16575
rect 9582 16572 9588 16584
rect 8711 16544 9588 16572
rect 8711 16541 8723 16544
rect 8665 16535 8723 16541
rect 7926 16504 7932 16516
rect 7839 16476 7932 16504
rect 7926 16464 7932 16476
rect 7984 16504 7990 16516
rect 8680 16504 8708 16535
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10226 16532 10232 16584
rect 10284 16572 10290 16584
rect 10284 16544 10329 16572
rect 10284 16532 10290 16544
rect 7984 16476 8708 16504
rect 13832 16504 13860 16612
rect 13909 16609 13921 16643
rect 13955 16640 13967 16643
rect 13998 16640 14004 16652
rect 13955 16612 14004 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14366 16600 14372 16652
rect 14424 16640 14430 16652
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 14424 16612 15669 16640
rect 14424 16600 14430 16612
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 17034 16640 17040 16652
rect 16995 16612 17040 16640
rect 15657 16603 15715 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 19392 16612 19533 16640
rect 19392 16600 19398 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 20530 16640 20536 16652
rect 20491 16612 20536 16640
rect 19521 16603 19579 16609
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 23474 16640 23480 16652
rect 23387 16612 23480 16640
rect 15838 16572 15844 16584
rect 15799 16544 15844 16572
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16572 20223 16575
rect 20438 16572 20444 16584
rect 20211 16544 20444 16572
rect 20211 16541 20223 16544
rect 20165 16535 20223 16541
rect 20438 16532 20444 16544
rect 20496 16572 20502 16584
rect 20806 16572 20812 16584
rect 20496 16544 20812 16572
rect 20496 16532 20502 16544
rect 20806 16532 20812 16544
rect 20864 16572 20870 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20864 16544 20913 16572
rect 20864 16532 20870 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 23290 16532 23296 16584
rect 23348 16572 23354 16584
rect 23400 16572 23428 16612
rect 23474 16600 23480 16612
rect 23532 16640 23538 16652
rect 24026 16649 24032 16652
rect 23569 16643 23627 16649
rect 23569 16640 23581 16643
rect 23532 16612 23581 16640
rect 23532 16600 23538 16612
rect 23569 16609 23581 16612
rect 23615 16640 23627 16643
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23615 16612 23765 16640
rect 23615 16609 23627 16612
rect 23569 16603 23627 16609
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 24020 16603 24032 16649
rect 24084 16640 24090 16652
rect 24084 16612 24120 16640
rect 24026 16600 24032 16603
rect 24084 16600 24090 16612
rect 23348 16544 23428 16572
rect 23348 16532 23354 16544
rect 14182 16504 14188 16516
rect 13832 16476 14188 16504
rect 7984 16464 7990 16476
rect 14182 16464 14188 16476
rect 14240 16464 14246 16516
rect 18417 16507 18475 16513
rect 18417 16473 18429 16507
rect 18463 16504 18475 16507
rect 18690 16504 18696 16516
rect 18463 16476 18696 16504
rect 18463 16473 18475 16476
rect 18417 16467 18475 16473
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 13817 16439 13875 16445
rect 13817 16405 13829 16439
rect 13863 16436 13875 16439
rect 14458 16436 14464 16448
rect 13863 16408 14464 16436
rect 13863 16405 13875 16408
rect 13817 16399 13875 16405
rect 14458 16396 14464 16408
rect 14516 16396 14522 16448
rect 16485 16439 16543 16445
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 16574 16436 16580 16448
rect 16531 16408 16580 16436
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 16574 16396 16580 16408
rect 16632 16396 16638 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2498 16232 2504 16244
rect 2459 16204 2504 16232
rect 2498 16192 2504 16204
rect 2556 16192 2562 16244
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 6270 16232 6276 16244
rect 2832 16204 2877 16232
rect 6231 16204 6276 16232
rect 2832 16192 2838 16204
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 6638 16232 6644 16244
rect 6599 16204 6644 16232
rect 6638 16192 6644 16204
rect 6696 16192 6702 16244
rect 7101 16235 7159 16241
rect 7101 16201 7113 16235
rect 7147 16232 7159 16235
rect 8202 16232 8208 16244
rect 7147 16204 8208 16232
rect 7147 16201 7159 16204
rect 7101 16195 7159 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9582 16232 9588 16244
rect 9543 16204 9588 16232
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 10134 16232 10140 16244
rect 10095 16204 10140 16232
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10502 16232 10508 16244
rect 10463 16204 10508 16232
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10778 16232 10784 16244
rect 10739 16204 10784 16232
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11790 16232 11796 16244
rect 11751 16204 11796 16232
rect 11790 16192 11796 16204
rect 11848 16232 11854 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 11848 16204 12173 16232
rect 11848 16192 11854 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 7742 16164 7748 16176
rect 7703 16136 7748 16164
rect 7742 16124 7748 16136
rect 7800 16124 7806 16176
rect 8018 16164 8024 16176
rect 7979 16136 8024 16164
rect 8018 16124 8024 16136
rect 8076 16124 8082 16176
rect 12176 16164 12204 16195
rect 12434 16192 12440 16244
rect 12492 16232 12498 16244
rect 12986 16232 12992 16244
rect 12492 16204 12992 16232
rect 12492 16192 12498 16204
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14366 16232 14372 16244
rect 14047 16204 14372 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 15381 16235 15439 16241
rect 15381 16201 15393 16235
rect 15427 16232 15439 16235
rect 15838 16232 15844 16244
rect 15427 16204 15844 16232
rect 15427 16201 15439 16204
rect 15381 16195 15439 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 16393 16235 16451 16241
rect 16393 16201 16405 16235
rect 16439 16232 16451 16235
rect 16482 16232 16488 16244
rect 16439 16204 16488 16232
rect 16439 16201 16451 16204
rect 16393 16195 16451 16201
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 18380 16204 19441 16232
rect 18380 16192 18386 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 20625 16235 20683 16241
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 20714 16232 20720 16244
rect 20671 16204 20720 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 20898 16232 20904 16244
rect 20859 16204 20904 16232
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 23750 16232 23756 16244
rect 23711 16204 23756 16232
rect 23750 16192 23756 16204
rect 23808 16192 23814 16244
rect 25498 16232 25504 16244
rect 25459 16204 25504 16232
rect 25498 16192 25504 16204
rect 25556 16192 25562 16244
rect 12176 16136 13124 16164
rect 13096 16108 13124 16136
rect 19334 16124 19340 16176
rect 19392 16164 19398 16176
rect 19981 16167 20039 16173
rect 19981 16164 19993 16167
rect 19392 16136 19993 16164
rect 19392 16124 19398 16136
rect 19981 16133 19993 16136
rect 20027 16133 20039 16167
rect 19981 16127 20039 16133
rect 3234 16096 3240 16108
rect 3195 16068 3240 16096
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 3421 16099 3479 16105
rect 3421 16065 3433 16099
rect 3467 16096 3479 16099
rect 3510 16096 3516 16108
rect 3467 16068 3516 16096
rect 3467 16065 3479 16068
rect 3421 16059 3479 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 4264 16068 5733 16096
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1854 16028 1860 16040
rect 1443 16000 1860 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 1854 15988 1860 16000
rect 1912 16028 1918 16040
rect 1912 16000 2728 16028
rect 1912 15988 1918 16000
rect 1670 15960 1676 15972
rect 1631 15932 1676 15960
rect 1670 15920 1676 15932
rect 1728 15920 1734 15972
rect 2222 15960 2228 15972
rect 2135 15932 2228 15960
rect 2222 15920 2228 15932
rect 2280 15960 2286 15972
rect 2700 15960 2728 16000
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 2924 16000 3157 16028
rect 2924 15988 2930 16000
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3145 15991 3203 15997
rect 3789 15963 3847 15969
rect 3789 15960 3801 15963
rect 2280 15932 2636 15960
rect 2700 15932 3801 15960
rect 2280 15920 2286 15932
rect 2608 15892 2636 15932
rect 3789 15929 3801 15932
rect 3835 15929 3847 15963
rect 3789 15923 3847 15929
rect 4264 15901 4292 16068
rect 5721 16065 5733 16068
rect 5767 16096 5779 16099
rect 6086 16096 6092 16108
rect 5767 16068 6092 16096
rect 5767 16065 5779 16068
rect 5721 16059 5779 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16096 7251 16099
rect 7466 16096 7472 16108
rect 7239 16068 7472 16096
rect 7239 16065 7251 16068
rect 7193 16059 7251 16065
rect 7466 16056 7472 16068
rect 7524 16056 7530 16108
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8205 16099 8263 16105
rect 8205 16096 8217 16099
rect 8168 16068 8217 16096
rect 8168 16056 8174 16068
rect 8205 16065 8217 16068
rect 8251 16065 8263 16099
rect 11422 16096 11428 16108
rect 11383 16068 11428 16096
rect 8205 16059 8263 16065
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 12897 16099 12955 16105
rect 12897 16096 12909 16099
rect 12860 16068 12909 16096
rect 12860 16056 12866 16068
rect 12897 16065 12909 16068
rect 12943 16065 12955 16099
rect 13078 16096 13084 16108
rect 13039 16068 13084 16096
rect 12897 16059 12955 16065
rect 13078 16056 13084 16068
rect 13136 16056 13142 16108
rect 14090 16096 14096 16108
rect 13832 16068 14096 16096
rect 4982 15988 4988 16040
rect 5040 16028 5046 16040
rect 5629 16031 5687 16037
rect 5629 16028 5641 16031
rect 5040 16000 5641 16028
rect 5040 15988 5046 16000
rect 5629 15997 5641 16000
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 8472 16031 8530 16037
rect 8472 15997 8484 16031
rect 8518 16028 8530 16031
rect 9490 16028 9496 16040
rect 8518 16000 9496 16028
rect 8518 15997 8530 16000
rect 8472 15991 8530 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 4709 15963 4767 15969
rect 4709 15929 4721 15963
rect 4755 15960 4767 15963
rect 5537 15963 5595 15969
rect 5537 15960 5549 15963
rect 4755 15932 5549 15960
rect 4755 15929 4767 15932
rect 4709 15923 4767 15929
rect 5537 15929 5549 15932
rect 5583 15960 5595 15963
rect 6822 15960 6828 15972
rect 5583 15932 6828 15960
rect 5583 15929 5595 15932
rect 5537 15923 5595 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 10778 15920 10784 15972
rect 10836 15960 10842 15972
rect 11241 15963 11299 15969
rect 11241 15960 11253 15963
rect 10836 15932 11253 15960
rect 10836 15920 10842 15932
rect 11241 15929 11253 15932
rect 11287 15960 11299 15963
rect 11287 15932 12480 15960
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 4249 15895 4307 15901
rect 4249 15892 4261 15895
rect 2608 15864 4261 15892
rect 4249 15861 4261 15864
rect 4295 15861 4307 15895
rect 4982 15892 4988 15904
rect 4943 15864 4988 15892
rect 4249 15855 4307 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 11146 15892 11152 15904
rect 11059 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15892 11210 15904
rect 12250 15892 12256 15904
rect 11204 15864 12256 15892
rect 11204 15852 11210 15864
rect 12250 15852 12256 15864
rect 12308 15852 12314 15904
rect 12452 15901 12480 15932
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15861 12495 15895
rect 12802 15892 12808 15904
rect 12715 15864 12808 15892
rect 12437 15855 12495 15861
rect 12802 15852 12808 15864
rect 12860 15892 12866 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12860 15864 13461 15892
rect 12860 15852 12866 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 13832 15901 13860 16068
rect 14090 16056 14096 16068
rect 14148 16096 14154 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14148 16068 14565 16096
rect 14148 16056 14154 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16096 15991 16099
rect 17037 16099 17095 16105
rect 17037 16096 17049 16099
rect 15979 16068 17049 16096
rect 15979 16065 15991 16068
rect 15933 16059 15991 16065
rect 17037 16065 17049 16068
rect 17083 16096 17095 16099
rect 17494 16096 17500 16108
rect 17083 16068 17500 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 17865 16099 17923 16105
rect 17865 16065 17877 16099
rect 17911 16096 17923 16099
rect 20916 16096 20944 16192
rect 17911 16068 18184 16096
rect 20916 16068 21220 16096
rect 17911 16065 17923 16068
rect 17865 16059 17923 16065
rect 16574 15988 16580 16040
rect 16632 16028 16638 16040
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 16632 16000 16773 16028
rect 16632 15988 16638 16000
rect 16761 15997 16773 16000
rect 16807 16028 16819 16031
rect 17402 16028 17408 16040
rect 16807 16000 17408 16028
rect 16807 15997 16819 16000
rect 16761 15991 16819 15997
rect 17402 15988 17408 16000
rect 17460 15988 17466 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18156 16028 18184 16068
rect 18316 16031 18374 16037
rect 18316 16028 18328 16031
rect 18156 16000 18328 16028
rect 18316 15997 18328 16000
rect 18362 16028 18374 16031
rect 18690 16028 18696 16040
rect 18362 16000 18696 16028
rect 18362 15997 18374 16000
rect 18316 15991 18374 15997
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 21085 16031 21143 16037
rect 21085 16028 21097 16031
rect 20772 16000 21097 16028
rect 20772 15988 20778 16000
rect 21085 15997 21097 16000
rect 21131 15997 21143 16031
rect 21192 16028 21220 16068
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22830 16096 22836 16108
rect 22520 16068 22836 16096
rect 22520 16056 22526 16068
rect 22830 16056 22836 16068
rect 22888 16056 22894 16108
rect 24026 16056 24032 16108
rect 24084 16096 24090 16108
rect 24305 16099 24363 16105
rect 24305 16096 24317 16099
rect 24084 16068 24317 16096
rect 24084 16056 24090 16068
rect 24305 16065 24317 16068
rect 24351 16096 24363 16099
rect 24762 16096 24768 16108
rect 24351 16068 24768 16096
rect 24351 16065 24363 16068
rect 24305 16059 24363 16065
rect 24762 16056 24768 16068
rect 24820 16096 24826 16108
rect 25133 16099 25191 16105
rect 25133 16096 25145 16099
rect 24820 16068 25145 16096
rect 24820 16056 24826 16068
rect 25133 16065 25145 16068
rect 25179 16065 25191 16099
rect 25133 16059 25191 16065
rect 21341 16031 21399 16037
rect 21341 16028 21353 16031
rect 21192 16000 21353 16028
rect 21085 15991 21143 15997
rect 21341 15997 21353 16000
rect 21387 15997 21399 16031
rect 21341 15991 21399 15997
rect 25222 15988 25228 16040
rect 25280 16028 25286 16040
rect 25317 16031 25375 16037
rect 25317 16028 25329 16031
rect 25280 16000 25329 16028
rect 25280 15988 25286 16000
rect 25317 15997 25329 16000
rect 25363 16028 25375 16031
rect 25869 16031 25927 16037
rect 25869 16028 25881 16031
rect 25363 16000 25881 16028
rect 25363 15997 25375 16000
rect 25317 15991 25375 15997
rect 25869 15997 25881 16000
rect 25915 15997 25927 16031
rect 25869 15991 25927 15997
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 16850 15960 16856 15972
rect 16347 15932 16856 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 22830 15920 22836 15972
rect 22888 15960 22894 15972
rect 23017 15963 23075 15969
rect 23017 15960 23029 15963
rect 22888 15932 23029 15960
rect 22888 15920 22894 15932
rect 23017 15929 23029 15932
rect 23063 15960 23075 15963
rect 24121 15963 24179 15969
rect 24121 15960 24133 15963
rect 23063 15932 24133 15960
rect 23063 15929 23075 15932
rect 23017 15923 23075 15929
rect 24121 15929 24133 15932
rect 24167 15929 24179 15963
rect 24121 15923 24179 15929
rect 13817 15895 13875 15901
rect 13817 15892 13829 15895
rect 13688 15864 13829 15892
rect 13688 15852 13694 15864
rect 13817 15861 13829 15864
rect 13863 15861 13875 15895
rect 13817 15855 13875 15861
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14369 15895 14427 15901
rect 14369 15892 14381 15895
rect 14240 15864 14381 15892
rect 14240 15852 14246 15864
rect 14369 15861 14381 15864
rect 14415 15861 14427 15895
rect 14369 15855 14427 15861
rect 14458 15852 14464 15904
rect 14516 15892 14522 15904
rect 17494 15892 17500 15904
rect 14516 15864 14561 15892
rect 17455 15864 17500 15892
rect 14516 15852 14522 15864
rect 17494 15852 17500 15864
rect 17552 15852 17558 15904
rect 22465 15895 22523 15901
rect 22465 15861 22477 15895
rect 22511 15892 22523 15895
rect 22922 15892 22928 15904
rect 22511 15864 22928 15892
rect 22511 15861 22523 15864
rect 22465 15855 22523 15861
rect 22922 15852 22928 15864
rect 22980 15852 22986 15904
rect 23474 15892 23480 15904
rect 23387 15864 23480 15892
rect 23474 15852 23480 15864
rect 23532 15892 23538 15904
rect 24213 15895 24271 15901
rect 24213 15892 24225 15895
rect 23532 15864 24225 15892
rect 23532 15852 23538 15864
rect 24213 15861 24225 15864
rect 24259 15892 24271 15895
rect 25498 15892 25504 15904
rect 24259 15864 25504 15892
rect 24259 15861 24271 15864
rect 24213 15855 24271 15861
rect 25498 15852 25504 15864
rect 25556 15852 25562 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 3292 15660 3525 15688
rect 3292 15648 3298 15660
rect 3513 15657 3525 15660
rect 3559 15657 3571 15691
rect 3513 15651 3571 15657
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 4028 15660 4261 15688
rect 4028 15648 4034 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 4249 15651 4307 15657
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 4488 15660 4997 15688
rect 4488 15648 4494 15660
rect 4985 15657 4997 15660
rect 5031 15657 5043 15691
rect 4985 15651 5043 15657
rect 5442 15648 5448 15700
rect 5500 15688 5506 15700
rect 5997 15691 6055 15697
rect 5997 15688 6009 15691
rect 5500 15660 6009 15688
rect 5500 15648 5506 15660
rect 5997 15657 6009 15660
rect 6043 15688 6055 15691
rect 6730 15688 6736 15700
rect 6043 15660 6736 15688
rect 6043 15657 6055 15660
rect 5997 15651 6055 15657
rect 6730 15648 6736 15660
rect 6788 15648 6794 15700
rect 9125 15691 9183 15697
rect 9125 15657 9137 15691
rect 9171 15688 9183 15691
rect 9490 15688 9496 15700
rect 9171 15660 9496 15688
rect 9171 15657 9183 15660
rect 9125 15651 9183 15657
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9858 15688 9864 15700
rect 9819 15660 9864 15688
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10192 15660 10333 15688
rect 10192 15648 10198 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10778 15688 10784 15700
rect 10739 15660 10784 15688
rect 10321 15651 10379 15657
rect 10778 15648 10784 15660
rect 10836 15648 10842 15700
rect 12894 15688 12900 15700
rect 12855 15660 12900 15688
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 13998 15648 14004 15700
rect 14056 15688 14062 15700
rect 14737 15691 14795 15697
rect 14737 15688 14749 15691
rect 14056 15660 14749 15688
rect 14056 15648 14062 15660
rect 14737 15657 14749 15660
rect 14783 15657 14795 15691
rect 18230 15688 18236 15700
rect 18191 15660 18236 15688
rect 14737 15651 14795 15657
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15688 20959 15691
rect 21082 15688 21088 15700
rect 20947 15660 21088 15688
rect 20947 15657 20959 15660
rect 20901 15651 20959 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 22278 15688 22284 15700
rect 22239 15660 22284 15688
rect 22278 15648 22284 15660
rect 22336 15648 22342 15700
rect 24762 15688 24768 15700
rect 24723 15660 24768 15688
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 6546 15620 6552 15632
rect 5368 15592 6552 15620
rect 2314 15552 2320 15564
rect 2275 15524 2320 15552
rect 2314 15512 2320 15524
rect 2372 15512 2378 15564
rect 3970 15512 3976 15564
rect 4028 15552 4034 15564
rect 5368 15561 5396 15592
rect 6546 15580 6552 15592
rect 6604 15580 6610 15632
rect 7368 15623 7426 15629
rect 7368 15589 7380 15623
rect 7414 15620 7426 15623
rect 7926 15620 7932 15632
rect 7414 15592 7932 15620
rect 7414 15589 7426 15592
rect 7368 15583 7426 15589
rect 7926 15580 7932 15592
rect 7984 15580 7990 15632
rect 11054 15580 11060 15632
rect 11112 15629 11118 15632
rect 11112 15623 11176 15629
rect 11112 15589 11130 15623
rect 11164 15589 11176 15623
rect 11112 15583 11176 15589
rect 18141 15623 18199 15629
rect 18141 15589 18153 15623
rect 18187 15620 18199 15623
rect 18322 15620 18328 15632
rect 18187 15592 18328 15620
rect 18187 15589 18199 15592
rect 18141 15583 18199 15589
rect 11112 15580 11118 15583
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 22922 15580 22928 15632
rect 22980 15620 22986 15632
rect 23630 15623 23688 15629
rect 23630 15620 23642 15623
rect 22980 15592 23642 15620
rect 22980 15580 22986 15592
rect 23630 15589 23642 15592
rect 23676 15620 23688 15623
rect 24026 15620 24032 15632
rect 23676 15592 24032 15620
rect 23676 15589 23688 15592
rect 23630 15583 23688 15589
rect 24026 15580 24032 15592
rect 24084 15580 24090 15632
rect 4065 15555 4123 15561
rect 4065 15552 4077 15555
rect 4028 15524 4077 15552
rect 4028 15512 4034 15524
rect 4065 15521 4077 15524
rect 4111 15521 4123 15555
rect 4065 15515 4123 15521
rect 5353 15555 5411 15561
rect 5353 15521 5365 15555
rect 5399 15521 5411 15555
rect 5353 15515 5411 15521
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5592 15524 5917 15552
rect 5592 15512 5598 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 7101 15555 7159 15561
rect 7101 15521 7113 15555
rect 7147 15552 7159 15555
rect 8110 15552 8116 15564
rect 7147 15524 8116 15552
rect 7147 15521 7159 15524
rect 7101 15515 7159 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9490 15552 9496 15564
rect 9451 15524 9496 15552
rect 9490 15512 9496 15524
rect 9548 15512 9554 15564
rect 13722 15552 13728 15564
rect 13683 15524 13728 15552
rect 13722 15512 13728 15524
rect 13780 15512 13786 15564
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 16016 15555 16074 15561
rect 16016 15552 16028 15555
rect 15703 15524 16028 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 16016 15521 16028 15524
rect 16062 15552 16074 15555
rect 16298 15552 16304 15564
rect 16062 15524 16304 15552
rect 16062 15521 16074 15524
rect 16016 15515 16074 15521
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18601 15555 18659 15561
rect 18601 15552 18613 15555
rect 18012 15524 18613 15552
rect 18012 15512 18018 15524
rect 18601 15521 18613 15524
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15552 20775 15555
rect 20898 15552 20904 15564
rect 20763 15524 20904 15552
rect 20763 15521 20775 15524
rect 20717 15515 20775 15521
rect 20898 15512 20904 15524
rect 20956 15552 20962 15564
rect 21269 15555 21327 15561
rect 21269 15552 21281 15555
rect 20956 15524 21281 15552
rect 20956 15512 20962 15524
rect 21269 15521 21281 15524
rect 21315 15521 21327 15555
rect 22646 15552 22652 15564
rect 22607 15524 22652 15552
rect 21269 15515 21327 15521
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 2406 15484 2412 15496
rect 2367 15456 2412 15484
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 6086 15484 6092 15496
rect 2556 15456 2601 15484
rect 6047 15456 6092 15484
rect 2556 15444 2562 15456
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 9674 15444 9680 15496
rect 9732 15484 9738 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 9732 15456 10885 15484
rect 9732 15444 9738 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 13814 15484 13820 15496
rect 13775 15456 13820 15484
rect 10873 15447 10931 15453
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 13906 15444 13912 15496
rect 13964 15484 13970 15496
rect 14369 15487 14427 15493
rect 14369 15484 14381 15487
rect 13964 15456 14381 15484
rect 13964 15444 13970 15456
rect 14369 15453 14381 15456
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15453 15807 15487
rect 18690 15484 18696 15496
rect 18651 15456 18696 15484
rect 15749 15447 15807 15453
rect 1946 15376 1952 15428
rect 2004 15416 2010 15428
rect 4617 15419 4675 15425
rect 4617 15416 4629 15419
rect 2004 15388 4629 15416
rect 2004 15376 2010 15388
rect 4617 15385 4629 15388
rect 4663 15385 4675 15419
rect 4617 15379 4675 15385
rect 5537 15419 5595 15425
rect 5537 15385 5549 15419
rect 5583 15416 5595 15419
rect 7006 15416 7012 15428
rect 5583 15388 7012 15416
rect 5583 15385 5595 15388
rect 5537 15379 5595 15385
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 12253 15419 12311 15425
rect 12253 15385 12265 15419
rect 12299 15416 12311 15419
rect 13078 15416 13084 15428
rect 12299 15388 13084 15416
rect 12299 15385 12311 15388
rect 12253 15379 12311 15385
rect 13078 15376 13084 15388
rect 13136 15376 13142 15428
rect 1673 15351 1731 15357
rect 1673 15317 1685 15351
rect 1719 15348 1731 15351
rect 2038 15348 2044 15360
rect 1719 15320 2044 15348
rect 1719 15317 1731 15320
rect 1673 15311 1731 15317
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 3234 15348 3240 15360
rect 3195 15320 3240 15348
rect 3234 15308 3240 15320
rect 3292 15308 3298 15360
rect 3694 15308 3700 15360
rect 3752 15348 3758 15360
rect 4154 15348 4160 15360
rect 3752 15320 4160 15348
rect 3752 15308 3758 15320
rect 4154 15308 4160 15320
rect 4212 15308 4218 15360
rect 5169 15351 5227 15357
rect 5169 15317 5181 15351
rect 5215 15348 5227 15351
rect 5350 15348 5356 15360
rect 5215 15320 5356 15348
rect 5215 15317 5227 15320
rect 5169 15311 5227 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15348 6975 15351
rect 7282 15348 7288 15360
rect 6963 15320 7288 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8481 15351 8539 15357
rect 8481 15348 8493 15351
rect 8352 15320 8493 15348
rect 8352 15308 8358 15320
rect 8481 15317 8493 15320
rect 8527 15317 8539 15351
rect 13170 15348 13176 15360
rect 13131 15320 13176 15348
rect 8481 15311 8539 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 15764 15348 15792 15447
rect 18690 15444 18696 15456
rect 18748 15444 18754 15496
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 18966 15484 18972 15496
rect 18923 15456 18972 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 17129 15419 17187 15425
rect 17129 15385 17141 15419
rect 17175 15416 17187 15419
rect 17494 15416 17500 15428
rect 17175 15388 17500 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17494 15376 17500 15388
rect 17552 15416 17558 15428
rect 18892 15416 18920 15447
rect 18966 15444 18972 15456
rect 19024 15444 19030 15496
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 20346 15484 20352 15496
rect 19843 15456 20352 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 21358 15484 21364 15496
rect 21319 15456 21364 15484
rect 21358 15444 21364 15456
rect 21416 15444 21422 15496
rect 21545 15487 21603 15493
rect 21545 15453 21557 15487
rect 21591 15484 21603 15487
rect 21818 15484 21824 15496
rect 21591 15456 21824 15484
rect 21591 15453 21603 15456
rect 21545 15447 21603 15453
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 23308 15456 23397 15484
rect 17552 15388 18920 15416
rect 17552 15376 17558 15388
rect 23308 15360 23336 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 16114 15348 16120 15360
rect 15764 15320 16120 15348
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16482 15308 16488 15360
rect 16540 15348 16546 15360
rect 17586 15348 17592 15360
rect 16540 15320 17592 15348
rect 16540 15308 16546 15320
rect 17586 15308 17592 15320
rect 17644 15348 17650 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 17644 15320 17693 15348
rect 17644 15308 17650 15320
rect 17681 15317 17693 15320
rect 17727 15348 17739 15351
rect 17770 15348 17776 15360
rect 17727 15320 17776 15348
rect 17727 15317 17739 15320
rect 17681 15311 17739 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 19334 15348 19340 15360
rect 19295 15320 19340 15348
rect 19334 15308 19340 15320
rect 19392 15348 19398 15360
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19392 15320 19625 15348
rect 19392 15308 19398 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15348 20407 15351
rect 20714 15348 20720 15360
rect 20395 15320 20720 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 20714 15308 20720 15320
rect 20772 15348 20778 15360
rect 21913 15351 21971 15357
rect 21913 15348 21925 15351
rect 20772 15320 21925 15348
rect 20772 15308 20778 15320
rect 21913 15317 21925 15320
rect 21959 15348 21971 15351
rect 22465 15351 22523 15357
rect 22465 15348 22477 15351
rect 21959 15320 22477 15348
rect 21959 15317 21971 15320
rect 21913 15311 21971 15317
rect 22465 15317 22477 15320
rect 22511 15348 22523 15351
rect 23290 15348 23296 15360
rect 22511 15320 23296 15348
rect 22511 15317 22523 15320
rect 22465 15311 22523 15317
rect 23290 15308 23296 15320
rect 23348 15308 23354 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 3053 15147 3111 15153
rect 3053 15113 3065 15147
rect 3099 15144 3111 15147
rect 4338 15144 4344 15156
rect 3099 15116 4344 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 1946 15036 1952 15088
rect 2004 15076 2010 15088
rect 2406 15076 2412 15088
rect 2004 15048 2412 15076
rect 2004 15036 2010 15048
rect 2406 15036 2412 15048
rect 2464 15076 2470 15088
rect 2593 15079 2651 15085
rect 2593 15076 2605 15079
rect 2464 15048 2605 15076
rect 2464 15036 2470 15048
rect 2593 15045 2605 15048
rect 2639 15045 2651 15079
rect 2593 15039 2651 15045
rect 2869 15079 2927 15085
rect 2869 15045 2881 15079
rect 2915 15076 2927 15079
rect 3068 15076 3096 15107
rect 4338 15104 4344 15116
rect 4396 15144 4402 15156
rect 5074 15144 5080 15156
rect 4396 15116 5080 15144
rect 4396 15104 4402 15116
rect 5074 15104 5080 15116
rect 5132 15104 5138 15156
rect 5169 15147 5227 15153
rect 5169 15113 5181 15147
rect 5215 15144 5227 15147
rect 5258 15144 5264 15156
rect 5215 15116 5264 15144
rect 5215 15113 5227 15116
rect 5169 15107 5227 15113
rect 5258 15104 5264 15116
rect 5316 15104 5322 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 7926 15144 7932 15156
rect 7887 15116 7932 15144
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 8849 15147 8907 15153
rect 8849 15144 8861 15147
rect 8168 15116 8861 15144
rect 8168 15104 8174 15116
rect 8849 15113 8861 15116
rect 8895 15113 8907 15147
rect 8849 15107 8907 15113
rect 10965 15147 11023 15153
rect 10965 15113 10977 15147
rect 11011 15144 11023 15147
rect 11054 15144 11060 15156
rect 11011 15116 11060 15144
rect 11011 15113 11023 15116
rect 10965 15107 11023 15113
rect 2915 15048 3096 15076
rect 2915 15045 2927 15048
rect 2869 15039 2927 15045
rect 4246 15036 4252 15088
rect 4304 15076 4310 15088
rect 4525 15079 4583 15085
rect 4525 15076 4537 15079
rect 4304 15048 4537 15076
rect 4304 15036 4310 15048
rect 4525 15045 4537 15048
rect 4571 15076 4583 15079
rect 6270 15076 6276 15088
rect 4571 15048 6276 15076
rect 4571 15045 4583 15048
rect 4525 15039 4583 15045
rect 6270 15036 6276 15048
rect 6328 15036 6334 15088
rect 2222 15008 2228 15020
rect 2183 14980 2228 15008
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 6144 14980 7389 15008
rect 6144 14968 6150 14980
rect 7377 14977 7389 14980
rect 7423 15008 7435 15011
rect 7558 15008 7564 15020
rect 7423 14980 7564 15008
rect 7423 14977 7435 14980
rect 7377 14971 7435 14977
rect 7558 14968 7564 14980
rect 7616 15008 7622 15020
rect 8202 15008 8208 15020
rect 7616 14980 8208 15008
rect 7616 14968 7622 14980
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8389 15011 8447 15017
rect 8389 14977 8401 15011
rect 8435 15008 8447 15011
rect 8478 15008 8484 15020
rect 8435 14980 8484 15008
rect 8435 14977 8447 14980
rect 8389 14971 8447 14977
rect 8478 14968 8484 14980
rect 8536 14968 8542 15020
rect 3050 14900 3056 14952
rect 3108 14940 3114 14952
rect 3145 14943 3203 14949
rect 3145 14940 3157 14943
rect 3108 14912 3157 14940
rect 3108 14900 3114 14912
rect 3145 14909 3157 14912
rect 3191 14909 3203 14943
rect 3145 14903 3203 14909
rect 5629 14943 5687 14949
rect 5629 14909 5641 14943
rect 5675 14909 5687 14943
rect 6638 14940 6644 14952
rect 6551 14912 6644 14940
rect 5629 14903 5687 14909
rect 1949 14875 2007 14881
rect 1949 14841 1961 14875
rect 1995 14872 2007 14875
rect 1995 14844 2728 14872
rect 1995 14841 2007 14844
rect 1949 14835 2007 14841
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 2700 14804 2728 14844
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 3234 14872 3240 14884
rect 2832 14844 3240 14872
rect 2832 14832 2838 14844
rect 3234 14832 3240 14844
rect 3292 14872 3298 14884
rect 3390 14875 3448 14881
rect 3390 14872 3402 14875
rect 3292 14844 3402 14872
rect 3292 14832 3298 14844
rect 3390 14841 3402 14844
rect 3436 14841 3448 14875
rect 5644 14872 5672 14903
rect 6638 14900 6644 14912
rect 6696 14940 6702 14952
rect 7190 14940 7196 14952
rect 6696 14912 7196 14940
rect 6696 14900 6702 14912
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 8864 14940 8892 15107
rect 11054 15104 11060 15116
rect 11112 15144 11118 15156
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11112 15116 11805 15144
rect 11112 15104 11118 15116
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 12437 15147 12495 15153
rect 12437 15113 12449 15147
rect 12483 15144 12495 15147
rect 12802 15144 12808 15156
rect 12483 15116 12808 15144
rect 12483 15113 12495 15116
rect 12437 15107 12495 15113
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 11808 15008 11836 15107
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 13541 15147 13599 15153
rect 13541 15113 13553 15147
rect 13587 15144 13599 15147
rect 13722 15144 13728 15156
rect 13587 15116 13728 15144
rect 13587 15113 13599 15116
rect 13541 15107 13599 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 14700 15116 15945 15144
rect 14700 15104 14706 15116
rect 15933 15113 15945 15116
rect 15979 15144 15991 15147
rect 17862 15144 17868 15156
rect 15979 15116 16896 15144
rect 17823 15116 17868 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 13170 15036 13176 15088
rect 13228 15076 13234 15088
rect 14001 15079 14059 15085
rect 14001 15076 14013 15079
rect 13228 15048 14013 15076
rect 13228 15036 13234 15048
rect 14001 15045 14013 15048
rect 14047 15045 14059 15079
rect 14001 15039 14059 15045
rect 16868 15076 16896 15116
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 20346 15144 20352 15156
rect 20307 15116 20352 15144
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20898 15144 20904 15156
rect 20859 15116 20904 15144
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 21818 15104 21824 15156
rect 21876 15144 21882 15156
rect 21913 15147 21971 15153
rect 21913 15144 21925 15147
rect 21876 15116 21925 15144
rect 21876 15104 21882 15116
rect 21913 15113 21925 15116
rect 21959 15113 21971 15147
rect 21913 15107 21971 15113
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22649 15147 22707 15153
rect 22152 15116 22324 15144
rect 22152 15104 22158 15116
rect 17310 15076 17316 15088
rect 16868 15048 17316 15076
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 9539 14980 9720 15008
rect 11808 14980 13001 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 9582 14940 9588 14952
rect 8812 14912 9588 14940
rect 8812 14900 8818 14912
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9692 14940 9720 14980
rect 12989 14977 13001 14980
rect 13035 15008 13047 15011
rect 13906 15008 13912 15020
rect 13035 14980 13912 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13906 14968 13912 14980
rect 13964 15008 13970 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 13964 14980 14565 15008
rect 13964 14968 13970 14980
rect 14553 14977 14565 14980
rect 14599 15008 14611 15011
rect 15013 15011 15071 15017
rect 15013 15008 15025 15011
rect 14599 14980 15025 15008
rect 14599 14977 14611 14980
rect 14553 14971 14611 14977
rect 15013 14977 15025 14980
rect 15059 14977 15071 15011
rect 15654 15008 15660 15020
rect 15567 14980 15660 15008
rect 15013 14971 15071 14977
rect 15654 14968 15660 14980
rect 15712 15008 15718 15020
rect 16868 15017 16896 15048
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 16853 15011 16911 15017
rect 15712 14980 16804 15008
rect 15712 14968 15718 14980
rect 16776 14952 16804 14980
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 16853 14971 16911 14977
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20530 15008 20536 15020
rect 20119 14980 20536 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 20530 14968 20536 14980
rect 20588 15008 20594 15020
rect 21453 15011 21511 15017
rect 21453 15008 21465 15011
rect 20588 14980 21465 15008
rect 20588 14968 20594 14980
rect 21453 14977 21465 14980
rect 21499 15008 21511 15011
rect 22094 15008 22100 15020
rect 21499 14980 22100 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 22094 14968 22100 14980
rect 22152 14968 22158 15020
rect 9852 14943 9910 14949
rect 9852 14940 9864 14943
rect 9692 14912 9864 14940
rect 9852 14909 9864 14912
rect 9898 14940 9910 14943
rect 10134 14940 10140 14952
rect 9898 14912 10140 14940
rect 9898 14909 9910 14912
rect 9852 14903 9910 14909
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 12253 14943 12311 14949
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12526 14940 12532 14952
rect 12299 14912 12532 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12526 14900 12532 14912
rect 12584 14940 12590 14952
rect 12894 14940 12900 14952
rect 12584 14912 12900 14940
rect 12584 14900 12590 14912
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 15930 14900 15936 14952
rect 15988 14940 15994 14952
rect 16301 14943 16359 14949
rect 16301 14940 16313 14943
rect 15988 14912 16313 14940
rect 15988 14900 15994 14912
rect 16301 14909 16313 14912
rect 16347 14940 16359 14943
rect 16482 14940 16488 14952
rect 16347 14912 16488 14940
rect 16347 14909 16359 14912
rect 16301 14903 16359 14909
rect 16482 14900 16488 14912
rect 16540 14900 16546 14952
rect 16758 14940 16764 14952
rect 16719 14912 16764 14940
rect 16758 14900 16764 14912
rect 16816 14900 16822 14952
rect 18046 14940 18052 14952
rect 18007 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 18322 14949 18328 14952
rect 18316 14940 18328 14949
rect 18283 14912 18328 14940
rect 18316 14903 18328 14912
rect 18322 14900 18328 14903
rect 18380 14900 18386 14952
rect 20346 14900 20352 14952
rect 20404 14940 20410 14952
rect 21269 14943 21327 14949
rect 21269 14940 21281 14943
rect 20404 14912 21281 14940
rect 20404 14900 20410 14912
rect 21269 14909 21281 14912
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 6273 14875 6331 14881
rect 6273 14872 6285 14875
rect 5644 14844 6285 14872
rect 3390 14835 3448 14841
rect 6273 14841 6285 14844
rect 6319 14872 6331 14875
rect 6319 14844 7328 14872
rect 6319 14841 6331 14844
rect 6273 14835 6331 14841
rect 7300 14816 7328 14844
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 13817 14875 13875 14881
rect 13817 14872 13829 14875
rect 12032 14844 13829 14872
rect 12032 14832 12038 14844
rect 13817 14841 13829 14844
rect 13863 14872 13875 14875
rect 14461 14875 14519 14881
rect 14461 14872 14473 14875
rect 13863 14844 14473 14872
rect 13863 14841 13875 14844
rect 13817 14835 13875 14841
rect 14461 14841 14473 14844
rect 14507 14872 14519 14875
rect 15286 14872 15292 14884
rect 14507 14844 15292 14872
rect 14507 14841 14519 14844
rect 14461 14835 14519 14841
rect 15286 14832 15292 14844
rect 15344 14832 15350 14884
rect 17954 14872 17960 14884
rect 17420 14844 17960 14872
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2700 14776 2881 14804
rect 2869 14773 2881 14776
rect 2915 14773 2927 14807
rect 5810 14804 5816 14816
rect 5771 14776 5816 14804
rect 2869 14767 2927 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14804 6883 14807
rect 6914 14804 6920 14816
rect 6871 14776 6920 14804
rect 6871 14773 6883 14776
rect 6825 14767 6883 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7282 14804 7288 14816
rect 7243 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 8202 14804 8208 14816
rect 8163 14776 8208 14804
rect 8202 14764 8208 14776
rect 8260 14764 8266 14816
rect 12802 14804 12808 14816
rect 12763 14776 12808 14804
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 14090 14764 14096 14816
rect 14148 14804 14154 14816
rect 14369 14807 14427 14813
rect 14369 14804 14381 14807
rect 14148 14776 14381 14804
rect 14148 14764 14154 14776
rect 14369 14773 14381 14776
rect 14415 14773 14427 14807
rect 16114 14804 16120 14816
rect 16075 14776 16120 14804
rect 14369 14767 14427 14773
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 16393 14807 16451 14813
rect 16393 14773 16405 14807
rect 16439 14804 16451 14807
rect 16666 14804 16672 14816
rect 16439 14776 16672 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16666 14764 16672 14776
rect 16724 14764 16730 14816
rect 16942 14764 16948 14816
rect 17000 14804 17006 14816
rect 17420 14813 17448 14844
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 22296 14872 22324 15116
rect 22649 15113 22661 15147
rect 22695 15144 22707 15147
rect 22738 15144 22744 15156
rect 22695 15116 22744 15144
rect 22695 15113 22707 15116
rect 22649 15107 22707 15113
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 22922 15104 22928 15156
rect 22980 15144 22986 15156
rect 23017 15147 23075 15153
rect 23017 15144 23029 15147
rect 22980 15116 23029 15144
rect 22980 15104 22986 15116
rect 23017 15113 23029 15116
rect 23063 15113 23075 15147
rect 23017 15107 23075 15113
rect 23753 15147 23811 15153
rect 23753 15113 23765 15147
rect 23799 15144 23811 15147
rect 24118 15144 24124 15156
rect 23799 15116 24124 15144
rect 23799 15113 23811 15116
rect 23753 15107 23811 15113
rect 24118 15104 24124 15116
rect 24176 15104 24182 15156
rect 24762 15144 24768 15156
rect 24723 15116 24768 15144
rect 24762 15104 24768 15116
rect 24820 15104 24826 15156
rect 25406 15104 25412 15156
rect 25464 15144 25470 15156
rect 25501 15147 25559 15153
rect 25501 15144 25513 15147
rect 25464 15116 25513 15144
rect 25464 15104 25470 15116
rect 25501 15113 25513 15116
rect 25547 15113 25559 15147
rect 25501 15107 25559 15113
rect 22373 15079 22431 15085
rect 22373 15045 22385 15079
rect 22419 15076 22431 15079
rect 23198 15076 23204 15088
rect 22419 15048 23204 15076
rect 22419 15045 22431 15048
rect 22373 15039 22431 15045
rect 22480 14949 22508 15048
rect 23198 15036 23204 15048
rect 23256 15036 23262 15088
rect 24397 15011 24455 15017
rect 24397 14977 24409 15011
rect 24443 15008 24455 15011
rect 24780 15008 24808 15104
rect 24443 14980 24808 15008
rect 24443 14977 24455 14980
rect 24397 14971 24455 14977
rect 22465 14943 22523 14949
rect 22465 14909 22477 14943
rect 22511 14909 22523 14943
rect 22465 14903 22523 14909
rect 25317 14943 25375 14949
rect 25317 14909 25329 14943
rect 25363 14940 25375 14943
rect 25682 14940 25688 14952
rect 25363 14912 25688 14940
rect 25363 14909 25375 14912
rect 25317 14903 25375 14909
rect 25682 14900 25688 14912
rect 25740 14940 25746 14952
rect 25869 14943 25927 14949
rect 25869 14940 25881 14943
rect 25740 14912 25881 14940
rect 25740 14900 25746 14912
rect 25869 14909 25881 14912
rect 25915 14909 25927 14943
rect 25869 14903 25927 14909
rect 22738 14872 22744 14884
rect 22296 14844 22744 14872
rect 22738 14832 22744 14844
rect 22796 14832 22802 14884
rect 24210 14872 24216 14884
rect 24123 14844 24216 14872
rect 24210 14832 24216 14844
rect 24268 14872 24274 14884
rect 25133 14875 25191 14881
rect 25133 14872 25145 14875
rect 24268 14844 25145 14872
rect 24268 14832 24274 14844
rect 25133 14841 25145 14844
rect 25179 14841 25191 14875
rect 25133 14835 25191 14841
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 17000 14776 17417 14804
rect 17000 14764 17006 14776
rect 17405 14773 17417 14776
rect 17451 14773 17463 14807
rect 19426 14804 19432 14816
rect 19387 14776 19432 14804
rect 17405 14767 17463 14773
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 20809 14807 20867 14813
rect 20809 14773 20821 14807
rect 20855 14804 20867 14807
rect 20990 14804 20996 14816
rect 20855 14776 20996 14804
rect 20855 14773 20867 14776
rect 20809 14767 20867 14773
rect 20990 14764 20996 14776
rect 21048 14804 21054 14816
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 21048 14776 21373 14804
rect 21048 14764 21054 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 23477 14807 23535 14813
rect 23477 14773 23489 14807
rect 23523 14804 23535 14807
rect 24121 14807 24179 14813
rect 24121 14804 24133 14807
rect 23523 14776 24133 14804
rect 23523 14773 23535 14776
rect 23477 14767 23535 14773
rect 24121 14773 24133 14776
rect 24167 14804 24179 14807
rect 24762 14804 24768 14816
rect 24167 14776 24768 14804
rect 24167 14773 24179 14776
rect 24121 14767 24179 14773
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 4525 14603 4583 14609
rect 4525 14600 4537 14603
rect 3927 14572 4537 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 4525 14569 4537 14572
rect 4571 14600 4583 14603
rect 5166 14600 5172 14612
rect 4571 14572 5172 14600
rect 4571 14569 4583 14572
rect 4525 14563 4583 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5261 14603 5319 14609
rect 5261 14569 5273 14603
rect 5307 14600 5319 14603
rect 5442 14600 5448 14612
rect 5307 14572 5448 14600
rect 5307 14569 5319 14572
rect 5261 14563 5319 14569
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 5629 14603 5687 14609
rect 5629 14569 5641 14603
rect 5675 14600 5687 14603
rect 6086 14600 6092 14612
rect 5675 14572 6092 14600
rect 5675 14569 5687 14572
rect 5629 14563 5687 14569
rect 4614 14532 4620 14544
rect 4575 14504 4620 14532
rect 4614 14492 4620 14504
rect 4672 14492 4678 14544
rect 6012 14541 6040 14572
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7156 14572 8217 14600
rect 7156 14560 7162 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8754 14600 8760 14612
rect 8715 14572 8760 14600
rect 8205 14563 8263 14569
rect 8754 14560 8760 14572
rect 8812 14600 8818 14612
rect 9033 14603 9091 14609
rect 9033 14600 9045 14603
rect 8812 14572 9045 14600
rect 8812 14560 8818 14572
rect 9033 14569 9045 14572
rect 9079 14600 9091 14603
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9079 14572 9413 14600
rect 9079 14569 9091 14572
rect 9033 14563 9091 14569
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 10965 14603 11023 14609
rect 10965 14569 10977 14603
rect 11011 14600 11023 14603
rect 11054 14600 11060 14612
rect 11011 14572 11060 14600
rect 11011 14569 11023 14572
rect 10965 14563 11023 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12308 14572 12725 14600
rect 12308 14560 12314 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 13081 14603 13139 14609
rect 13081 14569 13093 14603
rect 13127 14600 13139 14603
rect 13170 14600 13176 14612
rect 13127 14572 13176 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 18966 14600 18972 14612
rect 18923 14572 18972 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 21910 14560 21916 14612
rect 21968 14600 21974 14612
rect 22094 14600 22100 14612
rect 21968 14572 22100 14600
rect 21968 14560 21974 14572
rect 22094 14560 22100 14572
rect 22152 14600 22158 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 22152 14572 22293 14600
rect 22152 14560 22158 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 22646 14560 22652 14612
rect 22704 14600 22710 14612
rect 22833 14603 22891 14609
rect 22833 14600 22845 14603
rect 22704 14572 22845 14600
rect 22704 14560 22710 14572
rect 22833 14569 22845 14572
rect 22879 14569 22891 14603
rect 22833 14563 22891 14569
rect 23014 14560 23020 14612
rect 23072 14560 23078 14612
rect 23385 14603 23443 14609
rect 23385 14569 23397 14603
rect 23431 14600 23443 14603
rect 24210 14600 24216 14612
rect 23431 14572 24216 14600
rect 23431 14569 23443 14572
rect 23385 14563 23443 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 5988 14535 6046 14541
rect 5988 14501 6000 14535
rect 6034 14501 6046 14535
rect 5988 14495 6046 14501
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 7653 14535 7711 14541
rect 7653 14532 7665 14535
rect 7616 14504 7665 14532
rect 7616 14492 7622 14504
rect 7653 14501 7665 14504
rect 7699 14501 7711 14535
rect 10134 14532 10140 14544
rect 10095 14504 10140 14532
rect 7653 14495 7711 14501
rect 10134 14492 10140 14504
rect 10192 14492 10198 14544
rect 11609 14535 11667 14541
rect 11609 14501 11621 14535
rect 11655 14532 11667 14535
rect 12342 14532 12348 14544
rect 11655 14504 12348 14532
rect 11655 14501 11667 14504
rect 11609 14495 11667 14501
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 12618 14492 12624 14544
rect 12676 14532 12682 14544
rect 13262 14532 13268 14544
rect 12676 14504 13268 14532
rect 12676 14492 12682 14504
rect 13262 14492 13268 14504
rect 13320 14492 13326 14544
rect 14090 14532 14096 14544
rect 14051 14504 14096 14532
rect 14090 14492 14096 14504
rect 14148 14492 14154 14544
rect 19613 14535 19671 14541
rect 19260 14504 19472 14532
rect 1762 14473 1768 14476
rect 1756 14464 1768 14473
rect 1723 14436 1768 14464
rect 1756 14427 1768 14436
rect 1762 14424 1768 14427
rect 1820 14424 1826 14476
rect 8021 14467 8079 14473
rect 8021 14464 8033 14467
rect 5736 14436 8033 14464
rect 1486 14396 1492 14408
rect 1447 14368 1492 14396
rect 1486 14356 1492 14368
rect 1544 14356 1550 14408
rect 4706 14396 4712 14408
rect 4667 14368 4712 14396
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 5442 14356 5448 14408
rect 5500 14396 5506 14408
rect 5736 14405 5764 14436
rect 8021 14433 8033 14436
rect 8067 14464 8079 14467
rect 8202 14464 8208 14476
rect 8067 14436 8208 14464
rect 8067 14433 8079 14436
rect 8021 14427 8079 14433
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 10091 14436 11529 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 11517 14433 11529 14436
rect 11563 14464 11575 14467
rect 12434 14464 12440 14476
rect 11563 14436 12440 14464
rect 11563 14433 11575 14436
rect 11517 14427 11575 14433
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 13354 14464 13360 14476
rect 13219 14436 13360 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 13354 14424 13360 14436
rect 13412 14464 13418 14476
rect 14461 14467 14519 14473
rect 14461 14464 14473 14467
rect 13412 14436 14473 14464
rect 13412 14424 13418 14436
rect 14461 14433 14473 14436
rect 14507 14433 14519 14467
rect 14461 14427 14519 14433
rect 15556 14467 15614 14473
rect 15556 14433 15568 14467
rect 15602 14464 15614 14467
rect 15838 14464 15844 14476
rect 15602 14436 15844 14464
rect 15602 14433 15614 14436
rect 15556 14427 15614 14433
rect 15838 14424 15844 14436
rect 15896 14424 15902 14476
rect 17681 14467 17739 14473
rect 17681 14433 17693 14467
rect 17727 14464 17739 14467
rect 18138 14464 18144 14476
rect 17727 14436 18144 14464
rect 17727 14433 17739 14436
rect 17681 14427 17739 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5500 14368 5733 14396
rect 5500 14356 5506 14368
rect 5721 14365 5733 14368
rect 5767 14365 5779 14399
rect 11790 14396 11796 14408
rect 11751 14368 11796 14396
rect 5721 14359 5779 14365
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13136 14368 13277 14396
rect 13136 14356 13142 14368
rect 13265 14365 13277 14368
rect 13311 14396 13323 14399
rect 13814 14396 13820 14408
rect 13311 14368 13820 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 18230 14396 18236 14408
rect 18191 14368 18236 14396
rect 18230 14356 18236 14368
rect 18288 14356 18294 14408
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 19260 14396 19288 14504
rect 19337 14467 19395 14473
rect 19337 14433 19349 14467
rect 19383 14433 19395 14467
rect 19444 14464 19472 14504
rect 19613 14501 19625 14535
rect 19659 14532 19671 14535
rect 20162 14532 20168 14544
rect 19659 14504 20168 14532
rect 19659 14501 19671 14504
rect 19613 14495 19671 14501
rect 20162 14492 20168 14504
rect 20220 14492 20226 14544
rect 20717 14535 20775 14541
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 21358 14532 21364 14544
rect 20763 14504 21364 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 21358 14492 21364 14504
rect 21416 14492 21422 14544
rect 23032 14532 23060 14560
rect 22480 14504 23060 14532
rect 20254 14464 20260 14476
rect 19444 14436 20260 14464
rect 19337 14427 19395 14433
rect 18472 14368 19288 14396
rect 18472 14356 18478 14368
rect 19352 14340 19380 14427
rect 20254 14424 20260 14436
rect 20312 14464 20318 14476
rect 21168 14467 21226 14473
rect 21168 14464 21180 14467
rect 20312 14436 21180 14464
rect 20312 14424 20318 14436
rect 21168 14433 21180 14436
rect 21214 14464 21226 14467
rect 22278 14464 22284 14476
rect 21214 14436 22284 14464
rect 21214 14433 21226 14436
rect 21168 14427 21226 14433
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 20714 14356 20720 14408
rect 20772 14396 20778 14408
rect 20901 14399 20959 14405
rect 20901 14396 20913 14399
rect 20772 14368 20913 14396
rect 20772 14356 20778 14368
rect 20901 14365 20913 14368
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22480 14396 22508 14504
rect 23842 14492 23848 14544
rect 23900 14532 23906 14544
rect 24397 14535 24455 14541
rect 24397 14532 24409 14535
rect 23900 14504 24409 14532
rect 23900 14492 23906 14504
rect 24397 14501 24409 14504
rect 24443 14501 24455 14535
rect 24397 14495 24455 14501
rect 23566 14424 23572 14476
rect 23624 14464 23630 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23624 14436 23765 14464
rect 23624 14424 23630 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 23753 14427 23811 14433
rect 24949 14467 25007 14473
rect 24949 14433 24961 14467
rect 24995 14464 25007 14467
rect 25038 14464 25044 14476
rect 24995 14436 25044 14464
rect 24995 14433 25007 14436
rect 24949 14427 25007 14433
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 22152 14368 22508 14396
rect 22152 14356 22158 14368
rect 23474 14356 23480 14408
rect 23532 14396 23538 14408
rect 23845 14399 23903 14405
rect 23845 14396 23857 14399
rect 23532 14368 23857 14396
rect 23532 14356 23538 14368
rect 23845 14365 23857 14368
rect 23891 14365 23903 14399
rect 24026 14396 24032 14408
rect 23987 14368 24032 14396
rect 23845 14359 23903 14365
rect 24026 14356 24032 14368
rect 24084 14356 24090 14408
rect 25222 14396 25228 14408
rect 25183 14368 25228 14396
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 3513 14331 3571 14337
rect 3513 14297 3525 14331
rect 3559 14328 3571 14331
rect 17034 14328 17040 14340
rect 3559 14300 4200 14328
rect 3559 14297 3571 14300
rect 3513 14291 3571 14297
rect 4172 14272 4200 14300
rect 16224 14300 17040 14328
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 2869 14263 2927 14269
rect 2869 14260 2881 14263
rect 2832 14232 2881 14260
rect 2832 14220 2838 14232
rect 2869 14229 2881 14232
rect 2915 14229 2927 14263
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 2869 14223 2927 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 7098 14260 7104 14272
rect 7059 14232 7104 14260
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 11149 14263 11207 14269
rect 11149 14229 11161 14263
rect 11195 14260 11207 14263
rect 11330 14260 11336 14272
rect 11195 14232 11336 14260
rect 11195 14229 11207 14232
rect 11149 14223 11207 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12802 14260 12808 14272
rect 12575 14232 12808 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12802 14220 12808 14232
rect 12860 14260 12866 14272
rect 13170 14260 13176 14272
rect 12860 14232 13176 14260
rect 12860 14220 12866 14232
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13262 14220 13268 14272
rect 13320 14260 13326 14272
rect 13722 14260 13728 14272
rect 13320 14232 13728 14260
rect 13320 14220 13326 14232
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 13817 14263 13875 14269
rect 13817 14229 13829 14263
rect 13863 14260 13875 14263
rect 13906 14260 13912 14272
rect 13863 14232 13912 14260
rect 13863 14229 13875 14232
rect 13817 14223 13875 14229
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 14921 14263 14979 14269
rect 14921 14229 14933 14263
rect 14967 14260 14979 14263
rect 15470 14260 15476 14272
rect 14967 14232 15476 14260
rect 14967 14229 14979 14232
rect 14921 14223 14979 14229
rect 15470 14220 15476 14232
rect 15528 14260 15534 14272
rect 16224 14260 16252 14300
rect 17034 14288 17040 14300
rect 17092 14328 17098 14340
rect 17221 14331 17279 14337
rect 17221 14328 17233 14331
rect 17092 14300 17233 14328
rect 17092 14288 17098 14300
rect 17221 14297 17233 14300
rect 17267 14297 17279 14331
rect 17221 14291 17279 14297
rect 17773 14331 17831 14337
rect 17773 14297 17785 14331
rect 17819 14328 17831 14331
rect 19334 14328 19340 14340
rect 17819 14300 19340 14328
rect 17819 14297 17831 14300
rect 17773 14291 17831 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 23492 14328 23520 14356
rect 23256 14300 23520 14328
rect 23256 14288 23262 14300
rect 15528 14232 16252 14260
rect 15528 14220 15534 14232
rect 16298 14220 16304 14272
rect 16356 14260 16362 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16356 14232 16681 14260
rect 16356 14220 16362 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 18782 14220 18788 14272
rect 18840 14260 18846 14272
rect 19153 14263 19211 14269
rect 19153 14260 19165 14263
rect 18840 14232 19165 14260
rect 18840 14220 18846 14232
rect 19153 14229 19165 14232
rect 19199 14260 19211 14263
rect 19242 14260 19248 14272
rect 19199 14232 19248 14260
rect 19199 14229 19211 14232
rect 19153 14223 19211 14229
rect 19242 14220 19248 14232
rect 19300 14260 19306 14272
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19300 14232 20085 14260
rect 19300 14220 19306 14232
rect 20073 14229 20085 14232
rect 20119 14229 20131 14263
rect 23290 14260 23296 14272
rect 23251 14232 23296 14260
rect 20073 14223 20131 14229
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 26326 14220 26332 14272
rect 26384 14260 26390 14272
rect 27062 14260 27068 14272
rect 26384 14232 27068 14260
rect 26384 14220 26390 14232
rect 27062 14220 27068 14232
rect 27120 14220 27126 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2225 14059 2283 14065
rect 2225 14025 2237 14059
rect 2271 14056 2283 14059
rect 2314 14056 2320 14068
rect 2271 14028 2320 14056
rect 2271 14025 2283 14028
rect 2225 14019 2283 14025
rect 2314 14016 2320 14028
rect 2372 14016 2378 14068
rect 2409 14059 2467 14065
rect 2409 14025 2421 14059
rect 2455 14056 2467 14059
rect 3050 14056 3056 14068
rect 2455 14028 3056 14056
rect 2455 14025 2467 14028
rect 2409 14019 2467 14025
rect 3050 14016 3056 14028
rect 3108 14056 3114 14068
rect 3786 14056 3792 14068
rect 3108 14028 3792 14056
rect 3108 14016 3114 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 4706 14056 4712 14068
rect 4667 14028 4712 14056
rect 4706 14016 4712 14028
rect 4764 14056 4770 14068
rect 5994 14056 6000 14068
rect 4764 14028 6000 14056
rect 4764 14016 4770 14028
rect 5994 14016 6000 14028
rect 6052 14056 6058 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6052 14028 6561 14056
rect 6052 14016 6058 14028
rect 6549 14025 6561 14028
rect 6595 14056 6607 14059
rect 7098 14056 7104 14068
rect 6595 14028 7104 14056
rect 6595 14025 6607 14028
rect 6549 14019 6607 14025
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 8202 14056 8208 14068
rect 8163 14028 8208 14056
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 10042 14016 10048 14068
rect 10100 14056 10106 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 10100 14028 10241 14056
rect 10100 14016 10106 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12492 14028 12537 14056
rect 12492 14016 12498 14028
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13446 14056 13452 14068
rect 13044 14028 13452 14056
rect 13044 14016 13050 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14550 14056 14556 14068
rect 14332 14028 14556 14056
rect 14332 14016 14338 14028
rect 14550 14016 14556 14028
rect 14608 14056 14614 14068
rect 14645 14059 14703 14065
rect 14645 14056 14657 14059
rect 14608 14028 14657 14056
rect 14608 14016 14614 14028
rect 14645 14025 14657 14028
rect 14691 14056 14703 14059
rect 15838 14056 15844 14068
rect 14691 14028 14964 14056
rect 15799 14028 15844 14056
rect 14691 14025 14703 14028
rect 14645 14019 14703 14025
rect 2590 13988 2596 14000
rect 2551 13960 2596 13988
rect 2590 13948 2596 13960
rect 2648 13948 2654 14000
rect 3970 13948 3976 14000
rect 4028 13988 4034 14000
rect 5169 13991 5227 13997
rect 5169 13988 5181 13991
rect 4028 13960 5181 13988
rect 4028 13948 4034 13960
rect 5169 13957 5181 13960
rect 5215 13957 5227 13991
rect 5169 13951 5227 13957
rect 6089 13991 6147 13997
rect 6089 13957 6101 13991
rect 6135 13988 6147 13991
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 6135 13960 6837 13988
rect 6135 13957 6147 13960
rect 6089 13951 6147 13957
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 6825 13951 6883 13957
rect 7300 13960 7849 13988
rect 5077 13923 5135 13929
rect 1412 13892 2820 13920
rect 1412 13861 1440 13892
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13821 1455 13855
rect 1397 13815 1455 13821
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2590 13852 2596 13864
rect 1719 13824 2596 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13821 2743 13855
rect 2685 13815 2743 13821
rect 1486 13744 1492 13796
rect 1544 13784 1550 13796
rect 1946 13784 1952 13796
rect 1544 13756 1952 13784
rect 1544 13744 1550 13756
rect 1946 13744 1952 13756
rect 2004 13784 2010 13796
rect 2409 13787 2467 13793
rect 2409 13784 2421 13787
rect 2004 13756 2421 13784
rect 2004 13744 2010 13756
rect 2409 13753 2421 13756
rect 2455 13784 2467 13787
rect 2700 13784 2728 13815
rect 2455 13756 2728 13784
rect 2792 13784 2820 13892
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5721 13923 5779 13929
rect 5721 13920 5733 13923
rect 5123 13892 5733 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5721 13889 5733 13892
rect 5767 13920 5779 13923
rect 6730 13920 6736 13932
rect 5767 13892 6736 13920
rect 5767 13889 5779 13892
rect 5721 13883 5779 13889
rect 6730 13880 6736 13892
rect 6788 13880 6794 13932
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7300 13929 7328 13960
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 7837 13951 7895 13957
rect 12253 13991 12311 13997
rect 12253 13957 12265 13991
rect 12299 13988 12311 13991
rect 12894 13988 12900 14000
rect 12299 13960 12900 13988
rect 12299 13957 12311 13960
rect 12253 13951 12311 13957
rect 12894 13948 12900 13960
rect 12952 13948 12958 14000
rect 14829 13991 14887 13997
rect 14829 13957 14841 13991
rect 14875 13957 14887 13991
rect 14829 13951 14887 13957
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 7064 13892 7297 13920
rect 7064 13880 7070 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7377 13923 7435 13929
rect 7377 13889 7389 13923
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 11885 13923 11943 13929
rect 8803 13892 8984 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 2958 13861 2964 13864
rect 2952 13852 2964 13861
rect 2919 13824 2964 13852
rect 2952 13815 2964 13824
rect 2958 13812 2964 13815
rect 3016 13812 3022 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 5537 13855 5595 13861
rect 5537 13852 5549 13855
rect 4212 13824 5549 13852
rect 4212 13812 4218 13824
rect 5537 13821 5549 13824
rect 5583 13821 5595 13855
rect 5537 13815 5595 13821
rect 5629 13855 5687 13861
rect 5629 13821 5641 13855
rect 5675 13852 5687 13855
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 5675 13824 6009 13852
rect 5675 13821 5687 13824
rect 5629 13815 5687 13821
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 3234 13784 3240 13796
rect 2792 13756 3240 13784
rect 2455 13753 2467 13756
rect 2409 13747 2467 13753
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 3050 13676 3056 13728
rect 3108 13716 3114 13728
rect 4065 13719 4123 13725
rect 4065 13716 4077 13719
rect 3108 13688 4077 13716
rect 3108 13676 3114 13688
rect 4065 13685 4077 13688
rect 4111 13685 4123 13719
rect 4065 13679 4123 13685
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 5644 13716 5672 13815
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 6144 13824 6193 13852
rect 6144 13812 6150 13824
rect 6181 13821 6193 13824
rect 6227 13821 6239 13855
rect 6181 13815 6239 13821
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7392 13852 7420 13883
rect 7156 13824 7420 13852
rect 8849 13855 8907 13861
rect 7156 13812 7162 13824
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8956 13852 8984 13892
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 11931 13892 13093 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13538 13920 13544 13932
rect 13127 13892 13544 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13538 13880 13544 13892
rect 13596 13880 13602 13932
rect 9105 13855 9163 13861
rect 9105 13852 9117 13855
rect 8956 13824 9117 13852
rect 8849 13815 8907 13821
rect 9105 13821 9117 13824
rect 9151 13852 9163 13855
rect 9582 13852 9588 13864
rect 9151 13824 9588 13852
rect 9151 13821 9163 13824
rect 9105 13815 9163 13821
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 6972 13756 7205 13784
rect 6972 13744 6978 13756
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 8864 13784 8892 13815
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13852 10931 13855
rect 12342 13852 12348 13864
rect 10919 13824 12348 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13832 13824 14197 13852
rect 8812 13756 8892 13784
rect 11333 13787 11391 13793
rect 8812 13744 8818 13756
rect 11333 13753 11345 13787
rect 11379 13784 11391 13787
rect 12066 13784 12072 13796
rect 11379 13756 12072 13784
rect 11379 13753 11391 13756
rect 11333 13747 11391 13753
rect 12066 13744 12072 13756
rect 12124 13744 12130 13796
rect 13078 13744 13084 13796
rect 13136 13784 13142 13796
rect 13832 13784 13860 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14844 13852 14872 13951
rect 14936 13920 14964 14028
rect 15838 14016 15844 14028
rect 15896 14016 15902 14068
rect 16393 14059 16451 14065
rect 16393 14025 16405 14059
rect 16439 14056 16451 14059
rect 18230 14056 18236 14068
rect 16439 14028 18236 14056
rect 16439 14025 16451 14028
rect 16393 14019 16451 14025
rect 18230 14016 18236 14028
rect 18288 14016 18294 14068
rect 20165 14059 20223 14065
rect 20165 14025 20177 14059
rect 20211 14056 20223 14059
rect 20254 14056 20260 14068
rect 20211 14028 20260 14056
rect 20211 14025 20223 14028
rect 20165 14019 20223 14025
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 20806 14056 20812 14068
rect 20767 14028 20812 14056
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21269 14059 21327 14065
rect 21269 14025 21281 14059
rect 21315 14056 21327 14059
rect 21358 14056 21364 14068
rect 21315 14028 21364 14056
rect 21315 14025 21327 14028
rect 21269 14019 21327 14025
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 22278 14056 22284 14068
rect 22239 14028 22284 14056
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 15856 13988 15884 14016
rect 16022 13988 16028 14000
rect 15856 13960 16028 13988
rect 16022 13948 16028 13960
rect 16080 13988 16086 14000
rect 16482 13988 16488 14000
rect 16080 13960 16488 13988
rect 16080 13948 16086 13960
rect 16482 13948 16488 13960
rect 16540 13948 16546 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 16868 13960 17417 13988
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 14936 13892 15301 13920
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15470 13920 15476 13932
rect 15431 13892 15476 13920
rect 15289 13883 15347 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 16666 13880 16672 13932
rect 16724 13920 16730 13932
rect 16868 13929 16896 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 17865 13991 17923 13997
rect 17865 13957 17877 13991
rect 17911 13988 17923 13991
rect 18414 13988 18420 14000
rect 17911 13960 18420 13988
rect 17911 13957 17923 13960
rect 17865 13951 17923 13957
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 16853 13923 16911 13929
rect 16853 13920 16865 13923
rect 16724 13892 16865 13920
rect 16724 13880 16730 13892
rect 16853 13889 16865 13892
rect 16899 13889 16911 13923
rect 16853 13883 16911 13889
rect 16945 13923 17003 13929
rect 16945 13889 16957 13923
rect 16991 13920 17003 13923
rect 18601 13923 18659 13929
rect 18601 13920 18613 13923
rect 16991 13892 18613 13920
rect 16991 13889 17003 13892
rect 16945 13883 17003 13889
rect 18601 13889 18613 13892
rect 18647 13920 18659 13923
rect 20824 13920 20852 14016
rect 22649 13991 22707 13997
rect 22649 13957 22661 13991
rect 22695 13988 22707 13991
rect 22922 13988 22928 14000
rect 22695 13960 22928 13988
rect 22695 13957 22707 13960
rect 22649 13951 22707 13957
rect 22922 13948 22928 13960
rect 22980 13948 22986 14000
rect 23658 13948 23664 14000
rect 23716 13988 23722 14000
rect 24578 13988 24584 14000
rect 23716 13960 24584 13988
rect 23716 13948 23722 13960
rect 24578 13948 24584 13960
rect 24636 13948 24642 14000
rect 21729 13923 21787 13929
rect 21729 13920 21741 13923
rect 18647 13892 18920 13920
rect 20824 13892 21741 13920
rect 18647 13889 18659 13892
rect 18601 13883 18659 13889
rect 16301 13855 16359 13861
rect 14844 13824 15148 13852
rect 14185 13815 14243 13821
rect 13136 13756 13860 13784
rect 15120 13784 15148 13824
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16960 13852 16988 13883
rect 16347 13824 16988 13852
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18782 13852 18788 13864
rect 18012 13824 18788 13852
rect 18012 13812 18018 13824
rect 18782 13812 18788 13824
rect 18840 13812 18846 13864
rect 18892 13852 18920 13892
rect 21729 13889 21741 13892
rect 21775 13889 21787 13923
rect 21910 13920 21916 13932
rect 21871 13892 21916 13920
rect 21729 13883 21787 13889
rect 19058 13861 19064 13864
rect 19041 13855 19064 13861
rect 19041 13852 19053 13855
rect 18892 13824 19053 13852
rect 19041 13821 19053 13824
rect 19116 13852 19122 13864
rect 21744 13852 21772 13883
rect 21910 13880 21916 13892
rect 21968 13880 21974 13932
rect 22738 13880 22744 13932
rect 22796 13920 22802 13932
rect 23014 13920 23020 13932
rect 22796 13892 23020 13920
rect 22796 13880 22802 13892
rect 23014 13880 23020 13892
rect 23072 13880 23078 13932
rect 23474 13880 23480 13932
rect 23532 13920 23538 13932
rect 24213 13923 24271 13929
rect 24213 13920 24225 13923
rect 23532 13892 24225 13920
rect 23532 13880 23538 13892
rect 24213 13889 24225 13892
rect 24259 13920 24271 13923
rect 24673 13923 24731 13929
rect 24673 13920 24685 13923
rect 24259 13892 24685 13920
rect 24259 13889 24271 13892
rect 24213 13883 24271 13889
rect 24673 13889 24685 13892
rect 24719 13889 24731 13923
rect 25038 13920 25044 13932
rect 24999 13892 25044 13920
rect 24673 13883 24731 13889
rect 25038 13880 25044 13892
rect 25096 13880 25102 13932
rect 25406 13920 25412 13932
rect 25367 13892 25412 13920
rect 25406 13880 25412 13892
rect 25464 13880 25470 13932
rect 21818 13852 21824 13864
rect 19116 13824 19189 13852
rect 21744 13824 21824 13852
rect 19041 13815 19064 13821
rect 19058 13812 19064 13815
rect 19116 13812 19122 13824
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13852 23167 13855
rect 23566 13852 23572 13864
rect 23155 13824 23572 13852
rect 23155 13821 23167 13824
rect 23109 13815 23167 13821
rect 23566 13812 23572 13824
rect 23624 13852 23630 13864
rect 23750 13852 23756 13864
rect 23624 13824 23756 13852
rect 23624 13812 23630 13824
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 23842 13812 23848 13864
rect 23900 13852 23906 13864
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 23900 13824 24133 13852
rect 23900 13812 23906 13824
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 24121 13815 24179 13821
rect 24946 13812 24952 13864
rect 25004 13852 25010 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 25004 13824 25237 13852
rect 25004 13812 25010 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 25961 13855 26019 13861
rect 25961 13852 25973 13855
rect 25271 13824 25973 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25961 13821 25973 13824
rect 26007 13821 26019 13855
rect 25961 13815 26019 13821
rect 16761 13787 16819 13793
rect 16761 13784 16773 13787
rect 15120 13756 16773 13784
rect 13136 13744 13142 13756
rect 16761 13753 16773 13756
rect 16807 13784 16819 13787
rect 17218 13784 17224 13796
rect 16807 13756 17224 13784
rect 16807 13753 16819 13756
rect 16761 13747 16819 13753
rect 17218 13744 17224 13756
rect 17276 13744 17282 13796
rect 23385 13787 23443 13793
rect 23385 13753 23397 13787
rect 23431 13784 23443 13787
rect 24029 13787 24087 13793
rect 24029 13784 24041 13787
rect 23431 13756 24041 13784
rect 23431 13753 23443 13756
rect 23385 13747 23443 13753
rect 24029 13753 24041 13756
rect 24075 13784 24087 13787
rect 24670 13784 24676 13796
rect 24075 13756 24676 13784
rect 24075 13753 24087 13756
rect 24029 13747 24087 13753
rect 24670 13744 24676 13756
rect 24728 13744 24734 13796
rect 5592 13688 5672 13716
rect 11241 13719 11299 13725
rect 5592 13676 5598 13688
rect 11241 13685 11253 13719
rect 11287 13716 11299 13719
rect 11790 13716 11796 13728
rect 11287 13688 11796 13716
rect 11287 13685 11299 13688
rect 11241 13679 11299 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12526 13676 12532 13728
rect 12584 13716 12590 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12584 13688 12817 13716
rect 12584 13676 12590 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 13538 13716 13544 13728
rect 13499 13688 13544 13716
rect 12805 13679 12863 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 14734 13676 14740 13728
rect 14792 13716 14798 13728
rect 15197 13719 15255 13725
rect 15197 13716 15209 13719
rect 14792 13688 15209 13716
rect 14792 13676 14798 13688
rect 15197 13685 15209 13688
rect 15243 13685 15255 13719
rect 15197 13679 15255 13685
rect 21177 13719 21235 13725
rect 21177 13685 21189 13719
rect 21223 13716 21235 13719
rect 21634 13716 21640 13728
rect 21223 13688 21640 13716
rect 21223 13685 21235 13688
rect 21177 13679 21235 13685
rect 21634 13676 21640 13688
rect 21692 13676 21698 13728
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 23661 13719 23719 13725
rect 23661 13716 23673 13719
rect 23532 13688 23673 13716
rect 23532 13676 23538 13688
rect 23661 13685 23673 13688
rect 23707 13685 23719 13719
rect 23661 13679 23719 13685
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2041 13515 2099 13521
rect 2041 13512 2053 13515
rect 1912 13484 2053 13512
rect 1912 13472 1918 13484
rect 2041 13481 2053 13484
rect 2087 13481 2099 13515
rect 2041 13475 2099 13481
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 3234 13512 3240 13524
rect 3191 13484 3240 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3234 13472 3240 13484
rect 3292 13512 3298 13524
rect 3970 13512 3976 13524
rect 3292 13484 3976 13512
rect 3292 13472 3298 13484
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 4120 13484 4261 13512
rect 4120 13472 4126 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 4614 13512 4620 13524
rect 4575 13484 4620 13512
rect 4249 13475 4307 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 6972 13484 7481 13512
rect 6972 13472 6978 13484
rect 7469 13481 7481 13484
rect 7515 13481 7527 13515
rect 7469 13475 7527 13481
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7708 13484 8033 13512
rect 7708 13472 7714 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8386 13512 8392 13524
rect 8347 13484 8392 13512
rect 8021 13475 8079 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8570 13512 8576 13524
rect 8527 13484 8576 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8812 13484 9045 13512
rect 8812 13472 8818 13484
rect 9033 13481 9045 13484
rect 9079 13512 9091 13515
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9079 13484 9413 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 9766 13512 9772 13524
rect 9727 13484 9772 13512
rect 9401 13475 9459 13481
rect 2590 13404 2596 13456
rect 2648 13444 2654 13456
rect 5804 13447 5862 13453
rect 2648 13416 4108 13444
rect 2648 13404 2654 13416
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2409 13379 2467 13385
rect 2409 13376 2421 13379
rect 2280 13348 2421 13376
rect 2280 13336 2286 13348
rect 2409 13345 2421 13348
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2682 13376 2688 13388
rect 2547 13348 2688 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 4080 13385 4108 13416
rect 5804 13413 5816 13447
rect 5850 13444 5862 13447
rect 5994 13444 6000 13456
rect 5850 13416 6000 13444
rect 5850 13413 5862 13416
rect 5804 13407 5862 13413
rect 5994 13404 6000 13416
rect 6052 13404 6058 13456
rect 7929 13447 7987 13453
rect 7929 13413 7941 13447
rect 7975 13444 7987 13447
rect 8662 13444 8668 13456
rect 7975 13416 8668 13444
rect 7975 13413 7987 13416
rect 7929 13407 7987 13413
rect 8662 13404 8668 13416
rect 8720 13404 8726 13456
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4614 13376 4620 13388
rect 4111 13348 4620 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 9416 13376 9444 13475
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14792 13484 14841 13512
rect 14792 13472 14798 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 14829 13475 14887 13481
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 17218 13512 17224 13524
rect 17179 13484 17224 13512
rect 16669 13475 16727 13481
rect 17218 13472 17224 13484
rect 17276 13472 17282 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19889 13515 19947 13521
rect 19889 13512 19901 13515
rect 19392 13484 19901 13512
rect 19392 13472 19398 13484
rect 19889 13481 19901 13484
rect 19935 13481 19947 13515
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 19889 13475 19947 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 21910 13512 21916 13524
rect 21871 13484 21916 13512
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 22186 13472 22192 13524
rect 22244 13512 22250 13524
rect 22649 13515 22707 13521
rect 22649 13512 22661 13515
rect 22244 13484 22661 13512
rect 22244 13472 22250 13484
rect 22649 13481 22661 13484
rect 22695 13481 22707 13515
rect 22649 13475 22707 13481
rect 23198 13472 23204 13524
rect 23256 13512 23262 13524
rect 23477 13515 23535 13521
rect 23477 13512 23489 13515
rect 23256 13484 23489 13512
rect 23256 13472 23262 13484
rect 23477 13481 23489 13484
rect 23523 13481 23535 13515
rect 23477 13475 23535 13481
rect 24210 13472 24216 13524
rect 24268 13512 24274 13524
rect 25041 13515 25099 13521
rect 25041 13512 25053 13515
rect 24268 13484 25053 13512
rect 24268 13472 24274 13484
rect 25041 13481 25053 13484
rect 25087 13481 25099 13515
rect 25041 13475 25099 13481
rect 15470 13404 15476 13456
rect 15528 13453 15534 13456
rect 15528 13447 15592 13453
rect 15528 13413 15546 13447
rect 15580 13413 15592 13447
rect 15528 13407 15592 13413
rect 15528 13404 15534 13407
rect 17034 13404 17040 13456
rect 17092 13444 17098 13456
rect 17770 13444 17776 13456
rect 17092 13416 17776 13444
rect 17092 13404 17098 13416
rect 17770 13404 17776 13416
rect 17828 13444 17834 13456
rect 18202 13447 18260 13453
rect 18202 13444 18214 13447
rect 17828 13416 18214 13444
rect 17828 13404 17834 13416
rect 18202 13413 18214 13416
rect 18248 13413 18260 13447
rect 18202 13407 18260 13413
rect 21361 13447 21419 13453
rect 21361 13413 21373 13447
rect 21407 13444 21419 13447
rect 22738 13444 22744 13456
rect 21407 13416 22744 13444
rect 21407 13413 21419 13416
rect 21361 13407 21419 13413
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 23106 13404 23112 13456
rect 23164 13444 23170 13456
rect 23906 13447 23964 13453
rect 23906 13444 23918 13447
rect 23164 13416 23918 13444
rect 23164 13404 23170 13416
rect 23906 13413 23918 13416
rect 23952 13413 23964 13447
rect 23906 13407 23964 13413
rect 10134 13376 10140 13388
rect 9416 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13376 10198 13388
rect 10229 13379 10287 13385
rect 10229 13376 10241 13379
rect 10192 13348 10241 13376
rect 10192 13336 10198 13348
rect 10229 13345 10241 13348
rect 10275 13345 10287 13379
rect 10229 13339 10287 13345
rect 10318 13336 10324 13388
rect 10376 13376 10382 13388
rect 10496 13379 10554 13385
rect 10496 13376 10508 13379
rect 10376 13348 10508 13376
rect 10376 13336 10382 13348
rect 10496 13345 10508 13348
rect 10542 13376 10554 13379
rect 11790 13376 11796 13388
rect 10542 13348 11796 13376
rect 10542 13345 10554 13348
rect 10496 13339 10554 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12713 13379 12771 13385
rect 12713 13376 12725 13379
rect 12216 13348 12725 13376
rect 12216 13336 12222 13348
rect 12713 13345 12725 13348
rect 12759 13345 12771 13379
rect 12713 13339 12771 13345
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 15286 13376 15292 13388
rect 14332 13348 15292 13376
rect 14332 13336 14338 13348
rect 15286 13336 15292 13348
rect 15344 13376 15350 13388
rect 16114 13376 16120 13388
rect 15344 13348 16120 13376
rect 15344 13336 15350 13348
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 21266 13376 21272 13388
rect 21227 13348 21272 13376
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 22462 13376 22468 13388
rect 22423 13348 22468 13376
rect 22462 13336 22468 13348
rect 22520 13376 22526 13388
rect 23017 13379 23075 13385
rect 23017 13376 23029 13379
rect 22520 13348 23029 13376
rect 22520 13336 22526 13348
rect 23017 13345 23029 13348
rect 23063 13345 23075 13379
rect 25314 13376 25320 13388
rect 23017 13339 23075 13345
rect 23216 13348 25320 13376
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 3786 13268 3792 13320
rect 3844 13308 3850 13320
rect 5442 13308 5448 13320
rect 3844 13280 5448 13308
rect 3844 13268 3850 13280
rect 5442 13268 5448 13280
rect 5500 13308 5506 13320
rect 5537 13311 5595 13317
rect 5537 13308 5549 13311
rect 5500 13280 5549 13308
rect 5500 13268 5506 13280
rect 5537 13277 5549 13280
rect 5583 13277 5595 13311
rect 5537 13271 5595 13277
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 8573 13311 8631 13317
rect 8573 13308 8585 13311
rect 8536 13280 8585 13308
rect 8536 13268 8542 13280
rect 8573 13277 8585 13280
rect 8619 13277 8631 13311
rect 17954 13308 17960 13320
rect 17915 13280 17960 13308
rect 8573 13271 8631 13277
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 21358 13308 21364 13320
rect 20864 13280 21364 13308
rect 20864 13268 20870 13280
rect 21358 13268 21364 13280
rect 21416 13308 21422 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21416 13280 21465 13308
rect 21416 13268 21422 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 3697 13243 3755 13249
rect 3697 13209 3709 13243
rect 3743 13240 3755 13243
rect 4062 13240 4068 13252
rect 3743 13212 4068 13240
rect 3743 13209 3755 13212
rect 3697 13203 3755 13209
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 6730 13200 6736 13252
rect 6788 13240 6794 13252
rect 6917 13243 6975 13249
rect 6917 13240 6929 13243
rect 6788 13212 6929 13240
rect 6788 13200 6794 13212
rect 6917 13209 6929 13212
rect 6963 13209 6975 13243
rect 6917 13203 6975 13209
rect 12250 13200 12256 13252
rect 12308 13240 12314 13252
rect 14001 13243 14059 13249
rect 14001 13240 14013 13243
rect 12308 13212 14013 13240
rect 12308 13200 12314 13212
rect 14001 13209 14013 13212
rect 14047 13209 14059 13243
rect 14001 13203 14059 13209
rect 1673 13175 1731 13181
rect 1673 13141 1685 13175
rect 1719 13172 1731 13175
rect 1762 13172 1768 13184
rect 1719 13144 1768 13172
rect 1719 13141 1731 13144
rect 1673 13135 1731 13141
rect 1762 13132 1768 13144
rect 1820 13172 1826 13184
rect 3050 13172 3056 13184
rect 1820 13144 3056 13172
rect 1820 13132 1826 13144
rect 3050 13132 3056 13144
rect 3108 13132 3114 13184
rect 5258 13172 5264 13184
rect 5219 13144 5264 13172
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 11606 13172 11612 13184
rect 11567 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 12526 13172 12532 13184
rect 12487 13144 12532 13172
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 14016 13172 14044 13203
rect 19058 13200 19064 13252
rect 19116 13240 19122 13252
rect 19337 13243 19395 13249
rect 19337 13240 19349 13243
rect 19116 13212 19349 13240
rect 19116 13200 19122 13212
rect 19337 13209 19349 13212
rect 19383 13209 19395 13243
rect 19337 13203 19395 13209
rect 20901 13243 20959 13249
rect 20901 13209 20913 13243
rect 20947 13240 20959 13243
rect 23216 13240 23244 13348
rect 25314 13336 25320 13348
rect 25372 13336 25378 13388
rect 23290 13268 23296 13320
rect 23348 13308 23354 13320
rect 23661 13311 23719 13317
rect 23661 13308 23673 13311
rect 23348 13280 23673 13308
rect 23348 13268 23354 13280
rect 23661 13277 23673 13280
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 20947 13212 23244 13240
rect 20947 13209 20959 13212
rect 20901 13203 20959 13209
rect 15930 13172 15936 13184
rect 14016 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 17862 13172 17868 13184
rect 17823 13144 17868 13172
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 23676 13172 23704 13271
rect 23842 13172 23848 13184
rect 23676 13144 23848 13172
rect 23842 13132 23848 13144
rect 23900 13132 23906 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2590 12968 2596 12980
rect 1995 12940 2596 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 3326 12928 3332 12980
rect 3384 12968 3390 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 3384 12940 3433 12968
rect 3384 12928 3390 12940
rect 3421 12937 3433 12940
rect 3467 12937 3479 12971
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3421 12931 3479 12937
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 6052 12940 6193 12968
rect 6052 12928 6058 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6730 12968 6736 12980
rect 6687 12940 6736 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 8536 12940 9137 12968
rect 8536 12928 8542 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10318 12968 10324 12980
rect 10275 12940 10324 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10778 12968 10784 12980
rect 10739 12940 10784 12968
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 12342 12928 12348 12980
rect 12400 12968 12406 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 12400 12940 13277 12968
rect 12400 12928 12406 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 15378 12928 15384 12980
rect 15436 12968 15442 12980
rect 15654 12968 15660 12980
rect 15436 12940 15660 12968
rect 15436 12928 15442 12940
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 17770 12968 17776 12980
rect 17731 12940 17776 12968
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18138 12968 18144 12980
rect 18099 12940 18144 12968
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 20806 12968 20812 12980
rect 20767 12940 20812 12968
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 21266 12968 21272 12980
rect 21227 12940 21272 12968
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22738 12968 22744 12980
rect 22651 12940 22744 12968
rect 22738 12928 22744 12940
rect 22796 12968 22802 12980
rect 23382 12968 23388 12980
rect 22796 12940 23388 12968
rect 22796 12928 22802 12940
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 25590 12968 25596 12980
rect 23492 12940 25596 12968
rect 2406 12860 2412 12912
rect 2464 12900 2470 12912
rect 3145 12903 3203 12909
rect 3145 12900 3157 12903
rect 2464 12872 3157 12900
rect 2464 12860 2470 12872
rect 3145 12869 3157 12872
rect 3191 12900 3203 12903
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 3191 12872 5181 12900
rect 3191 12869 3203 12872
rect 3145 12863 3203 12869
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12832 2743 12835
rect 2774 12832 2780 12844
rect 2731 12804 2780 12832
rect 2731 12801 2743 12804
rect 2685 12795 2743 12801
rect 2774 12792 2780 12804
rect 2832 12832 2838 12844
rect 3050 12832 3056 12844
rect 2832 12804 3056 12832
rect 2832 12792 2838 12804
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3326 12792 3332 12844
rect 3384 12832 3390 12844
rect 3970 12832 3976 12844
rect 3384 12804 3976 12832
rect 3384 12792 3390 12804
rect 3970 12792 3976 12804
rect 4028 12832 4034 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 4028 12804 4077 12832
rect 4028 12792 4034 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4246 12832 4252 12844
rect 4207 12804 4252 12832
rect 4065 12795 4123 12801
rect 2409 12767 2467 12773
rect 2409 12733 2421 12767
rect 2455 12764 2467 12767
rect 2498 12764 2504 12776
rect 2455 12736 2504 12764
rect 2455 12733 2467 12736
rect 2409 12727 2467 12733
rect 2498 12724 2504 12736
rect 2556 12724 2562 12776
rect 4080 12764 4108 12795
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 5258 12832 5264 12844
rect 4672 12804 5264 12832
rect 4672 12792 4678 12804
rect 5258 12792 5264 12804
rect 5316 12832 5322 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5316 12804 5825 12832
rect 5316 12792 5322 12804
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 6748 12832 6776 12928
rect 8386 12860 8392 12912
rect 8444 12900 8450 12912
rect 8757 12903 8815 12909
rect 8757 12900 8769 12903
rect 8444 12872 8769 12900
rect 8444 12860 8450 12872
rect 8757 12869 8769 12872
rect 8803 12869 8815 12903
rect 8757 12863 8815 12869
rect 9861 12903 9919 12909
rect 9861 12869 9873 12903
rect 9907 12900 9919 12903
rect 12894 12900 12900 12912
rect 9907 12872 12900 12900
rect 9907 12869 9919 12872
rect 9861 12863 9919 12869
rect 12894 12860 12900 12872
rect 12952 12860 12958 12912
rect 17788 12900 17816 12928
rect 18966 12900 18972 12912
rect 17788 12872 18972 12900
rect 18966 12860 18972 12872
rect 19024 12900 19030 12912
rect 19153 12903 19211 12909
rect 19153 12900 19165 12903
rect 19024 12872 19165 12900
rect 19024 12860 19030 12872
rect 19153 12869 19165 12872
rect 19199 12900 19211 12903
rect 19426 12900 19432 12912
rect 19199 12872 19432 12900
rect 19199 12869 19211 12872
rect 19153 12863 19211 12869
rect 19426 12860 19432 12872
rect 19484 12860 19490 12912
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 21177 12903 21235 12909
rect 21177 12900 21189 12903
rect 20680 12872 21189 12900
rect 20680 12860 20686 12872
rect 21177 12869 21189 12872
rect 21223 12900 21235 12903
rect 23492 12900 23520 12940
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 21223 12872 23520 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 5859 12804 6132 12832
rect 6748 12804 6960 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 4985 12767 5043 12773
rect 4985 12764 4997 12767
rect 4080 12736 4997 12764
rect 4985 12733 4997 12736
rect 5031 12764 5043 12767
rect 5629 12767 5687 12773
rect 5629 12764 5641 12767
rect 5031 12736 5641 12764
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5629 12733 5641 12736
rect 5675 12733 5687 12767
rect 5629 12727 5687 12733
rect 2222 12696 2228 12708
rect 2056 12668 2228 12696
rect 2056 12637 2084 12668
rect 2222 12656 2228 12668
rect 2280 12696 2286 12708
rect 2866 12696 2872 12708
rect 2280 12668 2872 12696
rect 2280 12656 2286 12668
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 3694 12656 3700 12708
rect 3752 12696 3758 12708
rect 3973 12699 4031 12705
rect 3973 12696 3985 12699
rect 3752 12668 3985 12696
rect 3752 12656 3758 12668
rect 3973 12665 3985 12668
rect 4019 12696 4031 12699
rect 4338 12696 4344 12708
rect 4019 12668 4344 12696
rect 4019 12665 4031 12668
rect 3973 12659 4031 12665
rect 4338 12656 4344 12668
rect 4396 12656 4402 12708
rect 6104 12696 6132 12804
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6932 12764 6960 12804
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 9088 12804 9321 12832
rect 9088 12792 9094 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 11330 12832 11336 12844
rect 11287 12804 11336 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11425 12835 11483 12841
rect 11425 12801 11437 12835
rect 11471 12832 11483 12835
rect 11606 12832 11612 12844
rect 11471 12804 11612 12832
rect 11471 12801 11483 12804
rect 11425 12795 11483 12801
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11790 12832 11796 12844
rect 11751 12804 11796 12832
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13596 12804 13921 12832
rect 13596 12792 13602 12804
rect 13909 12801 13921 12804
rect 13955 12832 13967 12835
rect 13998 12832 14004 12844
rect 13955 12804 14004 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 13998 12792 14004 12804
rect 14056 12792 14062 12844
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12832 18843 12835
rect 19058 12832 19064 12844
rect 18831 12804 19064 12832
rect 18831 12801 18843 12804
rect 18785 12795 18843 12801
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 19444 12832 19472 12860
rect 21744 12841 21772 12872
rect 20257 12835 20315 12841
rect 20257 12832 20269 12835
rect 19444 12804 20269 12832
rect 20257 12801 20269 12804
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 21729 12835 21787 12841
rect 21729 12801 21741 12835
rect 21775 12801 21787 12835
rect 21729 12795 21787 12801
rect 21913 12835 21971 12841
rect 21913 12801 21925 12835
rect 21959 12832 21971 12835
rect 22002 12832 22008 12844
rect 21959 12804 22008 12832
rect 21959 12801 21971 12804
rect 21913 12795 21971 12801
rect 22002 12792 22008 12804
rect 22060 12832 22066 12844
rect 22281 12835 22339 12841
rect 22281 12832 22293 12835
rect 22060 12804 22293 12832
rect 22060 12792 22066 12804
rect 22281 12801 22293 12804
rect 22327 12801 22339 12835
rect 22281 12795 22339 12801
rect 23106 12792 23112 12844
rect 23164 12832 23170 12844
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 23164 12804 23397 12832
rect 23164 12792 23170 12804
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23385 12795 23443 12801
rect 7081 12767 7139 12773
rect 7081 12764 7093 12767
rect 6932 12736 7093 12764
rect 7081 12733 7093 12736
rect 7127 12733 7139 12767
rect 7081 12727 7139 12733
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 9456 12736 10517 12764
rect 9456 12724 9462 12736
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 12250 12764 12256 12776
rect 10551 12736 12256 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12492 12736 12817 12764
rect 12492 12724 12498 12736
rect 12805 12733 12817 12736
rect 12851 12764 12863 12767
rect 13078 12764 13084 12776
rect 12851 12736 13084 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13354 12724 13360 12776
rect 13412 12764 13418 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13412 12736 13645 12764
rect 13412 12724 13418 12736
rect 13633 12733 13645 12736
rect 13679 12733 13691 12767
rect 13633 12727 13691 12733
rect 17862 12724 17868 12776
rect 17920 12764 17926 12776
rect 18414 12764 18420 12776
rect 17920 12736 18420 12764
rect 17920 12724 17926 12736
rect 18414 12724 18420 12736
rect 18472 12764 18478 12776
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18472 12736 18521 12764
rect 18472 12724 18478 12736
rect 18509 12733 18521 12736
rect 18555 12733 18567 12767
rect 18509 12727 18567 12733
rect 19426 12724 19432 12776
rect 19484 12764 19490 12776
rect 20162 12764 20168 12776
rect 19484 12736 20168 12764
rect 19484 12724 19490 12736
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 23842 12764 23848 12776
rect 23803 12736 23848 12764
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 6104 12668 7972 12696
rect 7944 12640 7972 12668
rect 11164 12668 12480 12696
rect 2041 12631 2099 12637
rect 2041 12597 2053 12631
rect 2087 12597 2099 12631
rect 2041 12591 2099 12597
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2501 12631 2559 12637
rect 2501 12628 2513 12631
rect 2464 12600 2513 12628
rect 2464 12588 2470 12600
rect 2501 12597 2513 12600
rect 2547 12597 2559 12631
rect 2501 12591 2559 12597
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 5224 12600 5549 12628
rect 5224 12588 5230 12600
rect 5537 12597 5549 12600
rect 5583 12628 5595 12631
rect 6362 12628 6368 12640
rect 5583 12600 6368 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8205 12631 8263 12637
rect 8205 12628 8217 12631
rect 7984 12600 8217 12628
rect 7984 12588 7990 12600
rect 8205 12597 8217 12600
rect 8251 12597 8263 12631
rect 8205 12591 8263 12597
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 10192 12600 10333 12628
rect 10192 12588 10198 12600
rect 10321 12597 10333 12600
rect 10367 12628 10379 12631
rect 10778 12628 10784 12640
rect 10367 12600 10784 12628
rect 10367 12597 10379 12600
rect 10321 12591 10379 12597
rect 10778 12588 10784 12600
rect 10836 12588 10842 12640
rect 11054 12588 11060 12640
rect 11112 12628 11118 12640
rect 11164 12637 11192 12668
rect 11149 12631 11207 12637
rect 11149 12628 11161 12631
rect 11112 12600 11161 12628
rect 11112 12588 11118 12600
rect 11149 12597 11161 12600
rect 11195 12597 11207 12631
rect 12158 12628 12164 12640
rect 12119 12600 12164 12628
rect 11149 12591 11207 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12452 12637 12480 12668
rect 12986 12656 12992 12708
rect 13044 12696 13050 12708
rect 13725 12699 13783 12705
rect 13725 12696 13737 12699
rect 13044 12668 13737 12696
rect 13044 12656 13050 12668
rect 13725 12665 13737 12668
rect 13771 12665 13783 12699
rect 13725 12659 13783 12665
rect 14366 12656 14372 12708
rect 14424 12696 14430 12708
rect 14522 12699 14580 12705
rect 14522 12696 14534 12699
rect 14424 12668 14534 12696
rect 14424 12656 14430 12668
rect 14522 12665 14534 12668
rect 14568 12665 14580 12699
rect 14522 12659 14580 12665
rect 17497 12699 17555 12705
rect 17497 12665 17509 12699
rect 17543 12696 17555 12699
rect 18601 12699 18659 12705
rect 18601 12696 18613 12699
rect 17543 12668 18613 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 18601 12665 18613 12668
rect 18647 12696 18659 12699
rect 18647 12668 19748 12696
rect 18647 12665 18659 12668
rect 18601 12659 18659 12665
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 12894 12628 12900 12640
rect 12855 12600 12900 12628
rect 12437 12591 12495 12597
rect 12894 12588 12900 12600
rect 12952 12588 12958 12640
rect 15470 12588 15476 12640
rect 15528 12628 15534 12640
rect 15657 12631 15715 12637
rect 15657 12628 15669 12631
rect 15528 12600 15669 12628
rect 15528 12588 15534 12600
rect 15657 12597 15669 12600
rect 15703 12628 15715 12631
rect 16209 12631 16267 12637
rect 16209 12628 16221 12631
rect 15703 12600 16221 12628
rect 15703 12597 15715 12600
rect 15657 12591 15715 12597
rect 16209 12597 16221 12600
rect 16255 12597 16267 12631
rect 16574 12628 16580 12640
rect 16535 12600 16580 12628
rect 16209 12591 16267 12597
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19720 12637 19748 12668
rect 21818 12656 21824 12708
rect 21876 12696 21882 12708
rect 22002 12696 22008 12708
rect 21876 12668 22008 12696
rect 21876 12656 21882 12668
rect 22002 12656 22008 12668
rect 22060 12656 22066 12708
rect 23109 12699 23167 12705
rect 23109 12665 23121 12699
rect 23155 12696 23167 12699
rect 24112 12699 24170 12705
rect 24112 12696 24124 12699
rect 23155 12668 24124 12696
rect 23155 12665 23167 12668
rect 23109 12659 23167 12665
rect 24112 12665 24124 12668
rect 24158 12696 24170 12699
rect 24210 12696 24216 12708
rect 24158 12668 24216 12696
rect 24158 12665 24170 12668
rect 24112 12659 24170 12665
rect 24210 12656 24216 12668
rect 24268 12656 24274 12708
rect 19521 12631 19579 12637
rect 19521 12628 19533 12631
rect 19484 12600 19533 12628
rect 19484 12588 19490 12600
rect 19521 12597 19533 12600
rect 19567 12597 19579 12631
rect 19521 12591 19579 12597
rect 19705 12631 19763 12637
rect 19705 12597 19717 12631
rect 19751 12597 19763 12631
rect 20070 12628 20076 12640
rect 20031 12600 20076 12628
rect 19705 12591 19763 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21637 12631 21695 12637
rect 21637 12628 21649 12631
rect 21416 12600 21649 12628
rect 21416 12588 21422 12600
rect 21637 12597 21649 12600
rect 21683 12597 21695 12631
rect 21637 12591 21695 12597
rect 23566 12588 23572 12640
rect 23624 12628 23630 12640
rect 24762 12628 24768 12640
rect 23624 12600 24768 12628
rect 23624 12588 23630 12600
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 24854 12588 24860 12640
rect 24912 12628 24918 12640
rect 25225 12631 25283 12637
rect 25225 12628 25237 12631
rect 24912 12600 25237 12628
rect 24912 12588 24918 12600
rect 25225 12597 25237 12600
rect 25271 12597 25283 12631
rect 25225 12591 25283 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 2314 12424 2320 12436
rect 1443 12396 2320 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 2409 12427 2467 12433
rect 2409 12393 2421 12427
rect 2455 12424 2467 12427
rect 2682 12424 2688 12436
rect 2455 12396 2688 12424
rect 2455 12393 2467 12396
rect 2409 12387 2467 12393
rect 2682 12384 2688 12396
rect 2740 12384 2746 12436
rect 3234 12384 3240 12436
rect 3292 12424 3298 12436
rect 3694 12424 3700 12436
rect 3292 12396 3700 12424
rect 3292 12384 3298 12396
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 4065 12427 4123 12433
rect 4065 12424 4077 12427
rect 3936 12396 4077 12424
rect 3936 12384 3942 12396
rect 4065 12393 4077 12396
rect 4111 12393 4123 12427
rect 5534 12424 5540 12436
rect 5495 12396 5540 12424
rect 4065 12387 4123 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 7374 12424 7380 12436
rect 7335 12396 7380 12424
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 8570 12424 8576 12436
rect 8527 12396 8576 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9398 12424 9404 12436
rect 9359 12396 9404 12424
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 10781 12427 10839 12433
rect 10781 12424 10793 12427
rect 10744 12396 10793 12424
rect 10744 12384 10750 12396
rect 10781 12393 10793 12396
rect 10827 12393 10839 12427
rect 10781 12387 10839 12393
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 12345 12427 12403 12433
rect 12345 12424 12357 12427
rect 11848 12396 12357 12424
rect 11848 12384 11854 12396
rect 12345 12393 12357 12396
rect 12391 12393 12403 12427
rect 12345 12387 12403 12393
rect 12894 12384 12900 12436
rect 12952 12424 12958 12436
rect 13449 12427 13507 12433
rect 13449 12424 13461 12427
rect 12952 12396 13461 12424
rect 12952 12384 12958 12396
rect 13449 12393 13461 12396
rect 13495 12393 13507 12427
rect 13449 12387 13507 12393
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 13872 12396 13952 12424
rect 13872 12384 13878 12396
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 4525 12359 4583 12365
rect 4525 12356 4537 12359
rect 3016 12328 4537 12356
rect 3016 12316 3022 12328
rect 4525 12325 4537 12328
rect 4571 12325 4583 12359
rect 4525 12319 4583 12325
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 5905 12359 5963 12365
rect 5905 12356 5917 12359
rect 5500 12328 5917 12356
rect 5500 12316 5506 12328
rect 5905 12325 5917 12328
rect 5951 12356 5963 12359
rect 6822 12356 6828 12368
rect 5951 12328 6828 12356
rect 5951 12325 5963 12328
rect 5905 12319 5963 12325
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 7834 12356 7840 12368
rect 7747 12328 7840 12356
rect 7834 12316 7840 12328
rect 7892 12356 7898 12368
rect 8846 12356 8852 12368
rect 7892 12328 8852 12356
rect 7892 12316 7898 12328
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 10137 12359 10195 12365
rect 10137 12325 10149 12359
rect 10183 12356 10195 12359
rect 10870 12356 10876 12368
rect 10183 12328 10876 12356
rect 10183 12325 10195 12328
rect 10137 12319 10195 12325
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 11330 12356 11336 12368
rect 10980 12328 11336 12356
rect 2314 12248 2320 12300
rect 2372 12288 2378 12300
rect 2590 12288 2596 12300
rect 2372 12260 2596 12288
rect 2372 12248 2378 12260
rect 2590 12248 2596 12260
rect 2648 12288 2654 12300
rect 2777 12291 2835 12297
rect 2777 12288 2789 12291
rect 2648 12260 2789 12288
rect 2648 12248 2654 12260
rect 2777 12257 2789 12260
rect 2823 12257 2835 12291
rect 2777 12251 2835 12257
rect 2869 12291 2927 12297
rect 2869 12257 2881 12291
rect 2915 12288 2927 12291
rect 3050 12288 3056 12300
rect 2915 12260 3056 12288
rect 2915 12257 2927 12260
rect 2869 12251 2927 12257
rect 3050 12248 3056 12260
rect 3108 12248 3114 12300
rect 4430 12288 4436 12300
rect 4391 12260 4436 12288
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 7742 12288 7748 12300
rect 7703 12260 7748 12288
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 10980 12288 11008 12328
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 12986 12356 12992 12368
rect 12947 12328 12992 12356
rect 12986 12316 12992 12328
rect 13044 12316 13050 12368
rect 13924 12365 13952 12396
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 14550 12424 14556 12436
rect 14332 12396 14556 12424
rect 14332 12384 14338 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15470 12384 15476 12436
rect 15528 12424 15534 12436
rect 16758 12424 16764 12436
rect 15528 12396 16764 12424
rect 15528 12384 15534 12396
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 18414 12424 18420 12436
rect 18375 12396 18420 12424
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 18877 12427 18935 12433
rect 18877 12424 18889 12427
rect 18840 12396 18889 12424
rect 18840 12384 18846 12396
rect 18877 12393 18889 12396
rect 18923 12393 18935 12427
rect 18877 12387 18935 12393
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 21266 12424 21272 12436
rect 20763 12396 21272 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21726 12424 21732 12436
rect 21683 12396 21732 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 22738 12424 22744 12436
rect 22699 12396 22744 12424
rect 22738 12384 22744 12396
rect 22796 12384 22802 12436
rect 23750 12384 23756 12436
rect 23808 12424 23814 12436
rect 24762 12424 24768 12436
rect 23808 12396 24768 12424
rect 23808 12384 23814 12396
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 13909 12359 13967 12365
rect 13909 12325 13921 12359
rect 13955 12356 13967 12359
rect 15562 12356 15568 12368
rect 13955 12328 15568 12356
rect 13955 12325 13967 12328
rect 13909 12319 13967 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 16574 12356 16580 12368
rect 15672 12328 16580 12356
rect 10551 12260 11008 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11232 12291 11290 12297
rect 11232 12288 11244 12291
rect 11112 12260 11244 12288
rect 11112 12248 11118 12260
rect 11232 12257 11244 12260
rect 11278 12288 11290 12291
rect 13078 12288 13084 12300
rect 11278 12260 13084 12288
rect 11278 12257 11290 12260
rect 11232 12251 11290 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13722 12248 13728 12300
rect 13780 12288 13786 12300
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13780 12260 13829 12288
rect 13780 12248 13786 12260
rect 13817 12257 13829 12260
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 14550 12248 14556 12300
rect 14608 12288 14614 12300
rect 15672 12297 15700 12328
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 18233 12359 18291 12365
rect 18233 12325 18245 12359
rect 18279 12356 18291 12359
rect 19058 12356 19064 12368
rect 18279 12328 19064 12356
rect 18279 12325 18291 12328
rect 18233 12319 18291 12325
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 23928 12359 23986 12365
rect 23928 12325 23940 12359
rect 23974 12356 23986 12359
rect 24854 12356 24860 12368
rect 23974 12328 24860 12356
rect 23974 12325 23986 12328
rect 23928 12319 23986 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14608 12260 15669 12288
rect 14608 12248 14614 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 15804 12260 16681 12288
rect 15804 12248 15810 12260
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 17092 12260 17233 12288
rect 17092 12248 17098 12260
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 17221 12251 17279 12257
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 17586 12288 17592 12300
rect 17368 12260 17592 12288
rect 17368 12248 17374 12260
rect 17586 12248 17592 12260
rect 17644 12248 17650 12300
rect 18414 12248 18420 12300
rect 18472 12288 18478 12300
rect 18785 12291 18843 12297
rect 18785 12288 18797 12291
rect 18472 12260 18797 12288
rect 18472 12248 18478 12260
rect 18785 12257 18797 12260
rect 18831 12257 18843 12291
rect 21450 12288 21456 12300
rect 21363 12260 21456 12288
rect 18785 12251 18843 12257
rect 21450 12248 21456 12260
rect 21508 12288 21514 12300
rect 21818 12288 21824 12300
rect 21508 12260 21824 12288
rect 21508 12248 21514 12260
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 22557 12291 22615 12297
rect 22557 12257 22569 12291
rect 22603 12288 22615 12291
rect 22922 12288 22928 12300
rect 22603 12260 22928 12288
rect 22603 12257 22615 12260
rect 22557 12251 22615 12257
rect 22922 12248 22928 12260
rect 22980 12248 22986 12300
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 2961 12183 3019 12189
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2976 12152 3004 12183
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7984 12192 8033 12220
rect 7984 12180 7990 12192
rect 8021 12189 8033 12192
rect 8067 12220 8079 12223
rect 8110 12220 8116 12232
rect 8067 12192 8116 12220
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 10962 12220 10968 12232
rect 10836 12192 10968 12220
rect 10836 12180 10842 12192
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 13354 12220 13360 12232
rect 13315 12192 13360 12220
rect 13354 12180 13360 12192
rect 13412 12180 13418 12232
rect 13998 12220 14004 12232
rect 13959 12192 14004 12220
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 15838 12220 15844 12232
rect 15799 12192 15844 12220
rect 15838 12180 15844 12192
rect 15896 12220 15902 12232
rect 16298 12220 16304 12232
rect 15896 12192 16304 12220
rect 15896 12180 15902 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 16816 12192 17417 12220
rect 16816 12180 16822 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 18966 12220 18972 12232
rect 18927 12192 18972 12220
rect 17405 12183 17463 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 2832 12124 3004 12152
rect 2832 12112 2838 12124
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4724 12152 4752 12180
rect 4304 12124 4752 12152
rect 4304 12112 4310 12124
rect 14826 12112 14832 12164
rect 14884 12152 14890 12164
rect 14921 12155 14979 12161
rect 14921 12152 14933 12155
rect 14884 12124 14933 12152
rect 14884 12112 14890 12124
rect 14921 12121 14933 12124
rect 14967 12152 14979 12155
rect 16853 12155 16911 12161
rect 16853 12152 16865 12155
rect 14967 12124 16865 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 16853 12121 16865 12124
rect 16899 12121 16911 12155
rect 16853 12115 16911 12121
rect 2133 12087 2191 12093
rect 2133 12053 2145 12087
rect 2179 12084 2191 12087
rect 2406 12084 2412 12096
rect 2179 12056 2412 12084
rect 2179 12053 2191 12056
rect 2133 12047 2191 12053
rect 2406 12044 2412 12056
rect 2464 12084 2470 12096
rect 2792 12084 2820 12112
rect 5166 12084 5172 12096
rect 2464 12056 2820 12084
rect 5127 12056 5172 12084
rect 2464 12044 2470 12056
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14424 12056 14473 12084
rect 14424 12044 14430 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 16298 12084 16304 12096
rect 16259 12056 16304 12084
rect 14461 12047 14519 12053
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12084 19855 12087
rect 20070 12084 20076 12096
rect 19843 12056 20076 12084
rect 19843 12053 19855 12056
rect 19797 12047 19855 12053
rect 20070 12044 20076 12056
rect 20128 12044 20134 12096
rect 20898 12044 20904 12096
rect 20956 12084 20962 12096
rect 21269 12087 21327 12093
rect 21269 12084 21281 12087
rect 20956 12056 21281 12084
rect 20956 12044 20962 12056
rect 21269 12053 21281 12056
rect 21315 12084 21327 12087
rect 21358 12084 21364 12096
rect 21315 12056 21364 12084
rect 21315 12053 21327 12056
rect 21269 12047 21327 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 23201 12087 23259 12093
rect 23201 12053 23213 12087
rect 23247 12084 23259 12087
rect 23569 12087 23627 12093
rect 23569 12084 23581 12087
rect 23247 12056 23581 12084
rect 23247 12053 23259 12056
rect 23201 12047 23259 12053
rect 23569 12053 23581 12056
rect 23615 12084 23627 12087
rect 23676 12084 23704 12183
rect 23842 12084 23848 12096
rect 23615 12056 23848 12084
rect 23615 12053 23627 12056
rect 23569 12047 23627 12053
rect 23842 12044 23848 12056
rect 23900 12084 23906 12096
rect 24026 12084 24032 12096
rect 23900 12056 24032 12084
rect 23900 12044 23906 12056
rect 24026 12044 24032 12056
rect 24084 12044 24090 12096
rect 25038 12084 25044 12096
rect 24999 12056 25044 12084
rect 25038 12044 25044 12056
rect 25096 12044 25102 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2222 11840 2228 11892
rect 2280 11880 2286 11892
rect 2317 11883 2375 11889
rect 2317 11880 2329 11883
rect 2280 11852 2329 11880
rect 2280 11840 2286 11852
rect 2317 11849 2329 11852
rect 2363 11849 2375 11883
rect 2317 11843 2375 11849
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1670 11676 1676 11688
rect 1443 11648 1676 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1670 11636 1676 11648
rect 1728 11636 1734 11688
rect 2332 11676 2360 11843
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3513 11883 3571 11889
rect 3513 11880 3525 11883
rect 3016 11852 3525 11880
rect 3016 11840 3022 11852
rect 3513 11849 3525 11852
rect 3559 11849 3571 11883
rect 3513 11843 3571 11849
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 4764 11852 5457 11880
rect 4764 11840 4770 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 5445 11843 5503 11849
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7742 11880 7748 11892
rect 7515 11852 7748 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 7834 11840 7840 11892
rect 7892 11880 7898 11892
rect 8110 11880 8116 11892
rect 7892 11852 7937 11880
rect 8071 11852 8116 11880
rect 7892 11840 7898 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 11054 11880 11060 11892
rect 10735 11852 11060 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12492 11852 12537 11880
rect 12492 11840 12498 11852
rect 12802 11840 12808 11892
rect 12860 11880 12866 11892
rect 13814 11880 13820 11892
rect 12860 11852 13820 11880
rect 12860 11840 12866 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14550 11880 14556 11892
rect 14511 11852 14556 11880
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 14936 11852 16129 11880
rect 2590 11772 2596 11824
rect 2648 11812 2654 11824
rect 4065 11815 4123 11821
rect 4065 11812 4077 11815
rect 2648 11784 4077 11812
rect 2648 11772 2654 11784
rect 4065 11781 4077 11784
rect 4111 11781 4123 11815
rect 4065 11775 4123 11781
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 12710 11812 12716 11824
rect 4672 11784 4752 11812
rect 4672 11772 4678 11784
rect 3142 11744 3148 11756
rect 3055 11716 3148 11744
rect 3142 11704 3148 11716
rect 3200 11744 3206 11756
rect 4724 11753 4752 11784
rect 11256 11784 12716 11812
rect 11256 11753 11284 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 3200 11716 4721 11744
rect 3200 11704 3206 11716
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 11241 11747 11299 11753
rect 11241 11744 11253 11747
rect 10367 11716 11253 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 11241 11713 11253 11716
rect 11287 11713 11299 11747
rect 11241 11707 11299 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11698 11744 11704 11756
rect 11388 11716 11704 11744
rect 11388 11704 11394 11716
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 13078 11744 13084 11756
rect 12991 11716 13084 11744
rect 13078 11704 13084 11716
rect 13136 11744 13142 11756
rect 13998 11744 14004 11756
rect 13136 11716 14004 11744
rect 13136 11704 13142 11716
rect 13998 11704 14004 11716
rect 14056 11744 14062 11756
rect 14277 11747 14335 11753
rect 14277 11744 14289 11747
rect 14056 11716 14289 11744
rect 14056 11704 14062 11716
rect 14277 11713 14289 11716
rect 14323 11744 14335 11747
rect 14550 11744 14556 11756
rect 14323 11716 14556 11744
rect 14323 11713 14335 11716
rect 14277 11707 14335 11713
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 2958 11676 2964 11688
rect 2332 11648 2964 11676
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 4430 11636 4436 11688
rect 4488 11676 4494 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 4488 11648 5089 11676
rect 4488 11636 4494 11648
rect 5077 11645 5089 11648
rect 5123 11645 5135 11679
rect 12066 11676 12072 11688
rect 5077 11639 5135 11645
rect 11164 11648 12072 11676
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2590 11608 2596 11620
rect 2087 11580 2596 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2590 11568 2596 11580
rect 2648 11608 2654 11620
rect 2869 11611 2927 11617
rect 2869 11608 2881 11611
rect 2648 11580 2881 11608
rect 2648 11568 2654 11580
rect 2869 11577 2881 11580
rect 2915 11577 2927 11611
rect 4522 11608 4528 11620
rect 4483 11580 4528 11608
rect 2869 11571 2927 11577
rect 4522 11568 4528 11580
rect 4580 11568 4586 11620
rect 11164 11617 11192 11648
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 14936 11685 14964 11852
rect 16117 11849 16129 11852
rect 16163 11880 16175 11883
rect 16298 11880 16304 11892
rect 16163 11852 16304 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16298 11840 16304 11852
rect 16356 11840 16362 11892
rect 18414 11880 18420 11892
rect 18375 11852 18420 11880
rect 18414 11840 18420 11852
rect 18472 11880 18478 11892
rect 21266 11880 21272 11892
rect 18472 11852 18552 11880
rect 21227 11852 21272 11880
rect 18472 11840 18478 11852
rect 15194 11744 15200 11756
rect 15107 11716 15200 11744
rect 15194 11704 15200 11716
rect 15252 11744 15258 11756
rect 16022 11744 16028 11756
rect 15252 11716 16028 11744
rect 15252 11704 15258 11716
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16577 11747 16635 11753
rect 16577 11744 16589 11747
rect 16540 11716 16589 11744
rect 16540 11704 16546 11716
rect 16577 11713 16589 11716
rect 16623 11713 16635 11747
rect 16758 11744 16764 11756
rect 16719 11716 16764 11744
rect 16577 11707 16635 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 18524 11753 18552 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 21542 11880 21548 11892
rect 21503 11852 21548 11880
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 21818 11840 21824 11892
rect 21876 11880 21882 11892
rect 21913 11883 21971 11889
rect 21913 11880 21925 11883
rect 21876 11852 21925 11880
rect 21876 11840 21882 11852
rect 21913 11849 21925 11852
rect 21959 11849 21971 11883
rect 22278 11880 22284 11892
rect 22239 11852 22284 11880
rect 21913 11843 21971 11849
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 22649 11883 22707 11889
rect 22649 11849 22661 11883
rect 22695 11880 22707 11883
rect 23014 11880 23020 11892
rect 22695 11852 23020 11880
rect 22695 11849 22707 11852
rect 22649 11843 22707 11849
rect 23014 11840 23020 11852
rect 23072 11840 23078 11892
rect 23477 11883 23535 11889
rect 23477 11849 23489 11883
rect 23523 11880 23535 11883
rect 23937 11883 23995 11889
rect 23523 11852 23888 11880
rect 23523 11849 23535 11852
rect 23477 11843 23535 11849
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 19518 11744 19524 11756
rect 19479 11716 19524 11744
rect 18509 11707 18567 11713
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 23860 11744 23888 11852
rect 23937 11849 23949 11883
rect 23983 11880 23995 11883
rect 24946 11880 24952 11892
rect 23983 11852 24952 11880
rect 23983 11849 23995 11852
rect 23937 11843 23995 11849
rect 24946 11840 24952 11852
rect 25004 11840 25010 11892
rect 25130 11840 25136 11892
rect 25188 11880 25194 11892
rect 25685 11883 25743 11889
rect 25685 11880 25697 11883
rect 25188 11852 25697 11880
rect 25188 11840 25194 11852
rect 25685 11849 25697 11852
rect 25731 11849 25743 11883
rect 25685 11843 25743 11849
rect 24026 11772 24032 11824
rect 24084 11812 24090 11824
rect 25317 11815 25375 11821
rect 25317 11812 25329 11815
rect 24084 11784 25329 11812
rect 24084 11772 24090 11784
rect 25317 11781 25329 11784
rect 25363 11781 25375 11815
rect 25317 11775 25375 11781
rect 24581 11747 24639 11753
rect 24581 11744 24593 11747
rect 23860 11716 24593 11744
rect 24581 11713 24593 11716
rect 24627 11744 24639 11747
rect 24854 11744 24860 11756
rect 24627 11716 24860 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24854 11704 24860 11716
rect 24912 11704 24918 11756
rect 14921 11679 14979 11685
rect 14921 11645 14933 11679
rect 14967 11645 14979 11679
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 14921 11639 14979 11645
rect 15120 11648 15945 11676
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 11149 11611 11207 11617
rect 11149 11608 11161 11611
rect 9999 11580 11161 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 11149 11577 11161 11580
rect 11195 11577 11207 11611
rect 12805 11611 12863 11617
rect 12805 11608 12817 11611
rect 11149 11571 11207 11577
rect 11808 11580 12817 11608
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 2498 11540 2504 11552
rect 2188 11512 2504 11540
rect 2188 11500 2194 11512
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 3418 11500 3424 11552
rect 3476 11540 3482 11552
rect 3973 11543 4031 11549
rect 3973 11540 3985 11543
rect 3476 11512 3985 11540
rect 3476 11500 3482 11512
rect 3973 11509 3985 11512
rect 4019 11540 4031 11543
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4019 11512 4445 11540
rect 4019 11509 4031 11512
rect 3973 11503 4031 11509
rect 4433 11509 4445 11512
rect 4479 11540 4491 11543
rect 4982 11540 4988 11552
rect 4479 11512 4988 11540
rect 4479 11509 4491 11512
rect 4433 11503 4491 11509
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 11808 11549 11836 11580
rect 12805 11577 12817 11580
rect 12851 11577 12863 11611
rect 12805 11571 12863 11577
rect 13541 11611 13599 11617
rect 13541 11577 13553 11611
rect 13587 11608 13599 11611
rect 13722 11608 13728 11620
rect 13587 11580 13728 11608
rect 13587 11577 13599 11580
rect 13541 11571 13599 11577
rect 13722 11568 13728 11580
rect 13780 11608 13786 11620
rect 13780 11580 14780 11608
rect 13780 11568 13786 11580
rect 11793 11543 11851 11549
rect 11793 11540 11805 11543
rect 11756 11512 11805 11540
rect 11756 11500 11762 11512
rect 11793 11509 11805 11512
rect 11839 11509 11851 11543
rect 11793 11503 11851 11509
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12342 11540 12348 11552
rect 12299 11512 12348 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12342 11500 12348 11512
rect 12400 11540 12406 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12400 11512 12909 11540
rect 12400 11500 12406 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 14752 11540 14780 11580
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14884 11580 15025 11608
rect 14884 11568 14890 11580
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15013 11571 15071 11577
rect 15120 11540 15148 11648
rect 15933 11645 15945 11648
rect 15979 11676 15991 11679
rect 16500 11676 16528 11704
rect 15979 11648 16528 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 21266 11636 21272 11688
rect 21324 11676 21330 11688
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 21324 11648 21373 11676
rect 21324 11636 21330 11648
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 22278 11636 22284 11688
rect 22336 11676 22342 11688
rect 22465 11679 22523 11685
rect 22465 11676 22477 11679
rect 22336 11648 22477 11676
rect 22336 11636 22342 11648
rect 22465 11645 22477 11648
rect 22511 11645 22523 11679
rect 25498 11676 25504 11688
rect 25459 11648 25504 11676
rect 22465 11639 22523 11645
rect 25498 11636 25504 11648
rect 25556 11676 25562 11688
rect 26053 11679 26111 11685
rect 26053 11676 26065 11679
rect 25556 11648 26065 11676
rect 25556 11636 25562 11648
rect 26053 11645 26065 11648
rect 26099 11645 26111 11679
rect 26053 11639 26111 11645
rect 16485 11611 16543 11617
rect 16485 11608 16497 11611
rect 15580 11580 16497 11608
rect 14752 11512 15148 11540
rect 12897 11503 12955 11509
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 15580 11549 15608 11580
rect 16485 11577 16497 11580
rect 16531 11577 16543 11611
rect 16485 11571 16543 11577
rect 17954 11568 17960 11620
rect 18012 11608 18018 11620
rect 19337 11611 19395 11617
rect 19337 11608 19349 11611
rect 18012 11580 19349 11608
rect 18012 11568 18018 11580
rect 19337 11577 19349 11580
rect 19383 11577 19395 11611
rect 19337 11571 19395 11577
rect 24026 11568 24032 11620
rect 24084 11608 24090 11620
rect 24397 11611 24455 11617
rect 24397 11608 24409 11611
rect 24084 11580 24409 11608
rect 24084 11568 24090 11580
rect 24397 11577 24409 11580
rect 24443 11608 24455 11611
rect 24949 11611 25007 11617
rect 24949 11608 24961 11611
rect 24443 11580 24961 11608
rect 24443 11577 24455 11580
rect 24397 11571 24455 11577
rect 24949 11577 24961 11580
rect 24995 11577 25007 11611
rect 24949 11571 25007 11577
rect 15565 11543 15623 11549
rect 15565 11540 15577 11543
rect 15344 11512 15577 11540
rect 15344 11500 15350 11512
rect 15565 11509 15577 11512
rect 15611 11509 15623 11543
rect 15565 11503 15623 11509
rect 17034 11500 17040 11552
rect 17092 11540 17098 11552
rect 17129 11543 17187 11549
rect 17129 11540 17141 11543
rect 17092 11512 17141 11540
rect 17092 11500 17098 11512
rect 17129 11509 17141 11512
rect 17175 11509 17187 11543
rect 17586 11540 17592 11552
rect 17547 11512 17592 11540
rect 17129 11503 17187 11509
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 18969 11543 19027 11549
rect 18969 11540 18981 11543
rect 18840 11512 18981 11540
rect 18840 11500 18846 11512
rect 18969 11509 18981 11512
rect 19015 11509 19027 11543
rect 23014 11540 23020 11552
rect 22975 11512 23020 11540
rect 18969 11503 19027 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 23934 11500 23940 11552
rect 23992 11540 23998 11552
rect 24305 11543 24363 11549
rect 24305 11540 24317 11543
rect 23992 11512 24317 11540
rect 23992 11500 23998 11512
rect 24305 11509 24317 11512
rect 24351 11509 24363 11543
rect 24305 11503 24363 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2406 11336 2412 11348
rect 2367 11308 2412 11336
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 2501 11339 2559 11345
rect 2501 11305 2513 11339
rect 2547 11336 2559 11339
rect 2590 11336 2596 11348
rect 2547 11308 2596 11336
rect 2547 11305 2559 11308
rect 2501 11299 2559 11305
rect 2590 11296 2596 11308
rect 2648 11296 2654 11348
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 2924 11308 3341 11336
rect 2924 11296 2930 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 3697 11339 3755 11345
rect 3697 11336 3709 11339
rect 3660 11308 3709 11336
rect 3660 11296 3666 11308
rect 3697 11305 3709 11308
rect 3743 11305 3755 11339
rect 3697 11299 3755 11305
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4522 11336 4528 11348
rect 4387 11308 4528 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 11057 11339 11115 11345
rect 11057 11305 11069 11339
rect 11103 11336 11115 11339
rect 11698 11336 11704 11348
rect 11103 11308 11704 11336
rect 11103 11305 11115 11308
rect 11057 11299 11115 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 12492 11308 12541 11336
rect 12492 11296 12498 11308
rect 12529 11305 12541 11308
rect 12575 11336 12587 11339
rect 13170 11336 13176 11348
rect 12575 11308 13176 11336
rect 12575 11305 12587 11308
rect 12529 11299 12587 11305
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13814 11296 13820 11348
rect 13872 11336 13878 11348
rect 14001 11339 14059 11345
rect 14001 11336 14013 11339
rect 13872 11308 14013 11336
rect 13872 11296 13878 11308
rect 14001 11305 14013 11308
rect 14047 11336 14059 11339
rect 14274 11336 14280 11348
rect 14047 11308 14280 11336
rect 14047 11305 14059 11308
rect 14001 11299 14059 11305
rect 14274 11296 14280 11308
rect 14332 11296 14338 11348
rect 14737 11339 14795 11345
rect 14737 11305 14749 11339
rect 14783 11336 14795 11339
rect 15194 11336 15200 11348
rect 14783 11308 15200 11336
rect 14783 11305 14795 11308
rect 14737 11299 14795 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 15746 11336 15752 11348
rect 15335 11308 15752 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16850 11336 16856 11348
rect 16811 11308 16856 11336
rect 16850 11296 16856 11308
rect 16908 11296 16914 11348
rect 18601 11339 18659 11345
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 18874 11336 18880 11348
rect 18647 11308 18880 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 20898 11336 20904 11348
rect 20859 11308 20904 11336
rect 20898 11296 20904 11308
rect 20956 11296 20962 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23201 11339 23259 11345
rect 22152 11308 22197 11336
rect 22152 11296 22158 11308
rect 23201 11305 23213 11339
rect 23247 11336 23259 11339
rect 23566 11336 23572 11348
rect 23247 11308 23572 11336
rect 23247 11305 23259 11308
rect 23201 11299 23259 11305
rect 23566 11296 23572 11308
rect 23624 11296 23630 11348
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24765 11339 24823 11345
rect 24765 11336 24777 11339
rect 24176 11308 24777 11336
rect 24176 11296 24182 11308
rect 24765 11305 24777 11308
rect 24811 11305 24823 11339
rect 24765 11299 24823 11305
rect 2961 11271 3019 11277
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 3142 11268 3148 11280
rect 3007 11240 3148 11268
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 3142 11228 3148 11240
rect 3200 11228 3206 11280
rect 11146 11228 11152 11280
rect 11204 11268 11210 11280
rect 11885 11271 11943 11277
rect 11885 11268 11897 11271
rect 11204 11240 11897 11268
rect 11204 11228 11210 11240
rect 11885 11237 11897 11240
rect 11931 11237 11943 11271
rect 13078 11268 13084 11280
rect 13039 11240 13084 11268
rect 11885 11231 11943 11237
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 15105 11271 15163 11277
rect 15105 11237 15117 11271
rect 15151 11268 15163 11271
rect 15838 11268 15844 11280
rect 15151 11240 15844 11268
rect 15151 11237 15163 11240
rect 15105 11231 15163 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 16393 11271 16451 11277
rect 16393 11268 16405 11271
rect 16264 11240 16405 11268
rect 16264 11228 16270 11240
rect 16393 11237 16405 11240
rect 16439 11268 16451 11271
rect 16758 11268 16764 11280
rect 16439 11240 16764 11268
rect 16439 11237 16451 11240
rect 16393 11231 16451 11237
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 18509 11271 18567 11277
rect 18509 11237 18521 11271
rect 18555 11268 18567 11271
rect 18966 11268 18972 11280
rect 18555 11240 18972 11268
rect 18555 11237 18567 11240
rect 18509 11231 18567 11237
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 24486 11268 24492 11280
rect 24136 11240 24492 11268
rect 24136 11212 24164 11240
rect 24486 11228 24492 11240
rect 24544 11228 24550 11280
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 3050 11200 3056 11212
rect 2087 11172 3056 11200
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 12802 11200 12808 11212
rect 12483 11172 12808 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 13541 11203 13599 11209
rect 13541 11169 13553 11203
rect 13587 11200 13599 11203
rect 15654 11200 15660 11212
rect 13587 11172 14320 11200
rect 15615 11172 15660 11200
rect 13587 11169 13599 11172
rect 13541 11163 13599 11169
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3234 11132 3240 11144
rect 2924 11104 3240 11132
rect 2924 11092 2930 11104
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 14292 11141 14320 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 16850 11160 16856 11212
rect 16908 11200 16914 11212
rect 17221 11203 17279 11209
rect 17221 11200 17233 11203
rect 16908 11172 17233 11200
rect 16908 11160 16914 11172
rect 17221 11169 17233 11172
rect 17267 11200 17279 11203
rect 18782 11200 18788 11212
rect 17267 11172 18788 11200
rect 17267 11169 17279 11172
rect 17221 11163 17279 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 21910 11200 21916 11212
rect 21871 11172 21916 11200
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22554 11160 22560 11212
rect 22612 11200 22618 11212
rect 23017 11203 23075 11209
rect 23017 11200 23029 11203
rect 22612 11172 23029 11200
rect 22612 11160 22618 11172
rect 23017 11169 23029 11172
rect 23063 11200 23075 11203
rect 23106 11200 23112 11212
rect 23063 11172 23112 11200
rect 23063 11169 23075 11172
rect 23017 11163 23075 11169
rect 23106 11160 23112 11172
rect 23164 11160 23170 11212
rect 24118 11160 24124 11212
rect 24176 11160 24182 11212
rect 24578 11200 24584 11212
rect 24539 11172 24584 11200
rect 24578 11160 24584 11172
rect 24636 11200 24642 11212
rect 24854 11200 24860 11212
rect 24636 11172 24860 11200
rect 24636 11160 24642 11172
rect 24854 11160 24860 11172
rect 24912 11160 24918 11212
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13872 11104 14105 11132
rect 13872 11092 13878 11104
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 15470 11132 15476 11144
rect 14323 11104 15476 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16022 11132 16028 11144
rect 15979 11104 16028 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 11020 11036 11621 11064
rect 11020 11024 11026 11036
rect 11609 11033 11621 11036
rect 11655 11064 11667 11067
rect 11974 11064 11980 11076
rect 11655 11036 11980 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 13633 11067 13691 11073
rect 13633 11033 13645 11067
rect 13679 11064 13691 11067
rect 15764 11064 15792 11095
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11132 17555 11135
rect 17678 11132 17684 11144
rect 17543 11104 17684 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 17678 11092 17684 11104
rect 17736 11092 17742 11144
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11132 24455 11135
rect 24946 11132 24952 11144
rect 24443 11104 24952 11132
rect 24443 11101 24455 11104
rect 24397 11095 24455 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 16114 11064 16120 11076
rect 13679 11036 16120 11064
rect 13679 11033 13691 11036
rect 13633 11027 13691 11033
rect 16114 11024 16120 11036
rect 16172 11024 16178 11076
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16482 11064 16488 11076
rect 16356 11036 16488 11064
rect 16356 11024 16362 11036
rect 16482 11024 16488 11036
rect 16540 11064 16546 11076
rect 17954 11064 17960 11076
rect 16540 11036 17960 11064
rect 16540 11024 16546 11036
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 10873 10999 10931 11005
rect 10873 10965 10885 10999
rect 10919 10996 10931 10999
rect 11330 10996 11336 11008
rect 10919 10968 11336 10996
rect 10919 10965 10931 10968
rect 10873 10959 10931 10965
rect 11330 10956 11336 10968
rect 11388 10996 11394 11008
rect 14274 10996 14280 11008
rect 11388 10968 14280 10996
rect 11388 10956 11394 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 22554 10956 22560 11008
rect 22612 10996 22618 11008
rect 23934 10996 23940 11008
rect 22612 10968 23940 10996
rect 22612 10956 22618 10968
rect 23934 10956 23940 10968
rect 23992 10956 23998 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 2130 10792 2136 10804
rect 2091 10764 2136 10792
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2314 10752 2320 10804
rect 2372 10792 2378 10804
rect 2409 10795 2467 10801
rect 2409 10792 2421 10795
rect 2372 10764 2421 10792
rect 2372 10752 2378 10764
rect 2409 10761 2421 10764
rect 2455 10761 2467 10795
rect 2409 10755 2467 10761
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 12713 10795 12771 10801
rect 2832 10764 2877 10792
rect 2832 10752 2838 10764
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12802 10792 12808 10804
rect 12759 10764 12808 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13357 10795 13415 10801
rect 13357 10761 13369 10795
rect 13403 10792 13415 10795
rect 13722 10792 13728 10804
rect 13403 10764 13728 10792
rect 13403 10761 13415 10764
rect 13357 10755 13415 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 14792 10764 14841 10792
rect 14792 10752 14798 10764
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15654 10792 15660 10804
rect 15427 10764 15660 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 1673 10727 1731 10733
rect 1673 10693 1685 10727
rect 1719 10724 1731 10727
rect 1946 10724 1952 10736
rect 1719 10696 1952 10724
rect 1719 10693 1731 10696
rect 1673 10687 1731 10693
rect 1946 10684 1952 10696
rect 2004 10724 2010 10736
rect 3145 10727 3203 10733
rect 3145 10724 3157 10727
rect 2004 10696 3157 10724
rect 2004 10684 2010 10696
rect 3145 10693 3157 10696
rect 3191 10693 3203 10727
rect 3145 10687 3203 10693
rect 13633 10727 13691 10733
rect 13633 10693 13645 10727
rect 13679 10724 13691 10727
rect 14642 10724 14648 10736
rect 13679 10696 14648 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 566 10616 572 10668
rect 624 10656 630 10668
rect 5994 10656 6000 10668
rect 624 10628 6000 10656
rect 624 10616 630 10628
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 11793 10659 11851 10665
rect 11793 10625 11805 10659
rect 11839 10656 11851 10659
rect 11882 10656 11888 10668
rect 11839 10628 11888 10656
rect 11839 10625 11851 10628
rect 11793 10619 11851 10625
rect 11882 10616 11888 10628
rect 11940 10656 11946 10668
rect 12710 10656 12716 10668
rect 11940 10628 12716 10656
rect 11940 10616 11946 10628
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 14200 10588 14228 10696
rect 14642 10684 14648 10696
rect 14700 10684 14706 10736
rect 14366 10656 14372 10668
rect 14327 10628 14372 10656
rect 14366 10616 14372 10628
rect 14424 10616 14430 10668
rect 14844 10656 14872 10755
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 16022 10752 16028 10804
rect 16080 10792 16086 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 16080 10764 16405 10792
rect 16080 10752 16086 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 17678 10792 17684 10804
rect 17639 10764 17684 10792
rect 16393 10755 16451 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 21910 10792 21916 10804
rect 21871 10764 21916 10792
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 23106 10792 23112 10804
rect 23067 10764 23112 10792
rect 23106 10752 23112 10764
rect 23164 10752 23170 10804
rect 23658 10752 23664 10804
rect 23716 10792 23722 10804
rect 24765 10795 24823 10801
rect 24765 10792 24777 10795
rect 23716 10764 24777 10792
rect 23716 10752 23722 10764
rect 24765 10761 24777 10764
rect 24811 10761 24823 10795
rect 24765 10755 24823 10761
rect 24854 10752 24860 10804
rect 24912 10792 24918 10804
rect 25133 10795 25191 10801
rect 25133 10792 25145 10795
rect 24912 10764 25145 10792
rect 24912 10752 24918 10764
rect 25133 10761 25145 10764
rect 25179 10761 25191 10795
rect 25133 10755 25191 10761
rect 23934 10684 23940 10736
rect 23992 10724 23998 10736
rect 26142 10724 26148 10736
rect 23992 10696 26148 10724
rect 23992 10684 23998 10696
rect 26142 10684 26148 10696
rect 26200 10684 26206 10736
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 14844 10628 15853 10656
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10656 16083 10659
rect 16206 10656 16212 10668
rect 16071 10628 16212 10656
rect 16071 10625 16083 10628
rect 16025 10619 16083 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 22554 10656 22560 10668
rect 22515 10628 22560 10656
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14200 10560 14289 10588
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 14277 10551 14335 10557
rect 24412 10560 24593 10588
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 13906 10520 13912 10532
rect 12851 10492 13912 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13906 10480 13912 10492
rect 13964 10480 13970 10532
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 14185 10523 14243 10529
rect 14185 10520 14197 10523
rect 14056 10492 14197 10520
rect 14056 10480 14062 10492
rect 14185 10489 14197 10492
rect 14231 10520 14243 10523
rect 15378 10520 15384 10532
rect 14231 10492 15384 10520
rect 14231 10489 14243 10492
rect 14185 10483 14243 10489
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 24412 10464 24440 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 12161 10455 12219 10461
rect 12161 10421 12173 10455
rect 12207 10452 12219 10455
rect 12342 10452 12348 10464
rect 12207 10424 12348 10452
rect 12207 10421 12219 10424
rect 12161 10415 12219 10421
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 13814 10452 13820 10464
rect 13775 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 15746 10452 15752 10464
rect 15335 10424 15752 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17310 10452 17316 10464
rect 17271 10424 17316 10452
rect 17310 10412 17316 10424
rect 17368 10412 17374 10464
rect 24394 10452 24400 10464
rect 24355 10424 24400 10452
rect 24394 10412 24400 10424
rect 24452 10412 24458 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 12618 10208 12624 10260
rect 12676 10248 12682 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 12676 10220 12725 10248
rect 12676 10208 12682 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 12713 10211 12771 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 13228 10220 13273 10248
rect 13228 10208 13234 10220
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 13872 10220 14933 10248
rect 13872 10208 13878 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 15286 10248 15292 10260
rect 15247 10220 15292 10248
rect 14921 10211 14979 10217
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 16114 10248 16120 10260
rect 16075 10220 16120 10248
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 22465 10251 22523 10257
rect 22465 10217 22477 10251
rect 22511 10248 22523 10251
rect 22830 10248 22836 10260
rect 22511 10220 22836 10248
rect 22511 10217 22523 10220
rect 22465 10211 22523 10217
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 24765 10251 24823 10257
rect 24765 10248 24777 10251
rect 24728 10220 24777 10248
rect 24728 10208 24734 10220
rect 24765 10217 24777 10220
rect 24811 10217 24823 10251
rect 24765 10211 24823 10217
rect 13909 10183 13967 10189
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 13998 10180 14004 10192
rect 13955 10152 14004 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 13998 10140 14004 10152
rect 14056 10140 14062 10192
rect 15841 10183 15899 10189
rect 15841 10149 15853 10183
rect 15887 10180 15899 10183
rect 16206 10180 16212 10192
rect 15887 10152 16212 10180
rect 15887 10149 15899 10152
rect 15841 10143 15899 10149
rect 16206 10140 16212 10152
rect 16264 10140 16270 10192
rect 14274 10112 14280 10124
rect 14187 10084 14280 10112
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 17678 10112 17684 10124
rect 14332 10084 17684 10112
rect 14332 10072 14338 10084
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 23474 10112 23480 10124
rect 23435 10084 23480 10112
rect 23474 10072 23480 10084
rect 23532 10072 23538 10124
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 23808 10084 24593 10112
rect 23808 10072 23814 10084
rect 24581 10081 24593 10084
rect 24627 10112 24639 10115
rect 24946 10112 24952 10124
rect 24627 10084 24952 10112
rect 24627 10081 24639 10084
rect 24581 10075 24639 10081
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 13357 10047 13415 10053
rect 13357 10013 13369 10047
rect 13403 10044 13415 10047
rect 13630 10044 13636 10056
rect 13403 10016 13636 10044
rect 13403 10013 13415 10016
rect 13357 10007 13415 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13998 9936 14004 9988
rect 14056 9976 14062 9988
rect 14366 9976 14372 9988
rect 14056 9948 14372 9976
rect 14056 9936 14062 9948
rect 14366 9936 14372 9948
rect 14424 9976 14430 9988
rect 14553 9979 14611 9985
rect 14553 9976 14565 9979
rect 14424 9948 14565 9976
rect 14424 9936 14430 9948
rect 14553 9945 14565 9948
rect 14599 9945 14611 9979
rect 14553 9939 14611 9945
rect 23661 9979 23719 9985
rect 23661 9945 23673 9979
rect 23707 9976 23719 9979
rect 25774 9976 25780 9988
rect 23707 9948 25780 9976
rect 23707 9945 23719 9948
rect 23661 9939 23719 9945
rect 25774 9936 25780 9948
rect 25832 9936 25838 9988
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13449 9707 13507 9713
rect 13449 9704 13461 9707
rect 13136 9676 13461 9704
rect 13136 9664 13142 9676
rect 13449 9673 13461 9676
rect 13495 9673 13507 9707
rect 13449 9667 13507 9673
rect 15381 9707 15439 9713
rect 15381 9673 15393 9707
rect 15427 9704 15439 9707
rect 15654 9704 15660 9716
rect 15427 9676 15660 9704
rect 15427 9673 15439 9676
rect 15381 9667 15439 9673
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 23750 9664 23756 9716
rect 23808 9704 23814 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23808 9676 23857 9704
rect 23808 9664 23814 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 24946 9704 24952 9716
rect 23845 9667 23903 9673
rect 24780 9676 24952 9704
rect 12805 9639 12863 9645
rect 12805 9605 12817 9639
rect 12851 9636 12863 9639
rect 13630 9636 13636 9648
rect 12851 9608 13636 9636
rect 12851 9605 12863 9608
rect 12805 9599 12863 9605
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 14182 9636 14188 9648
rect 14143 9608 14188 9636
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 15749 9639 15807 9645
rect 14332 9608 14780 9636
rect 14332 9596 14338 9608
rect 13170 9568 13176 9580
rect 13131 9540 13176 9568
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 14090 9568 14096 9580
rect 14051 9540 14096 9568
rect 14090 9528 14096 9540
rect 14148 9568 14154 9580
rect 14752 9577 14780 9608
rect 15749 9605 15761 9639
rect 15795 9636 15807 9639
rect 16482 9636 16488 9648
rect 15795 9608 16488 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 16482 9596 16488 9608
rect 16540 9596 16546 9648
rect 24780 9636 24808 9676
rect 24946 9664 24952 9676
rect 25004 9664 25010 9716
rect 25133 9639 25191 9645
rect 25133 9636 25145 9639
rect 24780 9608 25145 9636
rect 25133 9605 25145 9608
rect 25179 9605 25191 9639
rect 25133 9599 25191 9605
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 14148 9540 14657 9568
rect 14148 9528 14154 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 14645 9531 14703 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9537 14795 9571
rect 14737 9531 14795 9537
rect 22738 9528 22744 9580
rect 22796 9568 22802 9580
rect 23750 9568 23756 9580
rect 22796 9540 23756 9568
rect 22796 9528 22802 9540
rect 23750 9528 23756 9540
rect 23808 9528 23814 9580
rect 24394 9568 24400 9580
rect 24355 9540 24400 9568
rect 24394 9528 24400 9540
rect 24452 9528 24458 9580
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14553 9503 14611 9509
rect 14553 9500 14565 9503
rect 13964 9472 14565 9500
rect 13964 9460 13970 9472
rect 14553 9469 14565 9472
rect 14599 9469 14611 9503
rect 24412 9500 24440 9528
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 24412 9472 24593 9500
rect 14553 9463 14611 9469
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 23934 9324 23940 9376
rect 23992 9364 23998 9376
rect 24765 9367 24823 9373
rect 24765 9364 24777 9367
rect 23992 9336 24777 9364
rect 23992 9324 23998 9336
rect 24765 9333 24777 9336
rect 24811 9333 24823 9367
rect 24765 9327 24823 9333
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 13964 9132 14197 9160
rect 13964 9120 13970 9132
rect 14185 9129 14197 9132
rect 14231 9129 14243 9163
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 14185 9123 14243 9129
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24946 9024 24952 9036
rect 24627 8996 24952 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24946 8984 24952 8996
rect 25004 9024 25010 9036
rect 25406 9024 25412 9036
rect 25004 8996 25412 9024
rect 25004 8984 25010 8996
rect 25406 8984 25412 8996
rect 25464 8984 25470 9036
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 24118 8616 24124 8628
rect 24079 8588 24124 8616
rect 24118 8576 24124 8588
rect 24176 8576 24182 8628
rect 24946 8616 24952 8628
rect 24907 8588 24952 8616
rect 24946 8576 24952 8588
rect 25004 8576 25010 8628
rect 19978 8508 19984 8560
rect 20036 8548 20042 8560
rect 24670 8548 24676 8560
rect 20036 8520 24676 8548
rect 20036 8508 20042 8520
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 23934 8412 23940 8424
rect 23895 8384 23940 8412
rect 23934 8372 23940 8384
rect 23992 8412 23998 8424
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 23992 8384 24501 8412
rect 23992 8372 23998 8384
rect 24489 8381 24501 8384
rect 24535 8381 24547 8415
rect 24489 8375 24547 8381
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 24670 5896 24676 5908
rect 24631 5868 24676 5896
rect 24670 5856 24676 5868
rect 24728 5856 24734 5908
rect 24486 5760 24492 5772
rect 24447 5732 24492 5760
rect 24486 5720 24492 5732
rect 24544 5720 24550 5772
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 24581 5355 24639 5361
rect 24581 5321 24593 5355
rect 24627 5352 24639 5355
rect 24670 5352 24676 5364
rect 24627 5324 24676 5352
rect 24627 5321 24639 5324
rect 24581 5315 24639 5321
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 24026 4768 24032 4820
rect 24084 4808 24090 4820
rect 24121 4811 24179 4817
rect 24121 4808 24133 4811
rect 24084 4780 24133 4808
rect 24084 4768 24090 4780
rect 24121 4777 24133 4780
rect 24167 4777 24179 4811
rect 24121 4771 24179 4777
rect 24581 4743 24639 4749
rect 24581 4709 24593 4743
rect 24627 4740 24639 4743
rect 24670 4740 24676 4752
rect 24627 4712 24676 4740
rect 24627 4709 24639 4712
rect 24581 4703 24639 4709
rect 24670 4700 24676 4712
rect 24728 4700 24734 4752
rect 24486 4672 24492 4684
rect 24447 4644 24492 4672
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 24210 4564 24216 4616
rect 24268 4604 24274 4616
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 24268 4576 24685 4604
rect 24268 4564 24274 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 24118 4264 24124 4276
rect 24079 4236 24124 4264
rect 24118 4224 24124 4236
rect 24176 4224 24182 4276
rect 24210 4156 24216 4208
rect 24268 4196 24274 4208
rect 24268 4168 24808 4196
rect 24268 4156 24274 4168
rect 24780 4128 24808 4168
rect 24857 4131 24915 4137
rect 24857 4128 24869 4131
rect 24780 4100 24869 4128
rect 24857 4097 24869 4100
rect 24903 4097 24915 4131
rect 24857 4091 24915 4097
rect 24578 3924 24584 3936
rect 24539 3896 24584 3924
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 11974 2632 11980 2644
rect 11935 2604 11980 2632
rect 11974 2592 11980 2604
rect 12032 2592 12038 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 13998 2632 14004 2644
rect 12492 2604 12537 2632
rect 13959 2604 14004 2632
rect 12492 2592 12498 2604
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 11992 2496 12020 2592
rect 12452 2564 12480 2592
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12452 2536 12878 2564
rect 12866 2533 12878 2536
rect 12912 2533 12924 2567
rect 12866 2527 12924 2533
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 11992 2468 12633 2496
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 18371 2468 19012 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 18506 2360 18512 2372
rect 18467 2332 18512 2360
rect 18506 2320 18512 2332
rect 18564 2320 18570 2372
rect 18984 2301 19012 2468
rect 18969 2295 19027 2301
rect 18969 2261 18981 2295
rect 19015 2292 19027 2295
rect 19518 2292 19524 2304
rect 19015 2264 19524 2292
rect 19015 2261 19027 2264
rect 18969 2255 19027 2261
rect 19518 2252 19524 2264
rect 19576 2252 19582 2304
rect 24213 2295 24271 2301
rect 24213 2261 24225 2295
rect 24259 2292 24271 2295
rect 25130 2292 25136 2304
rect 24259 2264 25136 2292
rect 24259 2261 24271 2264
rect 24213 2255 24271 2261
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 3332 26256 3384 26308
rect 4896 26256 4948 26308
rect 12992 25780 13044 25832
rect 20904 25780 20956 25832
rect 11612 25712 11664 25764
rect 20352 25712 20404 25764
rect 3056 25644 3108 25696
rect 7840 25644 7892 25696
rect 9496 25644 9548 25696
rect 22928 25644 22980 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 4160 25440 4212 25492
rect 7656 25440 7708 25492
rect 11612 25483 11664 25492
rect 11612 25449 11621 25483
rect 11621 25449 11655 25483
rect 11655 25449 11664 25483
rect 11612 25440 11664 25449
rect 16488 25440 16540 25492
rect 17040 25440 17092 25492
rect 27620 25440 27672 25492
rect 7472 25372 7524 25424
rect 2228 25304 2280 25356
rect 3516 25304 3568 25356
rect 5080 25304 5132 25356
rect 6276 25236 6328 25288
rect 7840 25372 7892 25424
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 11336 25304 11388 25356
rect 12716 25347 12768 25356
rect 12716 25313 12725 25347
rect 12725 25313 12759 25347
rect 12759 25313 12768 25347
rect 12716 25304 12768 25313
rect 14096 25304 14148 25356
rect 14280 25347 14332 25356
rect 14280 25313 14289 25347
rect 14289 25313 14323 25347
rect 14323 25313 14332 25347
rect 14280 25304 14332 25313
rect 14004 25236 14056 25288
rect 2780 25168 2832 25220
rect 1584 25143 1636 25152
rect 1584 25109 1593 25143
rect 1593 25109 1627 25143
rect 1627 25109 1636 25143
rect 1584 25100 1636 25109
rect 1676 25100 1728 25152
rect 2964 25100 3016 25152
rect 9128 25100 9180 25152
rect 12992 25168 13044 25220
rect 13360 25143 13412 25152
rect 13360 25109 13369 25143
rect 13369 25109 13403 25143
rect 13403 25109 13412 25143
rect 13360 25100 13412 25109
rect 13820 25143 13872 25152
rect 13820 25109 13829 25143
rect 13829 25109 13863 25143
rect 13863 25109 13872 25143
rect 13820 25100 13872 25109
rect 24308 25372 24360 25424
rect 16396 25304 16448 25356
rect 17868 25304 17920 25356
rect 19156 25304 19208 25356
rect 20444 25304 20496 25356
rect 21548 25347 21600 25356
rect 21548 25313 21557 25347
rect 21557 25313 21591 25347
rect 21591 25313 21600 25347
rect 21548 25304 21600 25313
rect 25044 25304 25096 25356
rect 16212 25279 16264 25288
rect 16212 25245 16221 25279
rect 16221 25245 16255 25279
rect 16255 25245 16264 25279
rect 16212 25236 16264 25245
rect 18880 25279 18932 25288
rect 15936 25168 15988 25220
rect 16764 25168 16816 25220
rect 18604 25168 18656 25220
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 21180 25236 21232 25288
rect 23020 25236 23072 25288
rect 18972 25168 19024 25220
rect 24768 25211 24820 25220
rect 14832 25143 14884 25152
rect 14832 25109 14841 25143
rect 14841 25109 14875 25143
rect 14875 25109 14884 25143
rect 14832 25100 14884 25109
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 17040 25100 17092 25152
rect 20076 25100 20128 25152
rect 21088 25100 21140 25152
rect 24768 25177 24777 25211
rect 24777 25177 24811 25211
rect 24811 25177 24820 25211
rect 24768 25168 24820 25177
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3792 24939 3844 24948
rect 3792 24905 3801 24939
rect 3801 24905 3835 24939
rect 3835 24905 3844 24939
rect 3792 24896 3844 24905
rect 4896 24939 4948 24948
rect 4896 24905 4905 24939
rect 4905 24905 4939 24939
rect 4939 24905 4948 24939
rect 4896 24896 4948 24905
rect 12256 24939 12308 24948
rect 12256 24905 12265 24939
rect 12265 24905 12299 24939
rect 12299 24905 12308 24939
rect 12256 24896 12308 24905
rect 2044 24692 2096 24744
rect 3424 24692 3476 24744
rect 4896 24760 4948 24812
rect 7656 24828 7708 24880
rect 9128 24828 9180 24880
rect 8208 24624 8260 24676
rect 12532 24760 12584 24812
rect 13544 24760 13596 24812
rect 18788 24896 18840 24948
rect 21548 24896 21600 24948
rect 24676 24896 24728 24948
rect 15752 24828 15804 24880
rect 20904 24828 20956 24880
rect 21088 24828 21140 24880
rect 14464 24760 14516 24812
rect 16764 24803 16816 24812
rect 16764 24769 16773 24803
rect 16773 24769 16807 24803
rect 16807 24769 16816 24803
rect 16764 24760 16816 24769
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 20352 24760 20404 24812
rect 20996 24760 21048 24812
rect 21916 24828 21968 24880
rect 22100 24760 22152 24812
rect 22744 24760 22796 24812
rect 9588 24692 9640 24744
rect 9496 24624 9548 24676
rect 1400 24556 1452 24608
rect 1676 24556 1728 24608
rect 2228 24556 2280 24608
rect 2688 24599 2740 24608
rect 2688 24565 2697 24599
rect 2697 24565 2731 24599
rect 2731 24565 2740 24599
rect 2688 24556 2740 24565
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 4712 24556 4764 24608
rect 5080 24556 5132 24608
rect 6276 24556 6328 24608
rect 7472 24556 7524 24608
rect 7656 24599 7708 24608
rect 7656 24565 7665 24599
rect 7665 24565 7699 24599
rect 7699 24565 7708 24599
rect 7656 24556 7708 24565
rect 8116 24599 8168 24608
rect 8116 24565 8125 24599
rect 8125 24565 8159 24599
rect 8159 24565 8168 24599
rect 8116 24556 8168 24565
rect 8760 24599 8812 24608
rect 8760 24565 8769 24599
rect 8769 24565 8803 24599
rect 8803 24565 8812 24599
rect 8760 24556 8812 24565
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 10324 24624 10376 24676
rect 10784 24624 10836 24676
rect 12072 24624 12124 24676
rect 13360 24692 13412 24744
rect 15844 24692 15896 24744
rect 17684 24692 17736 24744
rect 18972 24692 19024 24744
rect 21180 24692 21232 24744
rect 22192 24692 22244 24744
rect 23204 24692 23256 24744
rect 14832 24624 14884 24676
rect 16396 24624 16448 24676
rect 19156 24667 19208 24676
rect 19156 24633 19165 24667
rect 19165 24633 19199 24667
rect 19199 24633 19208 24667
rect 19156 24624 19208 24633
rect 20168 24624 20220 24676
rect 10692 24599 10744 24608
rect 10692 24565 10701 24599
rect 10701 24565 10735 24599
rect 10735 24565 10744 24599
rect 10692 24556 10744 24565
rect 11152 24599 11204 24608
rect 11152 24565 11161 24599
rect 11161 24565 11195 24599
rect 11195 24565 11204 24599
rect 11152 24556 11204 24565
rect 11428 24599 11480 24608
rect 11428 24565 11437 24599
rect 11437 24565 11471 24599
rect 11471 24565 11480 24599
rect 11428 24556 11480 24565
rect 12716 24556 12768 24608
rect 13360 24556 13412 24608
rect 13452 24556 13504 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 14280 24556 14332 24608
rect 14556 24556 14608 24608
rect 14740 24556 14792 24608
rect 15844 24556 15896 24608
rect 16120 24556 16172 24608
rect 16304 24556 16356 24608
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 17868 24556 17920 24608
rect 18972 24556 19024 24608
rect 19524 24556 19576 24608
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 20996 24556 21048 24608
rect 21364 24556 21416 24608
rect 23020 24599 23072 24608
rect 23020 24565 23029 24599
rect 23029 24565 23063 24599
rect 23063 24565 23072 24599
rect 23020 24556 23072 24565
rect 23204 24556 23256 24608
rect 23480 24556 23532 24608
rect 24860 24556 24912 24608
rect 25044 24556 25096 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 296 24352 348 24404
rect 1308 24352 1360 24404
rect 4160 24352 4212 24404
rect 6368 24352 6420 24404
rect 8116 24352 8168 24404
rect 9680 24395 9732 24404
rect 9680 24361 9689 24395
rect 9689 24361 9723 24395
rect 9723 24361 9732 24395
rect 9680 24352 9732 24361
rect 14004 24395 14056 24404
rect 14004 24361 14013 24395
rect 14013 24361 14047 24395
rect 14047 24361 14056 24395
rect 14004 24352 14056 24361
rect 18420 24352 18472 24404
rect 18880 24352 18932 24404
rect 20168 24395 20220 24404
rect 20168 24361 20177 24395
rect 20177 24361 20211 24395
rect 20211 24361 20220 24395
rect 20168 24352 20220 24361
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 24952 24352 25004 24404
rect 25964 24352 26016 24404
rect 9588 24284 9640 24336
rect 17684 24284 17736 24336
rect 21824 24284 21876 24336
rect 22284 24284 22336 24336
rect 1952 24216 2004 24268
rect 2504 24259 2556 24268
rect 2504 24225 2513 24259
rect 2513 24225 2547 24259
rect 2547 24225 2556 24259
rect 2504 24216 2556 24225
rect 3792 24216 3844 24268
rect 6368 24216 6420 24268
rect 8484 24259 8536 24268
rect 8484 24225 8493 24259
rect 8493 24225 8527 24259
rect 8527 24225 8536 24259
rect 8484 24216 8536 24225
rect 9864 24216 9916 24268
rect 2044 24191 2096 24200
rect 2044 24157 2053 24191
rect 2053 24157 2087 24191
rect 2087 24157 2096 24191
rect 2044 24148 2096 24157
rect 1492 24012 1544 24064
rect 2780 24012 2832 24064
rect 3608 24012 3660 24064
rect 4160 24012 4212 24064
rect 5264 24055 5316 24064
rect 5264 24021 5273 24055
rect 5273 24021 5307 24055
rect 5307 24021 5316 24055
rect 5264 24012 5316 24021
rect 9956 24148 10008 24200
rect 11520 24191 11572 24200
rect 10048 24080 10100 24132
rect 11520 24157 11529 24191
rect 11529 24157 11563 24191
rect 11563 24157 11572 24191
rect 11520 24148 11572 24157
rect 6092 24012 6144 24064
rect 6828 24012 6880 24064
rect 8208 24012 8260 24064
rect 8668 24055 8720 24064
rect 8668 24021 8677 24055
rect 8677 24021 8711 24055
rect 8711 24021 8720 24055
rect 8668 24012 8720 24021
rect 11060 24055 11112 24064
rect 11060 24021 11069 24055
rect 11069 24021 11103 24055
rect 11103 24021 11112 24055
rect 11060 24012 11112 24021
rect 13360 24216 13412 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 16672 24216 16724 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 20720 24216 20772 24268
rect 23020 24259 23072 24268
rect 23020 24225 23029 24259
rect 23029 24225 23063 24259
rect 23063 24225 23072 24259
rect 23020 24216 23072 24225
rect 24124 24216 24176 24268
rect 12808 24080 12860 24132
rect 12992 24080 13044 24132
rect 12348 24012 12400 24064
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 14648 24148 14700 24200
rect 15476 24191 15528 24200
rect 15476 24157 15485 24191
rect 15485 24157 15519 24191
rect 15519 24157 15528 24191
rect 15476 24148 15528 24157
rect 16580 24191 16632 24200
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 18972 24191 19024 24200
rect 18972 24157 18981 24191
rect 18981 24157 19015 24191
rect 19015 24157 19024 24191
rect 18972 24148 19024 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 21640 24191 21692 24200
rect 21640 24157 21649 24191
rect 21649 24157 21683 24191
rect 21683 24157 21692 24191
rect 23204 24191 23256 24200
rect 21640 24148 21692 24157
rect 23204 24157 23213 24191
rect 23213 24157 23247 24191
rect 23247 24157 23256 24191
rect 23204 24148 23256 24157
rect 21272 24080 21324 24132
rect 22652 24123 22704 24132
rect 22652 24089 22661 24123
rect 22661 24089 22695 24123
rect 22695 24089 22704 24123
rect 22652 24080 22704 24089
rect 14004 24055 14056 24064
rect 14004 24021 14013 24055
rect 14013 24021 14047 24055
rect 14047 24021 14056 24055
rect 14004 24012 14056 24021
rect 14464 24012 14516 24064
rect 14740 24012 14792 24064
rect 15568 24012 15620 24064
rect 16212 24012 16264 24064
rect 16304 24012 16356 24064
rect 17960 24055 18012 24064
rect 17960 24021 17969 24055
rect 17969 24021 18003 24055
rect 18003 24021 18012 24055
rect 17960 24012 18012 24021
rect 19064 24055 19116 24064
rect 19064 24021 19073 24055
rect 19073 24021 19107 24055
rect 19107 24021 19116 24055
rect 19064 24012 19116 24021
rect 20444 24055 20496 24064
rect 20444 24021 20453 24055
rect 20453 24021 20487 24055
rect 20487 24021 20496 24055
rect 20444 24012 20496 24021
rect 21364 24012 21416 24064
rect 23664 24055 23716 24064
rect 23664 24021 23673 24055
rect 23673 24021 23707 24055
rect 23707 24021 23716 24055
rect 23664 24012 23716 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 2504 23851 2556 23860
rect 2504 23817 2513 23851
rect 2513 23817 2547 23851
rect 2547 23817 2556 23851
rect 2504 23808 2556 23817
rect 2964 23851 3016 23860
rect 2964 23817 2973 23851
rect 2973 23817 3007 23851
rect 3007 23817 3016 23851
rect 2964 23808 3016 23817
rect 3976 23808 4028 23860
rect 4528 23740 4580 23792
rect 3792 23672 3844 23724
rect 4160 23715 4212 23724
rect 4160 23681 4169 23715
rect 4169 23681 4203 23715
rect 4203 23681 4212 23715
rect 4160 23672 4212 23681
rect 5632 23672 5684 23724
rect 6368 23808 6420 23860
rect 9036 23808 9088 23860
rect 11336 23808 11388 23860
rect 13820 23808 13872 23860
rect 8300 23740 8352 23792
rect 8760 23672 8812 23724
rect 10784 23672 10836 23724
rect 2964 23604 3016 23656
rect 3976 23647 4028 23656
rect 3976 23613 3985 23647
rect 3985 23613 4019 23647
rect 4019 23613 4028 23647
rect 3976 23604 4028 23613
rect 6092 23604 6144 23656
rect 7656 23604 7708 23656
rect 8024 23604 8076 23656
rect 9680 23604 9732 23656
rect 11060 23647 11112 23656
rect 11060 23613 11069 23647
rect 11069 23613 11103 23647
rect 11103 23613 11112 23647
rect 11060 23604 11112 23613
rect 3516 23536 3568 23588
rect 6368 23536 6420 23588
rect 7840 23536 7892 23588
rect 9864 23536 9916 23588
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 15292 23808 15344 23860
rect 16672 23851 16724 23860
rect 16672 23817 16681 23851
rect 16681 23817 16715 23851
rect 16715 23817 16724 23851
rect 16672 23808 16724 23817
rect 17040 23851 17092 23860
rect 17040 23817 17049 23851
rect 17049 23817 17083 23851
rect 17083 23817 17092 23851
rect 17040 23808 17092 23817
rect 17500 23851 17552 23860
rect 17500 23817 17509 23851
rect 17509 23817 17543 23851
rect 17543 23817 17552 23851
rect 17500 23808 17552 23817
rect 19616 23808 19668 23860
rect 21824 23808 21876 23860
rect 22284 23851 22336 23860
rect 22284 23817 22293 23851
rect 22293 23817 22327 23851
rect 22327 23817 22336 23851
rect 22284 23808 22336 23817
rect 22836 23808 22888 23860
rect 24124 23808 24176 23860
rect 25136 23851 25188 23860
rect 25136 23817 25145 23851
rect 25145 23817 25179 23851
rect 25179 23817 25188 23851
rect 25136 23808 25188 23817
rect 20720 23783 20772 23792
rect 20720 23749 20729 23783
rect 20729 23749 20763 23783
rect 20763 23749 20772 23783
rect 20720 23740 20772 23749
rect 16672 23672 16724 23724
rect 22008 23672 22060 23724
rect 12440 23604 12492 23613
rect 18052 23604 18104 23656
rect 20904 23604 20956 23656
rect 21088 23604 21140 23656
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 22468 23647 22520 23656
rect 22468 23613 22477 23647
rect 22477 23613 22511 23647
rect 22511 23613 22520 23647
rect 22468 23604 22520 23613
rect 23664 23740 23716 23792
rect 24860 23604 24912 23656
rect 1952 23468 2004 23520
rect 3700 23468 3752 23520
rect 5172 23511 5224 23520
rect 5172 23477 5181 23511
rect 5181 23477 5215 23511
rect 5215 23477 5224 23511
rect 5172 23468 5224 23477
rect 5264 23468 5316 23520
rect 6828 23468 6880 23520
rect 7380 23468 7432 23520
rect 9036 23468 9088 23520
rect 9956 23468 10008 23520
rect 12808 23536 12860 23588
rect 14188 23536 14240 23588
rect 15660 23536 15712 23588
rect 17040 23536 17092 23588
rect 17960 23536 18012 23588
rect 18972 23536 19024 23588
rect 21364 23579 21416 23588
rect 21364 23545 21373 23579
rect 21373 23545 21407 23579
rect 21407 23545 21416 23579
rect 21364 23536 21416 23545
rect 23480 23536 23532 23588
rect 12992 23468 13044 23520
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 15476 23511 15528 23520
rect 15476 23477 15485 23511
rect 15485 23477 15519 23511
rect 15519 23477 15528 23511
rect 15476 23468 15528 23477
rect 23020 23468 23072 23520
rect 23848 23468 23900 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5632 23307 5684 23316
rect 5632 23273 5641 23307
rect 5641 23273 5675 23307
rect 5675 23273 5684 23307
rect 5632 23264 5684 23273
rect 6092 23264 6144 23316
rect 7288 23264 7340 23316
rect 9588 23264 9640 23316
rect 3700 23239 3752 23248
rect 3700 23205 3709 23239
rect 3709 23205 3743 23239
rect 3743 23205 3752 23239
rect 3700 23196 3752 23205
rect 4252 23196 4304 23248
rect 8576 23239 8628 23248
rect 8576 23205 8585 23239
rect 8585 23205 8619 23239
rect 8619 23205 8628 23239
rect 8576 23196 8628 23205
rect 10968 23264 11020 23316
rect 13360 23307 13412 23316
rect 13360 23273 13369 23307
rect 13369 23273 13403 23307
rect 13403 23273 13412 23307
rect 13360 23264 13412 23273
rect 16672 23264 16724 23316
rect 19524 23264 19576 23316
rect 22100 23264 22152 23316
rect 22376 23264 22428 23316
rect 23664 23307 23716 23316
rect 23664 23273 23673 23307
rect 23673 23273 23707 23307
rect 23707 23273 23716 23307
rect 23664 23264 23716 23273
rect 25688 23264 25740 23316
rect 10232 23239 10284 23248
rect 10232 23205 10241 23239
rect 10241 23205 10275 23239
rect 10275 23205 10284 23239
rect 10232 23196 10284 23205
rect 10324 23196 10376 23248
rect 2596 23171 2648 23180
rect 2596 23137 2605 23171
rect 2605 23137 2639 23171
rect 2639 23137 2648 23171
rect 2596 23128 2648 23137
rect 3332 23128 3384 23180
rect 6552 23128 6604 23180
rect 8668 23128 8720 23180
rect 1768 23103 1820 23112
rect 1768 23069 1777 23103
rect 1777 23069 1811 23103
rect 1811 23069 1820 23103
rect 1768 23060 1820 23069
rect 2964 23060 3016 23112
rect 6644 23060 6696 23112
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 8208 23103 8260 23112
rect 8208 23069 8217 23103
rect 8217 23069 8251 23103
rect 8251 23069 8260 23103
rect 8208 23060 8260 23069
rect 9864 23060 9916 23112
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10324 23060 10376 23069
rect 11888 23196 11940 23248
rect 12256 23196 12308 23248
rect 12716 23196 12768 23248
rect 13912 23171 13964 23180
rect 13912 23137 13921 23171
rect 13921 23137 13955 23171
rect 13955 23137 13964 23171
rect 13912 23128 13964 23137
rect 16580 23196 16632 23248
rect 15660 23171 15712 23180
rect 15660 23137 15694 23171
rect 15694 23137 15712 23171
rect 15660 23128 15712 23137
rect 16856 23128 16908 23180
rect 17960 23171 18012 23180
rect 17960 23137 17969 23171
rect 17969 23137 18003 23171
rect 18003 23137 18012 23171
rect 17960 23128 18012 23137
rect 19064 23128 19116 23180
rect 19616 23171 19668 23180
rect 19616 23137 19625 23171
rect 19625 23137 19659 23171
rect 19659 23137 19668 23171
rect 19616 23128 19668 23137
rect 6736 23035 6788 23044
rect 6736 23001 6745 23035
rect 6745 23001 6779 23035
rect 6779 23001 6788 23035
rect 6736 22992 6788 23001
rect 2412 22924 2464 22976
rect 2872 22924 2924 22976
rect 6552 22967 6604 22976
rect 6552 22933 6561 22967
rect 6561 22933 6595 22967
rect 6595 22933 6604 22967
rect 6552 22924 6604 22933
rect 9404 22967 9456 22976
rect 9404 22933 9413 22967
rect 9413 22933 9447 22967
rect 9447 22933 9456 22967
rect 9404 22924 9456 22933
rect 9864 22967 9916 22976
rect 9864 22933 9873 22967
rect 9873 22933 9907 22967
rect 9907 22933 9916 22967
rect 9864 22924 9916 22933
rect 10968 22967 11020 22976
rect 10968 22933 10977 22967
rect 10977 22933 11011 22967
rect 11011 22933 11020 22967
rect 10968 22924 11020 22933
rect 11152 22924 11204 22976
rect 18144 23103 18196 23112
rect 18144 23069 18153 23103
rect 18153 23069 18187 23103
rect 18187 23069 18196 23103
rect 18144 23060 18196 23069
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20260 23128 20312 23180
rect 21640 23196 21692 23248
rect 21916 23196 21968 23248
rect 23112 23128 23164 23180
rect 25780 23128 25832 23180
rect 19892 23060 19944 23112
rect 20904 23060 20956 23112
rect 23664 23060 23716 23112
rect 24124 23103 24176 23112
rect 24124 23069 24133 23103
rect 24133 23069 24167 23103
rect 24167 23069 24176 23103
rect 24124 23060 24176 23069
rect 24216 23103 24268 23112
rect 24216 23069 24225 23103
rect 24225 23069 24259 23103
rect 24259 23069 24268 23103
rect 24216 23060 24268 23069
rect 19156 22992 19208 23044
rect 19432 22992 19484 23044
rect 12440 22924 12492 22976
rect 12808 22967 12860 22976
rect 12808 22933 12817 22967
rect 12817 22933 12851 22967
rect 12851 22933 12860 22967
rect 12808 22924 12860 22933
rect 18052 22924 18104 22976
rect 18972 22924 19024 22976
rect 19248 22967 19300 22976
rect 19248 22933 19257 22967
rect 19257 22933 19291 22967
rect 19291 22933 19300 22967
rect 19248 22924 19300 22933
rect 22468 22924 22520 22976
rect 23204 22924 23256 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 572 22720 624 22772
rect 7380 22720 7432 22772
rect 9680 22720 9732 22772
rect 10048 22720 10100 22772
rect 10324 22763 10376 22772
rect 10324 22729 10333 22763
rect 10333 22729 10367 22763
rect 10367 22729 10376 22763
rect 10324 22720 10376 22729
rect 11888 22763 11940 22772
rect 11888 22729 11897 22763
rect 11897 22729 11931 22763
rect 11931 22729 11940 22763
rect 11888 22720 11940 22729
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 10232 22652 10284 22704
rect 2412 22516 2464 22568
rect 2780 22516 2832 22568
rect 5356 22516 5408 22568
rect 7288 22516 7340 22568
rect 11428 22627 11480 22636
rect 11428 22593 11437 22627
rect 11437 22593 11471 22627
rect 11471 22593 11480 22627
rect 14004 22652 14056 22704
rect 15660 22720 15712 22772
rect 19156 22720 19208 22772
rect 19616 22720 19668 22772
rect 21640 22720 21692 22772
rect 22652 22720 22704 22772
rect 23112 22763 23164 22772
rect 23112 22729 23121 22763
rect 23121 22729 23155 22763
rect 23155 22729 23164 22763
rect 23112 22720 23164 22729
rect 25596 22720 25648 22772
rect 16856 22695 16908 22704
rect 16856 22661 16865 22695
rect 16865 22661 16899 22695
rect 16899 22661 16908 22695
rect 16856 22652 16908 22661
rect 18420 22652 18472 22704
rect 12440 22627 12492 22636
rect 11428 22584 11480 22593
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 17592 22584 17644 22636
rect 18788 22584 18840 22636
rect 18972 22584 19024 22636
rect 19524 22584 19576 22636
rect 10600 22559 10652 22568
rect 10600 22525 10609 22559
rect 10609 22525 10643 22559
rect 10643 22525 10652 22559
rect 10600 22516 10652 22525
rect 10968 22516 11020 22568
rect 12164 22516 12216 22568
rect 1768 22491 1820 22500
rect 1768 22457 1777 22491
rect 1777 22457 1811 22491
rect 1811 22457 1820 22491
rect 1768 22448 1820 22457
rect 11244 22491 11296 22500
rect 11244 22457 11253 22491
rect 11253 22457 11287 22491
rect 11287 22457 11296 22491
rect 11244 22448 11296 22457
rect 12256 22491 12308 22500
rect 12256 22457 12265 22491
rect 12265 22457 12299 22491
rect 12299 22457 12308 22491
rect 13728 22516 13780 22568
rect 15108 22516 15160 22568
rect 16580 22516 16632 22568
rect 19432 22516 19484 22568
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 19800 22516 19852 22525
rect 20076 22559 20128 22568
rect 20076 22525 20099 22559
rect 20099 22525 20128 22559
rect 20076 22516 20128 22525
rect 12256 22448 12308 22457
rect 12992 22448 13044 22500
rect 15752 22491 15804 22500
rect 15752 22457 15786 22491
rect 15786 22457 15804 22491
rect 15752 22448 15804 22457
rect 17408 22448 17460 22500
rect 23480 22559 23532 22568
rect 23480 22525 23489 22559
rect 23489 22525 23523 22559
rect 23523 22525 23532 22559
rect 23480 22516 23532 22525
rect 24860 22516 24912 22568
rect 22560 22491 22612 22500
rect 22560 22457 22569 22491
rect 22569 22457 22603 22491
rect 22603 22457 22612 22491
rect 22560 22448 22612 22457
rect 23572 22448 23624 22500
rect 2964 22380 3016 22432
rect 4252 22380 4304 22432
rect 5540 22380 5592 22432
rect 6644 22423 6696 22432
rect 6644 22389 6653 22423
rect 6653 22389 6687 22423
rect 6687 22389 6696 22423
rect 6644 22380 6696 22389
rect 7472 22380 7524 22432
rect 7840 22380 7892 22432
rect 8760 22423 8812 22432
rect 8760 22389 8769 22423
rect 8769 22389 8803 22423
rect 8803 22389 8812 22423
rect 8760 22380 8812 22389
rect 9128 22380 9180 22432
rect 10784 22423 10836 22432
rect 10784 22389 10793 22423
rect 10793 22389 10827 22423
rect 10827 22389 10836 22423
rect 10784 22380 10836 22389
rect 13912 22380 13964 22432
rect 14004 22380 14056 22432
rect 14280 22380 14332 22432
rect 22100 22423 22152 22432
rect 22100 22389 22109 22423
rect 22109 22389 22143 22423
rect 22143 22389 22152 22423
rect 22100 22380 22152 22389
rect 23388 22380 23440 22432
rect 25596 22516 25648 22568
rect 25228 22380 25280 22432
rect 25780 22423 25832 22432
rect 25780 22389 25789 22423
rect 25789 22389 25823 22423
rect 25823 22389 25832 22423
rect 25780 22380 25832 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2412 22219 2464 22228
rect 2412 22185 2421 22219
rect 2421 22185 2455 22219
rect 2455 22185 2464 22219
rect 2412 22176 2464 22185
rect 3148 22176 3200 22228
rect 4528 22219 4580 22228
rect 4528 22185 4537 22219
rect 4537 22185 4571 22219
rect 4571 22185 4580 22219
rect 4528 22176 4580 22185
rect 6552 22176 6604 22228
rect 6644 22176 6696 22228
rect 1400 22151 1452 22160
rect 1400 22117 1409 22151
rect 1409 22117 1443 22151
rect 1443 22117 1452 22151
rect 1400 22108 1452 22117
rect 2044 22040 2096 22092
rect 4620 22108 4672 22160
rect 7380 22151 7432 22160
rect 7380 22117 7389 22151
rect 7389 22117 7423 22151
rect 7423 22117 7432 22151
rect 7380 22108 7432 22117
rect 4252 22040 4304 22092
rect 6092 22040 6144 22092
rect 8208 22176 8260 22228
rect 10140 22176 10192 22228
rect 11428 22176 11480 22228
rect 12348 22219 12400 22228
rect 12348 22185 12357 22219
rect 12357 22185 12391 22219
rect 12391 22185 12400 22219
rect 12348 22176 12400 22185
rect 8024 22083 8076 22092
rect 8024 22049 8033 22083
rect 8033 22049 8067 22083
rect 8067 22049 8076 22083
rect 8024 22040 8076 22049
rect 11152 22040 11204 22092
rect 12624 22176 12676 22228
rect 15108 22219 15160 22228
rect 15108 22185 15117 22219
rect 15117 22185 15151 22219
rect 15151 22185 15160 22219
rect 15108 22176 15160 22185
rect 15384 22176 15436 22228
rect 16580 22176 16632 22228
rect 17960 22219 18012 22228
rect 17960 22185 17969 22219
rect 17969 22185 18003 22219
rect 18003 22185 18012 22219
rect 17960 22176 18012 22185
rect 20076 22176 20128 22228
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 24124 22219 24176 22228
rect 24124 22185 24133 22219
rect 24133 22185 24167 22219
rect 24167 22185 24176 22219
rect 24124 22176 24176 22185
rect 24584 22176 24636 22228
rect 12532 22108 12584 22160
rect 22376 22151 22428 22160
rect 22376 22117 22410 22151
rect 22410 22117 22428 22151
rect 22376 22108 22428 22117
rect 24216 22108 24268 22160
rect 14004 22040 14056 22092
rect 14832 22040 14884 22092
rect 15200 22040 15252 22092
rect 15292 22040 15344 22092
rect 15660 22083 15712 22092
rect 15660 22049 15669 22083
rect 15669 22049 15703 22083
rect 15703 22049 15712 22083
rect 15660 22040 15712 22049
rect 17132 22040 17184 22092
rect 17868 22040 17920 22092
rect 19064 22040 19116 22092
rect 20996 22083 21048 22092
rect 20996 22049 21005 22083
rect 21005 22049 21039 22083
rect 21039 22049 21048 22083
rect 20996 22040 21048 22049
rect 23388 22040 23440 22092
rect 26056 22040 26108 22092
rect 3056 22015 3108 22024
rect 3056 21981 3065 22015
rect 3065 21981 3099 22015
rect 3099 21981 3108 22015
rect 3056 21972 3108 21981
rect 4436 21904 4488 21956
rect 5172 21972 5224 22024
rect 6460 22015 6512 22024
rect 6460 21981 6469 22015
rect 6469 21981 6503 22015
rect 6503 21981 6512 22015
rect 6460 21972 6512 21981
rect 6828 21972 6880 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 10048 21972 10100 22024
rect 10508 22015 10560 22024
rect 10508 21981 10517 22015
rect 10517 21981 10551 22015
rect 10551 21981 10560 22015
rect 10508 21972 10560 21981
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 12440 21972 12492 22024
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 14188 22015 14240 22024
rect 14188 21981 14197 22015
rect 14197 21981 14231 22015
rect 14231 21981 14240 22015
rect 14188 21972 14240 21981
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 17316 22015 17368 22024
rect 17316 21981 17325 22015
rect 17325 21981 17359 22015
rect 17359 21981 17368 22015
rect 17316 21972 17368 21981
rect 17684 21972 17736 22024
rect 18972 22015 19024 22024
rect 18972 21981 18981 22015
rect 18981 21981 19015 22015
rect 19015 21981 19024 22015
rect 18972 21972 19024 21981
rect 14648 21904 14700 21956
rect 15200 21904 15252 21956
rect 18328 21947 18380 21956
rect 18328 21913 18337 21947
rect 18337 21913 18371 21947
rect 18371 21913 18380 21947
rect 18328 21904 18380 21913
rect 21272 21904 21324 21956
rect 3240 21836 3292 21888
rect 3792 21879 3844 21888
rect 3792 21845 3801 21879
rect 3801 21845 3835 21879
rect 3835 21845 3844 21879
rect 3792 21836 3844 21845
rect 5540 21836 5592 21888
rect 7288 21836 7340 21888
rect 8668 21879 8720 21888
rect 8668 21845 8677 21879
rect 8677 21845 8711 21879
rect 8711 21845 8720 21879
rect 8668 21836 8720 21845
rect 11244 21836 11296 21888
rect 16120 21836 16172 21888
rect 19432 21879 19484 21888
rect 19432 21845 19441 21879
rect 19441 21845 19475 21879
rect 19475 21845 19484 21879
rect 19432 21836 19484 21845
rect 20260 21836 20312 21888
rect 20904 21836 20956 21888
rect 22284 21836 22336 21888
rect 25044 22015 25096 22024
rect 25044 21981 25053 22015
rect 25053 21981 25087 22015
rect 25087 21981 25096 22015
rect 25044 21972 25096 21981
rect 25228 22015 25280 22024
rect 25228 21981 25237 22015
rect 25237 21981 25271 22015
rect 25271 21981 25280 22015
rect 25228 21972 25280 21981
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 25596 21972 25648 21981
rect 23480 21879 23532 21888
rect 23480 21845 23489 21879
rect 23489 21845 23523 21879
rect 23523 21845 23532 21879
rect 23480 21836 23532 21845
rect 23756 21836 23808 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 3056 21632 3108 21684
rect 4528 21632 4580 21684
rect 5356 21675 5408 21684
rect 5356 21641 5365 21675
rect 5365 21641 5399 21675
rect 5399 21641 5408 21675
rect 5356 21632 5408 21641
rect 6828 21632 6880 21684
rect 8116 21632 8168 21684
rect 9128 21675 9180 21684
rect 9128 21641 9137 21675
rect 9137 21641 9171 21675
rect 9171 21641 9180 21675
rect 9128 21632 9180 21641
rect 9588 21632 9640 21684
rect 10140 21675 10192 21684
rect 10140 21641 10149 21675
rect 10149 21641 10183 21675
rect 10183 21641 10192 21675
rect 10140 21632 10192 21641
rect 10508 21675 10560 21684
rect 10508 21641 10517 21675
rect 10517 21641 10551 21675
rect 10551 21641 10560 21675
rect 10508 21632 10560 21641
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12440 21675 12492 21684
rect 12440 21641 12449 21675
rect 12449 21641 12483 21675
rect 12483 21641 12492 21675
rect 14004 21675 14056 21684
rect 12440 21632 12492 21641
rect 14004 21641 14013 21675
rect 14013 21641 14047 21675
rect 14047 21641 14056 21675
rect 14004 21632 14056 21641
rect 14188 21632 14240 21684
rect 14372 21632 14424 21684
rect 14464 21632 14516 21684
rect 14648 21632 14700 21684
rect 15936 21632 15988 21684
rect 16212 21632 16264 21684
rect 18972 21632 19024 21684
rect 19156 21632 19208 21684
rect 22008 21675 22060 21684
rect 22008 21641 22017 21675
rect 22017 21641 22051 21675
rect 22051 21641 22060 21675
rect 22008 21632 22060 21641
rect 25228 21632 25280 21684
rect 2320 21564 2372 21616
rect 12808 21564 12860 21616
rect 17684 21564 17736 21616
rect 18144 21564 18196 21616
rect 22376 21564 22428 21616
rect 3056 21471 3108 21480
rect 3056 21437 3065 21471
rect 3065 21437 3099 21471
rect 3099 21437 3108 21471
rect 3056 21428 3108 21437
rect 7288 21496 7340 21548
rect 11244 21539 11296 21548
rect 11244 21505 11253 21539
rect 11253 21505 11287 21539
rect 11287 21505 11296 21539
rect 11244 21496 11296 21505
rect 11888 21496 11940 21548
rect 12900 21539 12952 21548
rect 12900 21505 12909 21539
rect 12909 21505 12943 21539
rect 12943 21505 12952 21539
rect 12900 21496 12952 21505
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 14004 21496 14056 21548
rect 14648 21496 14700 21548
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 3608 21428 3660 21480
rect 5356 21428 5408 21480
rect 12716 21428 12768 21480
rect 2044 21360 2096 21412
rect 8116 21360 8168 21412
rect 10692 21360 10744 21412
rect 11152 21403 11204 21412
rect 11152 21369 11161 21403
rect 11161 21369 11195 21403
rect 11195 21369 11204 21403
rect 11152 21360 11204 21369
rect 12348 21360 12400 21412
rect 14096 21360 14148 21412
rect 18052 21428 18104 21480
rect 18328 21428 18380 21480
rect 19432 21428 19484 21480
rect 22284 21428 22336 21480
rect 15936 21403 15988 21412
rect 15936 21369 15945 21403
rect 15945 21369 15979 21403
rect 15979 21369 15988 21403
rect 15936 21360 15988 21369
rect 1492 21335 1544 21344
rect 1492 21301 1501 21335
rect 1501 21301 1535 21335
rect 1535 21301 1544 21335
rect 1492 21292 1544 21301
rect 2136 21292 2188 21344
rect 4436 21335 4488 21344
rect 4436 21301 4445 21335
rect 4445 21301 4479 21335
rect 4479 21301 4488 21335
rect 4436 21292 4488 21301
rect 5724 21335 5776 21344
rect 5724 21301 5733 21335
rect 5733 21301 5767 21335
rect 5767 21301 5776 21335
rect 5724 21292 5776 21301
rect 6092 21335 6144 21344
rect 6092 21301 6101 21335
rect 6101 21301 6135 21335
rect 6135 21301 6144 21335
rect 6092 21292 6144 21301
rect 10784 21335 10836 21344
rect 10784 21301 10793 21335
rect 10793 21301 10827 21335
rect 10827 21301 10836 21335
rect 10784 21292 10836 21301
rect 11888 21335 11940 21344
rect 11888 21301 11897 21335
rect 11897 21301 11931 21335
rect 11931 21301 11940 21335
rect 11888 21292 11940 21301
rect 14004 21292 14056 21344
rect 14372 21335 14424 21344
rect 14372 21301 14381 21335
rect 14381 21301 14415 21335
rect 14415 21301 14424 21335
rect 14372 21292 14424 21301
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 15476 21292 15528 21344
rect 18420 21335 18472 21344
rect 18420 21301 18429 21335
rect 18429 21301 18463 21335
rect 18463 21301 18472 21335
rect 18420 21292 18472 21301
rect 19064 21292 19116 21344
rect 20996 21292 21048 21344
rect 21180 21292 21232 21344
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 23756 21428 23808 21480
rect 23480 21403 23532 21412
rect 23480 21369 23489 21403
rect 23489 21369 23523 21403
rect 23523 21369 23532 21403
rect 25228 21428 25280 21480
rect 23480 21360 23532 21369
rect 23756 21292 23808 21344
rect 26056 21292 26108 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1400 21131 1452 21140
rect 1400 21097 1409 21131
rect 1409 21097 1443 21131
rect 1443 21097 1452 21131
rect 1400 21088 1452 21097
rect 2320 21131 2372 21140
rect 2320 21097 2329 21131
rect 2329 21097 2363 21131
rect 2363 21097 2372 21131
rect 2320 21088 2372 21097
rect 3148 21088 3200 21140
rect 4620 21131 4672 21140
rect 4620 21097 4629 21131
rect 4629 21097 4663 21131
rect 4663 21097 4672 21131
rect 4620 21088 4672 21097
rect 3608 21020 3660 21072
rect 6460 21088 6512 21140
rect 7748 21131 7800 21140
rect 7748 21097 7757 21131
rect 7757 21097 7791 21131
rect 7791 21097 7800 21131
rect 7748 21088 7800 21097
rect 7840 21131 7892 21140
rect 7840 21097 7849 21131
rect 7849 21097 7883 21131
rect 7883 21097 7892 21131
rect 7840 21088 7892 21097
rect 8024 21088 8076 21140
rect 11152 21088 11204 21140
rect 11888 21088 11940 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 14096 21131 14148 21140
rect 14096 21097 14105 21131
rect 14105 21097 14139 21131
rect 14139 21097 14148 21131
rect 14096 21088 14148 21097
rect 15292 21088 15344 21140
rect 15660 21088 15712 21140
rect 17040 21131 17092 21140
rect 17040 21097 17049 21131
rect 17049 21097 17083 21131
rect 17083 21097 17092 21131
rect 17040 21088 17092 21097
rect 17132 21088 17184 21140
rect 18604 21088 18656 21140
rect 18972 21088 19024 21140
rect 19340 21088 19392 21140
rect 20720 21131 20772 21140
rect 20720 21097 20729 21131
rect 20729 21097 20763 21131
rect 20763 21097 20772 21131
rect 20720 21088 20772 21097
rect 12992 21020 13044 21072
rect 2688 20952 2740 21004
rect 5172 20995 5224 21004
rect 5172 20961 5206 20995
rect 5206 20961 5224 20995
rect 5172 20952 5224 20961
rect 10692 20952 10744 21004
rect 11152 20952 11204 21004
rect 12808 20952 12860 21004
rect 13728 20952 13780 21004
rect 23388 21088 23440 21140
rect 23112 21020 23164 21072
rect 23664 21088 23716 21140
rect 25044 21088 25096 21140
rect 23756 21063 23808 21072
rect 16488 20952 16540 21004
rect 18420 20952 18472 21004
rect 20168 20952 20220 21004
rect 20720 20952 20772 21004
rect 23756 21029 23790 21063
rect 23790 21029 23808 21063
rect 23756 21020 23808 21029
rect 2596 20884 2648 20936
rect 2780 20816 2832 20868
rect 4436 20884 4488 20936
rect 7932 20927 7984 20936
rect 7932 20893 7941 20927
rect 7941 20893 7975 20927
rect 7975 20893 7984 20927
rect 7932 20884 7984 20893
rect 10140 20884 10192 20936
rect 11980 20884 12032 20936
rect 14280 20884 14332 20936
rect 18696 20927 18748 20936
rect 18696 20893 18705 20927
rect 18705 20893 18739 20927
rect 18739 20893 18748 20927
rect 18696 20884 18748 20893
rect 21088 20884 21140 20936
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 9496 20816 9548 20868
rect 11704 20816 11756 20868
rect 14832 20816 14884 20868
rect 18328 20816 18380 20868
rect 20260 20859 20312 20868
rect 20260 20825 20269 20859
rect 20269 20825 20303 20859
rect 20303 20825 20312 20859
rect 20260 20816 20312 20825
rect 20812 20816 20864 20868
rect 20904 20816 20956 20868
rect 2136 20748 2188 20800
rect 3056 20748 3108 20800
rect 3792 20748 3844 20800
rect 4252 20748 4304 20800
rect 7288 20748 7340 20800
rect 9036 20748 9088 20800
rect 14464 20791 14516 20800
rect 14464 20757 14473 20791
rect 14473 20757 14507 20791
rect 14507 20757 14516 20791
rect 14464 20748 14516 20757
rect 16304 20748 16356 20800
rect 19248 20748 19300 20800
rect 23112 20816 23164 20868
rect 24584 20816 24636 20868
rect 22284 20748 22336 20800
rect 23480 20748 23532 20800
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 2688 20544 2740 20596
rect 7748 20544 7800 20596
rect 7840 20544 7892 20596
rect 10784 20587 10836 20596
rect 10784 20553 10793 20587
rect 10793 20553 10827 20587
rect 10827 20553 10836 20587
rect 10784 20544 10836 20553
rect 11152 20544 11204 20596
rect 14280 20587 14332 20596
rect 4252 20476 4304 20528
rect 11244 20476 11296 20528
rect 14280 20553 14289 20587
rect 14289 20553 14323 20587
rect 14323 20553 14332 20587
rect 14280 20544 14332 20553
rect 14648 20544 14700 20596
rect 15660 20544 15712 20596
rect 16672 20587 16724 20596
rect 16672 20553 16681 20587
rect 16681 20553 16715 20587
rect 16715 20553 16724 20587
rect 16672 20544 16724 20553
rect 18696 20544 18748 20596
rect 19432 20544 19484 20596
rect 23756 20544 23808 20596
rect 12808 20476 12860 20528
rect 17500 20519 17552 20528
rect 17500 20485 17509 20519
rect 17509 20485 17543 20519
rect 17543 20485 17552 20519
rect 17500 20476 17552 20485
rect 3608 20408 3660 20460
rect 5172 20408 5224 20460
rect 5540 20408 5592 20460
rect 7104 20451 7156 20460
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 8116 20451 8168 20460
rect 8116 20417 8125 20451
rect 8125 20417 8159 20451
rect 8159 20417 8168 20451
rect 8116 20408 8168 20417
rect 11428 20451 11480 20460
rect 11428 20417 11437 20451
rect 11437 20417 11471 20451
rect 11471 20417 11480 20451
rect 11428 20408 11480 20417
rect 11888 20408 11940 20460
rect 12716 20408 12768 20460
rect 13912 20408 13964 20460
rect 23572 20408 23624 20460
rect 2320 20272 2372 20324
rect 4804 20383 4856 20392
rect 4804 20349 4813 20383
rect 4813 20349 4847 20383
rect 4847 20349 4856 20383
rect 4804 20340 4856 20349
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 8392 20383 8444 20392
rect 8392 20349 8426 20383
rect 8426 20349 8444 20383
rect 8392 20340 8444 20349
rect 9128 20340 9180 20392
rect 15292 20340 15344 20392
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 2044 20247 2096 20256
rect 2044 20213 2053 20247
rect 2053 20213 2087 20247
rect 2087 20213 2096 20247
rect 2044 20204 2096 20213
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 5540 20247 5592 20256
rect 5540 20213 5549 20247
rect 5549 20213 5583 20247
rect 5583 20213 5592 20247
rect 5540 20204 5592 20213
rect 6000 20204 6052 20256
rect 9404 20204 9456 20256
rect 9772 20204 9824 20256
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 11336 20204 11388 20256
rect 12992 20272 13044 20324
rect 14924 20315 14976 20324
rect 14924 20281 14958 20315
rect 14958 20281 14976 20315
rect 14924 20272 14976 20281
rect 16212 20272 16264 20324
rect 18972 20383 19024 20392
rect 18972 20349 19006 20383
rect 19006 20349 19024 20383
rect 18972 20340 19024 20349
rect 20720 20340 20772 20392
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 12900 20247 12952 20256
rect 12900 20213 12909 20247
rect 12909 20213 12943 20247
rect 12943 20213 12952 20247
rect 12900 20204 12952 20213
rect 13912 20247 13964 20256
rect 13912 20213 13921 20247
rect 13921 20213 13955 20247
rect 13955 20213 13964 20247
rect 13912 20204 13964 20213
rect 17592 20204 17644 20256
rect 18328 20204 18380 20256
rect 20904 20247 20956 20256
rect 20904 20213 20913 20247
rect 20913 20213 20947 20247
rect 20947 20213 20956 20247
rect 20904 20204 20956 20213
rect 20996 20204 21048 20256
rect 21272 20204 21324 20256
rect 22008 20247 22060 20256
rect 22008 20213 22017 20247
rect 22017 20213 22051 20247
rect 22051 20213 22060 20247
rect 22008 20204 22060 20213
rect 22284 20272 22336 20324
rect 23756 20272 23808 20324
rect 25136 20272 25188 20324
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 24124 20247 24176 20256
rect 24124 20213 24133 20247
rect 24133 20213 24167 20247
rect 24167 20213 24176 20247
rect 24124 20204 24176 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 2964 20000 3016 20052
rect 2688 19932 2740 19984
rect 2780 19907 2832 19916
rect 2780 19873 2789 19907
rect 2789 19873 2823 19907
rect 2823 19873 2832 19907
rect 2780 19864 2832 19873
rect 3608 20000 3660 20052
rect 8392 20043 8444 20052
rect 8392 20009 8401 20043
rect 8401 20009 8435 20043
rect 8435 20009 8444 20043
rect 8392 20000 8444 20009
rect 11244 20000 11296 20052
rect 11980 20043 12032 20052
rect 11980 20009 11989 20043
rect 11989 20009 12023 20043
rect 12023 20009 12032 20043
rect 11980 20000 12032 20009
rect 12900 20000 12952 20052
rect 13636 20000 13688 20052
rect 14924 20000 14976 20052
rect 16672 20043 16724 20052
rect 16672 20009 16681 20043
rect 16681 20009 16715 20043
rect 16715 20009 16724 20043
rect 16672 20000 16724 20009
rect 18972 20000 19024 20052
rect 21364 20000 21416 20052
rect 22468 20000 22520 20052
rect 23112 20043 23164 20052
rect 23112 20009 23121 20043
rect 23121 20009 23155 20043
rect 23155 20009 23164 20043
rect 23112 20000 23164 20009
rect 8116 19932 8168 19984
rect 9036 19975 9088 19984
rect 9036 19941 9045 19975
rect 9045 19941 9079 19975
rect 9079 19941 9088 19975
rect 9036 19932 9088 19941
rect 11428 19932 11480 19984
rect 15660 19932 15712 19984
rect 19156 19932 19208 19984
rect 5080 19907 5132 19916
rect 5080 19873 5114 19907
rect 5114 19873 5132 19907
rect 5080 19864 5132 19873
rect 7656 19907 7708 19916
rect 7656 19873 7665 19907
rect 7665 19873 7699 19907
rect 7699 19873 7708 19907
rect 7656 19864 7708 19873
rect 7840 19864 7892 19916
rect 9496 19907 9548 19916
rect 9496 19873 9505 19907
rect 9505 19873 9539 19907
rect 9539 19873 9548 19907
rect 9496 19864 9548 19873
rect 12992 19864 13044 19916
rect 13268 19864 13320 19916
rect 13728 19864 13780 19916
rect 15384 19864 15436 19916
rect 17592 19864 17644 19916
rect 18328 19864 18380 19916
rect 20812 19864 20864 19916
rect 21272 19907 21324 19916
rect 21272 19873 21306 19907
rect 21306 19873 21324 19907
rect 21272 19864 21324 19873
rect 24308 20000 24360 20052
rect 24216 19932 24268 19984
rect 24860 19932 24912 19984
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 2872 19796 2924 19805
rect 3516 19796 3568 19848
rect 4252 19796 4304 19848
rect 7748 19839 7800 19848
rect 7748 19805 7757 19839
rect 7757 19805 7791 19839
rect 7791 19805 7800 19839
rect 7748 19796 7800 19805
rect 7932 19839 7984 19848
rect 7932 19805 7941 19839
rect 7941 19805 7975 19839
rect 7975 19805 7984 19839
rect 7932 19796 7984 19805
rect 9036 19796 9088 19848
rect 2596 19728 2648 19780
rect 3608 19660 3660 19712
rect 4344 19703 4396 19712
rect 4344 19669 4353 19703
rect 4353 19669 4387 19703
rect 4387 19669 4396 19703
rect 4344 19660 4396 19669
rect 4712 19703 4764 19712
rect 4712 19669 4721 19703
rect 4721 19669 4755 19703
rect 4755 19669 4764 19703
rect 4712 19660 4764 19669
rect 5448 19660 5500 19712
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 7196 19660 7248 19712
rect 8576 19660 8628 19712
rect 10140 19796 10192 19848
rect 13268 19728 13320 19780
rect 14556 19728 14608 19780
rect 17868 19728 17920 19780
rect 13084 19703 13136 19712
rect 13084 19669 13093 19703
rect 13093 19669 13127 19703
rect 13127 19669 13136 19703
rect 13084 19660 13136 19669
rect 14464 19660 14516 19712
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 2136 19456 2188 19508
rect 2596 19456 2648 19508
rect 3516 19456 3568 19508
rect 5540 19456 5592 19508
rect 6000 19456 6052 19508
rect 11428 19456 11480 19508
rect 12440 19499 12492 19508
rect 12440 19465 12449 19499
rect 12449 19465 12483 19499
rect 12483 19465 12492 19499
rect 12440 19456 12492 19465
rect 13636 19456 13688 19508
rect 15660 19456 15712 19508
rect 16856 19456 16908 19508
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 19340 19456 19392 19508
rect 23756 19499 23808 19508
rect 2872 19388 2924 19440
rect 3516 19320 3568 19372
rect 7932 19388 7984 19440
rect 10784 19388 10836 19440
rect 12624 19388 12676 19440
rect 15752 19388 15804 19440
rect 23756 19465 23765 19499
rect 23765 19465 23799 19499
rect 23799 19465 23808 19499
rect 23756 19456 23808 19465
rect 25780 19388 25832 19440
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 4252 19295 4304 19304
rect 4252 19261 4261 19295
rect 4261 19261 4295 19295
rect 4295 19261 4304 19295
rect 4252 19252 4304 19261
rect 1676 19227 1728 19236
rect 1676 19193 1685 19227
rect 1685 19193 1719 19227
rect 1719 19193 1728 19227
rect 1676 19184 1728 19193
rect 3884 19184 3936 19236
rect 4160 19227 4212 19236
rect 4160 19193 4169 19227
rect 4169 19193 4203 19227
rect 4203 19193 4212 19227
rect 5080 19252 5132 19304
rect 6828 19320 6880 19372
rect 9220 19363 9272 19372
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 11152 19320 11204 19372
rect 12716 19320 12768 19372
rect 14004 19320 14056 19372
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 16856 19320 16908 19372
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 20812 19363 20864 19372
rect 20812 19329 20821 19363
rect 20821 19329 20855 19363
rect 20855 19329 20864 19363
rect 20812 19320 20864 19329
rect 24308 19363 24360 19372
rect 24308 19329 24317 19363
rect 24317 19329 24351 19363
rect 24351 19329 24360 19363
rect 24308 19320 24360 19329
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 9864 19252 9916 19304
rect 4528 19227 4580 19236
rect 4160 19184 4212 19193
rect 4528 19193 4562 19227
rect 4562 19193 4580 19227
rect 4528 19184 4580 19193
rect 8944 19184 8996 19236
rect 10048 19227 10100 19236
rect 10048 19193 10057 19227
rect 10057 19193 10091 19227
rect 10091 19193 10100 19227
rect 10048 19184 10100 19193
rect 2872 19116 2924 19168
rect 3608 19116 3660 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 8668 19116 8720 19125
rect 9036 19159 9088 19168
rect 9036 19125 9045 19159
rect 9045 19125 9079 19159
rect 9079 19125 9088 19159
rect 9036 19116 9088 19125
rect 11980 19116 12032 19168
rect 13360 19252 13412 19304
rect 16028 19295 16080 19304
rect 14372 19227 14424 19236
rect 14372 19193 14381 19227
rect 14381 19193 14415 19227
rect 14415 19193 14424 19227
rect 14372 19184 14424 19193
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 18420 19295 18472 19304
rect 12440 19116 12492 19168
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 14096 19116 14148 19168
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 14740 19116 14792 19168
rect 17132 19116 17184 19168
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18512 19227 18564 19236
rect 18512 19193 18521 19227
rect 18521 19193 18555 19227
rect 18555 19193 18564 19227
rect 18512 19184 18564 19193
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 19708 19184 19760 19236
rect 21548 19184 21600 19236
rect 22468 19184 22520 19236
rect 25596 19227 25648 19236
rect 25596 19193 25605 19227
rect 25605 19193 25639 19227
rect 25639 19193 25648 19227
rect 25596 19184 25648 19193
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 18052 19116 18104 19125
rect 19524 19159 19576 19168
rect 19524 19125 19533 19159
rect 19533 19125 19567 19159
rect 19567 19125 19576 19159
rect 19524 19116 19576 19125
rect 21272 19116 21324 19168
rect 25780 19116 25832 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 2780 18912 2832 18964
rect 3332 18912 3384 18964
rect 4712 18912 4764 18964
rect 5080 18912 5132 18964
rect 6276 18912 6328 18964
rect 6736 18912 6788 18964
rect 7748 18912 7800 18964
rect 9220 18912 9272 18964
rect 9864 18912 9916 18964
rect 12808 18912 12860 18964
rect 13084 18912 13136 18964
rect 14372 18955 14424 18964
rect 14372 18921 14381 18955
rect 14381 18921 14415 18955
rect 14415 18921 14424 18955
rect 14372 18912 14424 18921
rect 15016 18955 15068 18964
rect 15016 18921 15025 18955
rect 15025 18921 15059 18955
rect 15059 18921 15068 18955
rect 15016 18912 15068 18921
rect 18144 18912 18196 18964
rect 20812 18912 20864 18964
rect 22468 18955 22520 18964
rect 22468 18921 22477 18955
rect 22477 18921 22511 18955
rect 22511 18921 22520 18955
rect 22468 18912 22520 18921
rect 24124 18912 24176 18964
rect 24860 18912 24912 18964
rect 4344 18844 4396 18896
rect 5172 18887 5224 18896
rect 5172 18853 5181 18887
rect 5181 18853 5215 18887
rect 5215 18853 5224 18887
rect 5172 18844 5224 18853
rect 7196 18844 7248 18896
rect 8024 18844 8076 18896
rect 8760 18844 8812 18896
rect 10508 18844 10560 18896
rect 10968 18844 11020 18896
rect 15660 18887 15712 18896
rect 15660 18853 15669 18887
rect 15669 18853 15703 18887
rect 15703 18853 15712 18887
rect 15660 18844 15712 18853
rect 17960 18844 18012 18896
rect 19248 18844 19300 18896
rect 23572 18844 23624 18896
rect 23756 18844 23808 18896
rect 1768 18776 1820 18828
rect 6736 18776 6788 18828
rect 8116 18776 8168 18828
rect 11796 18776 11848 18828
rect 12440 18776 12492 18828
rect 17500 18776 17552 18828
rect 19156 18776 19208 18828
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 20720 18819 20772 18828
rect 20720 18785 20729 18819
rect 20729 18785 20763 18819
rect 20763 18785 20772 18819
rect 20720 18776 20772 18785
rect 21548 18776 21600 18828
rect 24124 18776 24176 18828
rect 25136 18776 25188 18828
rect 1952 18683 2004 18692
rect 1952 18649 1961 18683
rect 1961 18649 1995 18683
rect 1995 18649 2004 18683
rect 1952 18640 2004 18649
rect 4528 18708 4580 18760
rect 5448 18751 5500 18760
rect 5448 18717 5457 18751
rect 5457 18717 5491 18751
rect 5491 18717 5500 18751
rect 5448 18708 5500 18717
rect 4804 18683 4856 18692
rect 4804 18649 4813 18683
rect 4813 18649 4847 18683
rect 4847 18649 4856 18683
rect 4804 18640 4856 18649
rect 6828 18640 6880 18692
rect 2044 18615 2096 18624
rect 2044 18581 2053 18615
rect 2053 18581 2087 18615
rect 2087 18581 2096 18615
rect 2044 18572 2096 18581
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 3884 18615 3936 18624
rect 3884 18581 3893 18615
rect 3893 18581 3927 18615
rect 3927 18581 3936 18615
rect 3884 18572 3936 18581
rect 6552 18572 6604 18624
rect 8300 18708 8352 18760
rect 10416 18751 10468 18760
rect 8668 18640 8720 18692
rect 8300 18572 8352 18624
rect 8576 18572 8628 18624
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 12532 18708 12584 18760
rect 12348 18640 12400 18692
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 9864 18615 9916 18624
rect 9864 18581 9873 18615
rect 9873 18581 9907 18615
rect 9907 18581 9916 18615
rect 9864 18572 9916 18581
rect 11060 18572 11112 18624
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12440 18572 12492 18581
rect 12716 18572 12768 18624
rect 13268 18640 13320 18692
rect 14740 18708 14792 18760
rect 18604 18708 18656 18760
rect 18512 18640 18564 18692
rect 14004 18615 14056 18624
rect 14004 18581 14013 18615
rect 14013 18581 14047 18615
rect 14047 18581 14056 18615
rect 14004 18572 14056 18581
rect 14096 18572 14148 18624
rect 18420 18572 18472 18624
rect 19432 18708 19484 18760
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 23112 18708 23164 18760
rect 23572 18640 23624 18692
rect 24308 18708 24360 18760
rect 18972 18572 19024 18624
rect 19248 18615 19300 18624
rect 19248 18581 19257 18615
rect 19257 18581 19291 18615
rect 19291 18581 19300 18615
rect 19248 18572 19300 18581
rect 21364 18572 21416 18624
rect 23296 18615 23348 18624
rect 23296 18581 23305 18615
rect 23305 18581 23339 18615
rect 23339 18581 23348 18615
rect 23296 18572 23348 18581
rect 23848 18572 23900 18624
rect 24216 18572 24268 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 1768 18411 1820 18420
rect 1768 18377 1777 18411
rect 1777 18377 1811 18411
rect 1811 18377 1820 18411
rect 1768 18368 1820 18377
rect 2504 18368 2556 18420
rect 4160 18368 4212 18420
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 6552 18411 6604 18420
rect 6552 18377 6561 18411
rect 6561 18377 6595 18411
rect 6595 18377 6604 18411
rect 6552 18368 6604 18377
rect 8116 18411 8168 18420
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 9220 18368 9272 18420
rect 10508 18411 10560 18420
rect 10508 18377 10517 18411
rect 10517 18377 10551 18411
rect 10551 18377 10560 18411
rect 10508 18368 10560 18377
rect 12164 18368 12216 18420
rect 12532 18368 12584 18420
rect 10416 18300 10468 18352
rect 11244 18300 11296 18352
rect 11612 18300 11664 18352
rect 15844 18368 15896 18420
rect 16856 18411 16908 18420
rect 16856 18377 16865 18411
rect 16865 18377 16899 18411
rect 16899 18377 16908 18411
rect 16856 18368 16908 18377
rect 17500 18411 17552 18420
rect 17500 18377 17509 18411
rect 17509 18377 17543 18411
rect 17543 18377 17552 18411
rect 17500 18368 17552 18377
rect 18144 18368 18196 18420
rect 4620 18232 4672 18284
rect 5448 18232 5500 18284
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 11888 18275 11940 18284
rect 2136 18164 2188 18216
rect 8576 18164 8628 18216
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 18052 18232 18104 18284
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 12440 18164 12492 18216
rect 12808 18164 12860 18216
rect 15384 18164 15436 18216
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 20720 18368 20772 18420
rect 20996 18411 21048 18420
rect 20996 18377 21005 18411
rect 21005 18377 21039 18411
rect 21039 18377 21048 18411
rect 20996 18368 21048 18377
rect 21456 18368 21508 18420
rect 21824 18368 21876 18420
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 23388 18368 23440 18420
rect 25044 18411 25096 18420
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 25136 18368 25188 18420
rect 25596 18411 25648 18420
rect 25596 18377 25605 18411
rect 25605 18377 25639 18411
rect 25639 18377 25648 18411
rect 25596 18368 25648 18377
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 20996 18164 21048 18216
rect 23296 18164 23348 18216
rect 23756 18164 23808 18216
rect 24768 18164 24820 18216
rect 1952 18096 2004 18148
rect 1768 18028 1820 18080
rect 4068 18028 4120 18080
rect 5724 18096 5776 18148
rect 7656 18096 7708 18148
rect 8668 18096 8720 18148
rect 9128 18096 9180 18148
rect 13728 18096 13780 18148
rect 14740 18096 14792 18148
rect 4988 18071 5040 18080
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 6828 18028 6880 18037
rect 7564 18028 7616 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11428 18071 11480 18080
rect 11428 18037 11437 18071
rect 11437 18037 11471 18071
rect 11471 18037 11480 18071
rect 11428 18028 11480 18037
rect 12532 18028 12584 18080
rect 14096 18028 14148 18080
rect 15108 18028 15160 18080
rect 15844 18028 15896 18080
rect 16488 18028 16540 18080
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 18972 18028 19024 18080
rect 19156 18028 19208 18080
rect 20444 18028 20496 18080
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 22284 18028 22336 18080
rect 23756 18028 23808 18080
rect 24124 18028 24176 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 1400 17824 1452 17876
rect 2044 17824 2096 17876
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 5448 17824 5500 17833
rect 5540 17824 5592 17876
rect 8024 17867 8076 17876
rect 8024 17833 8033 17867
rect 8033 17833 8067 17867
rect 8067 17833 8076 17867
rect 8024 17824 8076 17833
rect 8300 17824 8352 17876
rect 10140 17867 10192 17876
rect 10140 17833 10149 17867
rect 10149 17833 10183 17867
rect 10183 17833 10192 17867
rect 10140 17824 10192 17833
rect 10876 17824 10928 17876
rect 11704 17824 11756 17876
rect 13728 17824 13780 17876
rect 9128 17799 9180 17808
rect 9128 17765 9137 17799
rect 9137 17765 9171 17799
rect 9171 17765 9180 17799
rect 9128 17756 9180 17765
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 2780 17688 2832 17740
rect 4160 17688 4212 17740
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 8392 17731 8444 17740
rect 8392 17697 8401 17731
rect 8401 17697 8435 17731
rect 8435 17697 8444 17731
rect 8392 17688 8444 17697
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 4068 17663 4120 17672
rect 4068 17629 4077 17663
rect 4077 17629 4111 17663
rect 4111 17629 4120 17663
rect 4068 17620 4120 17629
rect 6736 17620 6788 17672
rect 8576 17620 8628 17672
rect 9220 17620 9272 17672
rect 11152 17756 11204 17808
rect 11888 17756 11940 17808
rect 13268 17756 13320 17808
rect 14740 17824 14792 17876
rect 16580 17824 16632 17876
rect 18052 17824 18104 17876
rect 18696 17824 18748 17876
rect 21548 17824 21600 17876
rect 22652 17867 22704 17876
rect 22652 17833 22661 17867
rect 22661 17833 22695 17867
rect 22695 17833 22704 17867
rect 22652 17824 22704 17833
rect 23572 17867 23624 17876
rect 23572 17833 23581 17867
rect 23581 17833 23615 17867
rect 23615 17833 23624 17867
rect 23572 17824 23624 17833
rect 24860 17824 24912 17876
rect 15200 17756 15252 17808
rect 15936 17756 15988 17808
rect 17868 17756 17920 17808
rect 18512 17756 18564 17808
rect 19524 17756 19576 17808
rect 21364 17799 21416 17808
rect 21364 17765 21373 17799
rect 21373 17765 21407 17799
rect 21407 17765 21416 17799
rect 21364 17756 21416 17765
rect 23848 17756 23900 17808
rect 9956 17688 10008 17740
rect 11244 17731 11296 17740
rect 11244 17697 11253 17731
rect 11253 17697 11287 17731
rect 11287 17697 11296 17731
rect 11244 17688 11296 17697
rect 12348 17688 12400 17740
rect 14556 17688 14608 17740
rect 15108 17688 15160 17740
rect 15384 17688 15436 17740
rect 17040 17688 17092 17740
rect 18052 17688 18104 17740
rect 19432 17688 19484 17740
rect 10968 17620 11020 17672
rect 18328 17663 18380 17672
rect 18328 17629 18337 17663
rect 18337 17629 18371 17663
rect 18371 17629 18380 17663
rect 18328 17620 18380 17629
rect 7656 17552 7708 17604
rect 8392 17552 8444 17604
rect 13820 17552 13872 17604
rect 14556 17552 14608 17604
rect 14924 17595 14976 17604
rect 14924 17561 14933 17595
rect 14933 17561 14967 17595
rect 14967 17561 14976 17595
rect 14924 17552 14976 17561
rect 17776 17595 17828 17604
rect 17776 17561 17785 17595
rect 17785 17561 17819 17595
rect 17819 17561 17828 17595
rect 17776 17552 17828 17561
rect 21088 17688 21140 17740
rect 22928 17688 22980 17740
rect 20996 17620 21048 17672
rect 23480 17620 23532 17672
rect 2964 17527 3016 17536
rect 2964 17493 2973 17527
rect 2973 17493 3007 17527
rect 3007 17493 3016 17527
rect 2964 17484 3016 17493
rect 3516 17484 3568 17536
rect 6736 17484 6788 17536
rect 7380 17484 7432 17536
rect 7564 17527 7616 17536
rect 7564 17493 7573 17527
rect 7573 17493 7607 17527
rect 7607 17493 7616 17527
rect 7564 17484 7616 17493
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 9220 17484 9272 17536
rect 9496 17484 9548 17536
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 20536 17484 20588 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2412 17280 2464 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 5080 17323 5132 17332
rect 5080 17289 5089 17323
rect 5089 17289 5123 17323
rect 5123 17289 5132 17323
rect 5080 17280 5132 17289
rect 6092 17323 6144 17332
rect 6092 17289 6101 17323
rect 6101 17289 6135 17323
rect 6135 17289 6144 17323
rect 6092 17280 6144 17289
rect 6184 17280 6236 17332
rect 5448 17144 5500 17196
rect 2136 17119 2188 17128
rect 2136 17085 2145 17119
rect 2145 17085 2179 17119
rect 2179 17085 2188 17119
rect 2136 17076 2188 17085
rect 4068 17076 4120 17128
rect 4896 17076 4948 17128
rect 9496 17280 9548 17332
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 10140 17280 10192 17332
rect 11152 17280 11204 17332
rect 13176 17280 13228 17332
rect 13820 17280 13872 17332
rect 15936 17323 15988 17332
rect 15936 17289 15945 17323
rect 15945 17289 15979 17323
rect 15979 17289 15988 17323
rect 15936 17280 15988 17289
rect 18328 17280 18380 17332
rect 21088 17280 21140 17332
rect 21364 17280 21416 17332
rect 23848 17280 23900 17332
rect 7012 17255 7064 17264
rect 7012 17221 7021 17255
rect 7021 17221 7055 17255
rect 7055 17221 7064 17255
rect 7012 17212 7064 17221
rect 14648 17212 14700 17264
rect 21824 17255 21876 17264
rect 10876 17144 10928 17196
rect 11060 17144 11112 17196
rect 12348 17144 12400 17196
rect 8576 17119 8628 17128
rect 8576 17085 8610 17119
rect 8610 17085 8628 17119
rect 2504 17008 2556 17060
rect 8116 17008 8168 17060
rect 8576 17076 8628 17085
rect 9680 17076 9732 17128
rect 10784 17076 10836 17128
rect 21824 17221 21833 17255
rect 21833 17221 21867 17255
rect 21867 17221 21876 17255
rect 21824 17212 21876 17221
rect 14832 17144 14884 17196
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 9864 17008 9916 17060
rect 10876 17008 10928 17060
rect 11428 17008 11480 17060
rect 12624 17008 12676 17060
rect 14924 17008 14976 17060
rect 20444 17119 20496 17128
rect 20444 17085 20453 17119
rect 20453 17085 20487 17119
rect 20487 17085 20496 17119
rect 20444 17076 20496 17085
rect 24308 17187 24360 17196
rect 24308 17153 24317 17187
rect 24317 17153 24351 17187
rect 24351 17153 24360 17187
rect 24308 17144 24360 17153
rect 17132 17008 17184 17060
rect 18236 17008 18288 17060
rect 20536 17008 20588 17060
rect 23756 17008 23808 17060
rect 25136 17008 25188 17060
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 5172 16940 5224 16992
rect 10140 16940 10192 16992
rect 10968 16940 11020 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 11888 16983 11940 16992
rect 11888 16949 11897 16983
rect 11897 16949 11931 16983
rect 11931 16949 11940 16983
rect 11888 16940 11940 16949
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 16304 16983 16356 16992
rect 16304 16949 16313 16983
rect 16313 16949 16347 16983
rect 16347 16949 16356 16983
rect 16304 16940 16356 16949
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 18512 16983 18564 16992
rect 18512 16949 18521 16983
rect 18521 16949 18555 16983
rect 18555 16949 18564 16983
rect 18512 16940 18564 16949
rect 20904 16940 20956 16992
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2228 16736 2280 16788
rect 2044 16668 2096 16720
rect 2504 16668 2556 16720
rect 2964 16736 3016 16788
rect 3516 16736 3568 16788
rect 4528 16736 4580 16788
rect 5172 16779 5224 16788
rect 5172 16745 5181 16779
rect 5181 16745 5215 16779
rect 5215 16745 5224 16779
rect 5172 16736 5224 16745
rect 6736 16779 6788 16788
rect 6736 16745 6745 16779
rect 6745 16745 6779 16779
rect 6779 16745 6788 16779
rect 6736 16736 6788 16745
rect 6920 16736 6972 16788
rect 8300 16736 8352 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 10140 16779 10192 16788
rect 10140 16745 10149 16779
rect 10149 16745 10183 16779
rect 10183 16745 10192 16779
rect 10140 16736 10192 16745
rect 10876 16779 10928 16788
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 14924 16779 14976 16788
rect 14924 16745 14933 16779
rect 14933 16745 14967 16779
rect 14967 16745 14976 16779
rect 14924 16736 14976 16745
rect 16304 16736 16356 16788
rect 18052 16736 18104 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 19984 16736 20036 16788
rect 20904 16736 20956 16788
rect 22928 16779 22980 16788
rect 22928 16745 22937 16779
rect 22937 16745 22971 16779
rect 22971 16745 22980 16779
rect 22928 16736 22980 16745
rect 23296 16779 23348 16788
rect 23296 16745 23305 16779
rect 23305 16745 23339 16779
rect 23339 16745 23348 16779
rect 23296 16736 23348 16745
rect 24308 16736 24360 16788
rect 1860 16600 1912 16652
rect 1952 16600 2004 16652
rect 2872 16668 2924 16720
rect 6552 16668 6604 16720
rect 8576 16668 8628 16720
rect 9956 16668 10008 16720
rect 10692 16668 10744 16720
rect 14832 16668 14884 16720
rect 15476 16668 15528 16720
rect 17500 16668 17552 16720
rect 20720 16668 20772 16720
rect 21824 16668 21876 16720
rect 3516 16532 3568 16584
rect 6184 16600 6236 16652
rect 4436 16532 4488 16584
rect 5356 16575 5408 16584
rect 5356 16541 5365 16575
rect 5365 16541 5399 16575
rect 5399 16541 5408 16575
rect 5356 16532 5408 16541
rect 7748 16532 7800 16584
rect 9312 16600 9364 16652
rect 10508 16600 10560 16652
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 11796 16600 11848 16652
rect 12624 16600 12676 16652
rect 12808 16600 12860 16652
rect 7932 16507 7984 16516
rect 7932 16473 7941 16507
rect 7941 16473 7975 16507
rect 7975 16473 7984 16507
rect 9588 16532 9640 16584
rect 10232 16575 10284 16584
rect 10232 16541 10241 16575
rect 10241 16541 10275 16575
rect 10275 16541 10284 16575
rect 10232 16532 10284 16541
rect 14004 16600 14056 16652
rect 14372 16600 14424 16652
rect 17040 16643 17092 16652
rect 17040 16609 17049 16643
rect 17049 16609 17083 16643
rect 17083 16609 17092 16643
rect 17040 16600 17092 16609
rect 19340 16600 19392 16652
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 20444 16532 20496 16584
rect 20812 16532 20864 16584
rect 23296 16532 23348 16584
rect 23480 16600 23532 16652
rect 24032 16643 24084 16652
rect 24032 16609 24066 16643
rect 24066 16609 24084 16643
rect 24032 16600 24084 16609
rect 7932 16464 7984 16473
rect 14188 16464 14240 16516
rect 18696 16464 18748 16516
rect 14464 16396 14516 16448
rect 16580 16396 16632 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2504 16235 2556 16244
rect 2504 16201 2513 16235
rect 2513 16201 2547 16235
rect 2547 16201 2556 16235
rect 2504 16192 2556 16201
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 6276 16235 6328 16244
rect 2780 16192 2832 16201
rect 6276 16201 6285 16235
rect 6285 16201 6319 16235
rect 6319 16201 6328 16235
rect 6276 16192 6328 16201
rect 6644 16235 6696 16244
rect 6644 16201 6653 16235
rect 6653 16201 6687 16235
rect 6687 16201 6696 16235
rect 6644 16192 6696 16201
rect 8208 16192 8260 16244
rect 9588 16235 9640 16244
rect 9588 16201 9597 16235
rect 9597 16201 9631 16235
rect 9631 16201 9640 16235
rect 9588 16192 9640 16201
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 10508 16235 10560 16244
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 11796 16235 11848 16244
rect 11796 16201 11805 16235
rect 11805 16201 11839 16235
rect 11839 16201 11848 16235
rect 11796 16192 11848 16201
rect 7748 16167 7800 16176
rect 7748 16133 7757 16167
rect 7757 16133 7791 16167
rect 7791 16133 7800 16167
rect 7748 16124 7800 16133
rect 8024 16167 8076 16176
rect 8024 16133 8033 16167
rect 8033 16133 8067 16167
rect 8067 16133 8076 16167
rect 8024 16124 8076 16133
rect 12440 16192 12492 16244
rect 12992 16192 13044 16244
rect 14372 16192 14424 16244
rect 15844 16192 15896 16244
rect 16488 16192 16540 16244
rect 18328 16192 18380 16244
rect 20720 16192 20772 16244
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 23756 16235 23808 16244
rect 23756 16201 23765 16235
rect 23765 16201 23799 16235
rect 23799 16201 23808 16235
rect 23756 16192 23808 16201
rect 25504 16235 25556 16244
rect 25504 16201 25513 16235
rect 25513 16201 25547 16235
rect 25547 16201 25556 16235
rect 25504 16192 25556 16201
rect 19340 16124 19392 16176
rect 3240 16099 3292 16108
rect 3240 16065 3249 16099
rect 3249 16065 3283 16099
rect 3283 16065 3292 16099
rect 3240 16056 3292 16065
rect 3516 16056 3568 16108
rect 1860 15988 1912 16040
rect 1676 15963 1728 15972
rect 1676 15929 1685 15963
rect 1685 15929 1719 15963
rect 1719 15929 1728 15963
rect 1676 15920 1728 15929
rect 2228 15963 2280 15972
rect 2228 15929 2237 15963
rect 2237 15929 2271 15963
rect 2271 15929 2280 15963
rect 2872 15988 2924 16040
rect 2228 15920 2280 15929
rect 6092 16056 6144 16108
rect 7472 16056 7524 16108
rect 8116 16056 8168 16108
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 12808 16056 12860 16108
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 4988 15988 5040 16040
rect 9496 15988 9548 16040
rect 6828 15920 6880 15972
rect 10784 15920 10836 15972
rect 4988 15895 5040 15904
rect 4988 15861 4997 15895
rect 4997 15861 5031 15895
rect 5031 15861 5040 15895
rect 4988 15852 5040 15861
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 12256 15852 12308 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13636 15852 13688 15904
rect 14096 16056 14148 16108
rect 17500 16056 17552 16108
rect 16580 15988 16632 16040
rect 17408 15988 17460 16040
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 18696 15988 18748 16040
rect 20720 15988 20772 16040
rect 22468 16056 22520 16108
rect 22836 16056 22888 16108
rect 24032 16056 24084 16108
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 25228 15988 25280 16040
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 22836 15920 22888 15972
rect 14188 15852 14240 15904
rect 14464 15895 14516 15904
rect 14464 15861 14473 15895
rect 14473 15861 14507 15895
rect 14507 15861 14516 15895
rect 17500 15895 17552 15904
rect 14464 15852 14516 15861
rect 17500 15861 17509 15895
rect 17509 15861 17543 15895
rect 17543 15861 17552 15895
rect 17500 15852 17552 15861
rect 22928 15852 22980 15904
rect 23480 15895 23532 15904
rect 23480 15861 23489 15895
rect 23489 15861 23523 15895
rect 23523 15861 23532 15895
rect 23480 15852 23532 15861
rect 25504 15852 25556 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 3240 15648 3292 15700
rect 3976 15648 4028 15700
rect 4436 15648 4488 15700
rect 5448 15648 5500 15700
rect 6736 15648 6788 15700
rect 9496 15648 9548 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10140 15648 10192 15700
rect 10784 15691 10836 15700
rect 10784 15657 10793 15691
rect 10793 15657 10827 15691
rect 10827 15657 10836 15691
rect 10784 15648 10836 15657
rect 12900 15691 12952 15700
rect 12900 15657 12909 15691
rect 12909 15657 12943 15691
rect 12943 15657 12952 15691
rect 12900 15648 12952 15657
rect 14004 15648 14056 15700
rect 18236 15691 18288 15700
rect 18236 15657 18245 15691
rect 18245 15657 18279 15691
rect 18279 15657 18288 15691
rect 18236 15648 18288 15657
rect 21088 15648 21140 15700
rect 22284 15691 22336 15700
rect 22284 15657 22293 15691
rect 22293 15657 22327 15691
rect 22327 15657 22336 15691
rect 22284 15648 22336 15657
rect 24768 15691 24820 15700
rect 24768 15657 24777 15691
rect 24777 15657 24811 15691
rect 24811 15657 24820 15691
rect 24768 15648 24820 15657
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 3976 15512 4028 15564
rect 6552 15580 6604 15632
rect 7932 15580 7984 15632
rect 11060 15580 11112 15632
rect 18328 15580 18380 15632
rect 22928 15580 22980 15632
rect 24032 15580 24084 15632
rect 5540 15512 5592 15564
rect 8116 15512 8168 15564
rect 9496 15555 9548 15564
rect 9496 15521 9505 15555
rect 9505 15521 9539 15555
rect 9539 15521 9548 15555
rect 9496 15512 9548 15521
rect 13728 15555 13780 15564
rect 13728 15521 13737 15555
rect 13737 15521 13771 15555
rect 13771 15521 13780 15555
rect 13728 15512 13780 15521
rect 16304 15512 16356 15564
rect 17960 15512 18012 15564
rect 20904 15512 20956 15564
rect 22652 15555 22704 15564
rect 22652 15521 22661 15555
rect 22661 15521 22695 15555
rect 22695 15521 22704 15555
rect 22652 15512 22704 15521
rect 2412 15487 2464 15496
rect 2412 15453 2421 15487
rect 2421 15453 2455 15487
rect 2455 15453 2464 15487
rect 2412 15444 2464 15453
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 6092 15487 6144 15496
rect 2504 15444 2556 15453
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 9680 15444 9732 15496
rect 13820 15487 13872 15496
rect 13820 15453 13829 15487
rect 13829 15453 13863 15487
rect 13863 15453 13872 15487
rect 13820 15444 13872 15453
rect 13912 15487 13964 15496
rect 13912 15453 13921 15487
rect 13921 15453 13955 15487
rect 13955 15453 13964 15487
rect 13912 15444 13964 15453
rect 18696 15487 18748 15496
rect 1952 15376 2004 15428
rect 7012 15376 7064 15428
rect 13084 15376 13136 15428
rect 2044 15308 2096 15360
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 3700 15308 3752 15360
rect 4160 15308 4212 15360
rect 5356 15308 5408 15360
rect 7288 15308 7340 15360
rect 8300 15308 8352 15360
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 13176 15308 13228 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 17500 15376 17552 15428
rect 18972 15444 19024 15496
rect 20352 15444 20404 15496
rect 21364 15487 21416 15496
rect 21364 15453 21373 15487
rect 21373 15453 21407 15487
rect 21407 15453 21416 15487
rect 21364 15444 21416 15453
rect 21824 15444 21876 15496
rect 16120 15308 16172 15360
rect 16488 15308 16540 15360
rect 17592 15308 17644 15360
rect 17776 15308 17828 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 20720 15308 20772 15360
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 1952 15036 2004 15088
rect 2412 15036 2464 15088
rect 4344 15104 4396 15156
rect 5080 15104 5132 15156
rect 5264 15104 5316 15156
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 8116 15104 8168 15156
rect 4252 15036 4304 15088
rect 6276 15036 6328 15088
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 6092 14968 6144 15020
rect 7564 14968 7616 15020
rect 8208 14968 8260 15020
rect 8484 14968 8536 15020
rect 3056 14900 3108 14952
rect 6644 14943 6696 14952
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 2780 14832 2832 14884
rect 3240 14832 3292 14884
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 7196 14943 7248 14952
rect 6644 14900 6696 14909
rect 7196 14909 7205 14943
rect 7205 14909 7239 14943
rect 7239 14909 7248 14943
rect 7196 14900 7248 14909
rect 8760 14900 8812 14952
rect 11060 15104 11112 15156
rect 12808 15104 12860 15156
rect 13728 15104 13780 15156
rect 14648 15104 14700 15156
rect 17868 15147 17920 15156
rect 13176 15036 13228 15088
rect 17868 15113 17877 15147
rect 17877 15113 17911 15147
rect 17911 15113 17920 15147
rect 17868 15104 17920 15113
rect 20352 15147 20404 15156
rect 20352 15113 20361 15147
rect 20361 15113 20395 15147
rect 20395 15113 20404 15147
rect 20352 15104 20404 15113
rect 20904 15147 20956 15156
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 21824 15104 21876 15156
rect 22100 15104 22152 15156
rect 9588 14943 9640 14952
rect 9588 14909 9597 14943
rect 9597 14909 9631 14943
rect 9631 14909 9640 14943
rect 9588 14900 9640 14909
rect 13912 14968 13964 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 17316 15036 17368 15088
rect 15660 14968 15712 14977
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 20536 14968 20588 15020
rect 22100 14968 22152 15020
rect 10140 14900 10192 14952
rect 12532 14900 12584 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 15936 14900 15988 14952
rect 16488 14900 16540 14952
rect 16764 14943 16816 14952
rect 16764 14909 16773 14943
rect 16773 14909 16807 14943
rect 16807 14909 16816 14943
rect 16764 14900 16816 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 18328 14943 18380 14952
rect 18328 14909 18362 14943
rect 18362 14909 18380 14943
rect 18328 14900 18380 14909
rect 20352 14900 20404 14952
rect 11980 14832 12032 14884
rect 15292 14832 15344 14884
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 6920 14764 6972 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 12808 14807 12860 14816
rect 12808 14773 12817 14807
rect 12817 14773 12851 14807
rect 12851 14773 12860 14807
rect 12808 14764 12860 14773
rect 14096 14764 14148 14816
rect 16120 14807 16172 14816
rect 16120 14773 16129 14807
rect 16129 14773 16163 14807
rect 16163 14773 16172 14807
rect 16120 14764 16172 14773
rect 16672 14764 16724 14816
rect 16948 14764 17000 14816
rect 17960 14832 18012 14884
rect 22744 15104 22796 15156
rect 22928 15104 22980 15156
rect 24124 15104 24176 15156
rect 24768 15147 24820 15156
rect 24768 15113 24777 15147
rect 24777 15113 24811 15147
rect 24811 15113 24820 15147
rect 24768 15104 24820 15113
rect 25412 15104 25464 15156
rect 23204 15036 23256 15088
rect 25688 14900 25740 14952
rect 22744 14832 22796 14884
rect 24216 14875 24268 14884
rect 24216 14841 24225 14875
rect 24225 14841 24259 14875
rect 24259 14841 24268 14875
rect 24216 14832 24268 14841
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 20996 14764 21048 14816
rect 24768 14764 24820 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 5172 14560 5224 14612
rect 5448 14560 5500 14612
rect 4620 14535 4672 14544
rect 4620 14501 4629 14535
rect 4629 14501 4663 14535
rect 4663 14501 4672 14535
rect 4620 14492 4672 14501
rect 6092 14560 6144 14612
rect 7104 14560 7156 14612
rect 8760 14603 8812 14612
rect 8760 14569 8769 14603
rect 8769 14569 8803 14603
rect 8803 14569 8812 14603
rect 8760 14560 8812 14569
rect 11060 14560 11112 14612
rect 12256 14560 12308 14612
rect 13176 14560 13228 14612
rect 18972 14560 19024 14612
rect 21916 14560 21968 14612
rect 22100 14560 22152 14612
rect 22652 14560 22704 14612
rect 23020 14560 23072 14612
rect 24216 14560 24268 14612
rect 7564 14492 7616 14544
rect 10140 14535 10192 14544
rect 10140 14501 10149 14535
rect 10149 14501 10183 14535
rect 10183 14501 10192 14535
rect 10140 14492 10192 14501
rect 12348 14492 12400 14544
rect 12624 14492 12676 14544
rect 13268 14492 13320 14544
rect 14096 14535 14148 14544
rect 14096 14501 14105 14535
rect 14105 14501 14139 14535
rect 14139 14501 14148 14535
rect 14096 14492 14148 14501
rect 1768 14467 1820 14476
rect 1768 14433 1802 14467
rect 1802 14433 1820 14467
rect 1768 14424 1820 14433
rect 1492 14399 1544 14408
rect 1492 14365 1501 14399
rect 1501 14365 1535 14399
rect 1535 14365 1544 14399
rect 1492 14356 1544 14365
rect 4712 14399 4764 14408
rect 4712 14365 4721 14399
rect 4721 14365 4755 14399
rect 4755 14365 4764 14399
rect 4712 14356 4764 14365
rect 5448 14356 5500 14408
rect 8208 14424 8260 14476
rect 12440 14424 12492 14476
rect 13360 14424 13412 14476
rect 15844 14424 15896 14476
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 13084 14356 13136 14408
rect 13820 14356 13872 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 20168 14492 20220 14544
rect 21364 14492 21416 14544
rect 18420 14356 18472 14365
rect 20260 14424 20312 14476
rect 22284 14424 22336 14476
rect 20720 14356 20772 14408
rect 22100 14356 22152 14408
rect 23848 14492 23900 14544
rect 23572 14424 23624 14476
rect 25044 14424 25096 14476
rect 23480 14356 23532 14408
rect 24032 14399 24084 14408
rect 24032 14365 24041 14399
rect 24041 14365 24075 14399
rect 24075 14365 24084 14399
rect 24032 14356 24084 14365
rect 25228 14399 25280 14408
rect 25228 14365 25237 14399
rect 25237 14365 25271 14399
rect 25271 14365 25280 14399
rect 25228 14356 25280 14365
rect 2780 14220 2832 14272
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 7104 14263 7156 14272
rect 7104 14229 7113 14263
rect 7113 14229 7147 14263
rect 7147 14229 7156 14263
rect 7104 14220 7156 14229
rect 11336 14220 11388 14272
rect 12808 14220 12860 14272
rect 13176 14220 13228 14272
rect 13268 14220 13320 14272
rect 13728 14220 13780 14272
rect 13912 14220 13964 14272
rect 15476 14220 15528 14272
rect 17040 14288 17092 14340
rect 19340 14288 19392 14340
rect 23204 14288 23256 14340
rect 16304 14220 16356 14272
rect 18788 14220 18840 14272
rect 19248 14220 19300 14272
rect 23296 14263 23348 14272
rect 23296 14229 23305 14263
rect 23305 14229 23339 14263
rect 23339 14229 23348 14263
rect 23296 14220 23348 14229
rect 26332 14220 26384 14272
rect 27068 14220 27120 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2320 14016 2372 14068
rect 3056 14016 3108 14068
rect 3792 14016 3844 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 6000 14016 6052 14068
rect 7104 14016 7156 14068
rect 8208 14059 8260 14068
rect 8208 14025 8217 14059
rect 8217 14025 8251 14059
rect 8251 14025 8260 14059
rect 8208 14016 8260 14025
rect 10048 14016 10100 14068
rect 12440 14059 12492 14068
rect 12440 14025 12449 14059
rect 12449 14025 12483 14059
rect 12483 14025 12492 14059
rect 12440 14016 12492 14025
rect 12992 14016 13044 14068
rect 13452 14016 13504 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 14280 14016 14332 14068
rect 14556 14016 14608 14068
rect 15844 14059 15896 14068
rect 2596 13991 2648 14000
rect 2596 13957 2605 13991
rect 2605 13957 2639 13991
rect 2639 13957 2648 13991
rect 2596 13948 2648 13957
rect 3976 13948 4028 14000
rect 2596 13812 2648 13864
rect 1492 13744 1544 13796
rect 1952 13744 2004 13796
rect 6736 13880 6788 13932
rect 7012 13880 7064 13932
rect 12900 13948 12952 14000
rect 2964 13855 3016 13864
rect 2964 13821 2998 13855
rect 2998 13821 3016 13855
rect 2964 13812 3016 13821
rect 4160 13812 4212 13864
rect 3240 13744 3292 13796
rect 3056 13676 3108 13728
rect 5540 13676 5592 13728
rect 6092 13812 6144 13864
rect 7104 13812 7156 13864
rect 13544 13880 13596 13932
rect 6920 13744 6972 13796
rect 8760 13744 8812 13796
rect 9588 13812 9640 13864
rect 12348 13812 12400 13864
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 12072 13744 12124 13796
rect 13084 13744 13136 13796
rect 15844 14025 15853 14059
rect 15853 14025 15887 14059
rect 15887 14025 15896 14059
rect 15844 14016 15896 14025
rect 18236 14059 18288 14068
rect 18236 14025 18245 14059
rect 18245 14025 18279 14059
rect 18279 14025 18288 14059
rect 18236 14016 18288 14025
rect 20260 14016 20312 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21364 14016 21416 14068
rect 22284 14059 22336 14068
rect 22284 14025 22293 14059
rect 22293 14025 22327 14059
rect 22327 14025 22336 14059
rect 22284 14016 22336 14025
rect 16028 13948 16080 14000
rect 16488 13948 16540 14000
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 16672 13880 16724 13932
rect 18420 13948 18472 14000
rect 22928 13948 22980 14000
rect 23664 13948 23716 14000
rect 24584 13948 24636 14000
rect 17960 13812 18012 13864
rect 18788 13855 18840 13864
rect 18788 13821 18797 13855
rect 18797 13821 18831 13855
rect 18831 13821 18840 13855
rect 18788 13812 18840 13821
rect 21916 13923 21968 13932
rect 19064 13855 19116 13864
rect 19064 13821 19087 13855
rect 19087 13821 19116 13855
rect 21916 13889 21925 13923
rect 21925 13889 21959 13923
rect 21959 13889 21968 13923
rect 21916 13880 21968 13889
rect 22744 13880 22796 13932
rect 23020 13880 23072 13932
rect 23480 13880 23532 13932
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25412 13923 25464 13932
rect 25412 13889 25421 13923
rect 25421 13889 25455 13923
rect 25455 13889 25464 13923
rect 25412 13880 25464 13889
rect 19064 13812 19116 13821
rect 21824 13812 21876 13864
rect 23572 13812 23624 13864
rect 23756 13812 23808 13864
rect 23848 13812 23900 13864
rect 24952 13812 25004 13864
rect 17224 13744 17276 13796
rect 24676 13744 24728 13796
rect 11796 13676 11848 13728
rect 12532 13676 12584 13728
rect 13544 13719 13596 13728
rect 13544 13685 13553 13719
rect 13553 13685 13587 13719
rect 13587 13685 13596 13719
rect 13544 13676 13596 13685
rect 14740 13676 14792 13728
rect 21640 13719 21692 13728
rect 21640 13685 21649 13719
rect 21649 13685 21683 13719
rect 21683 13685 21692 13719
rect 21640 13676 21692 13685
rect 23480 13676 23532 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 1860 13472 1912 13524
rect 3240 13472 3292 13524
rect 3976 13472 4028 13524
rect 4068 13472 4120 13524
rect 4620 13515 4672 13524
rect 4620 13481 4629 13515
rect 4629 13481 4663 13515
rect 4663 13481 4672 13515
rect 4620 13472 4672 13481
rect 6920 13472 6972 13524
rect 7656 13472 7708 13524
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 8576 13472 8628 13524
rect 8760 13472 8812 13524
rect 9772 13515 9824 13524
rect 2596 13404 2648 13456
rect 2228 13336 2280 13388
rect 2688 13336 2740 13388
rect 6000 13404 6052 13456
rect 8668 13404 8720 13456
rect 4620 13336 4672 13388
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 14740 13472 14792 13524
rect 16580 13472 16632 13524
rect 17224 13515 17276 13524
rect 17224 13481 17233 13515
rect 17233 13481 17267 13515
rect 17267 13481 17276 13515
rect 17224 13472 17276 13481
rect 19340 13472 19392 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 21916 13515 21968 13524
rect 21916 13481 21925 13515
rect 21925 13481 21959 13515
rect 21959 13481 21968 13515
rect 21916 13472 21968 13481
rect 22192 13472 22244 13524
rect 23204 13472 23256 13524
rect 24216 13472 24268 13524
rect 15476 13404 15528 13456
rect 17040 13404 17092 13456
rect 17776 13404 17828 13456
rect 22744 13404 22796 13456
rect 23112 13404 23164 13456
rect 10140 13336 10192 13388
rect 10324 13336 10376 13388
rect 11796 13336 11848 13388
rect 12164 13336 12216 13388
rect 14280 13336 14332 13388
rect 15292 13379 15344 13388
rect 15292 13345 15301 13379
rect 15301 13345 15335 13379
rect 15335 13345 15344 13379
rect 15292 13336 15344 13345
rect 16120 13336 16172 13388
rect 21272 13379 21324 13388
rect 21272 13345 21281 13379
rect 21281 13345 21315 13379
rect 21315 13345 21324 13379
rect 21272 13336 21324 13345
rect 22468 13379 22520 13388
rect 22468 13345 22477 13379
rect 22477 13345 22511 13379
rect 22511 13345 22520 13379
rect 22468 13336 22520 13345
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 3792 13268 3844 13320
rect 5448 13268 5500 13320
rect 8484 13268 8536 13320
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 20812 13268 20864 13320
rect 21364 13268 21416 13320
rect 4068 13200 4120 13252
rect 6736 13200 6788 13252
rect 12256 13200 12308 13252
rect 1768 13132 1820 13184
rect 3056 13132 3108 13184
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 11612 13175 11664 13184
rect 11612 13141 11621 13175
rect 11621 13141 11655 13175
rect 11655 13141 11664 13175
rect 11612 13132 11664 13141
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 19064 13200 19116 13252
rect 25320 13336 25372 13388
rect 23296 13268 23348 13320
rect 15936 13132 15988 13184
rect 17868 13175 17920 13184
rect 17868 13141 17877 13175
rect 17877 13141 17911 13175
rect 17911 13141 17920 13175
rect 17868 13132 17920 13141
rect 23848 13132 23900 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2596 12928 2648 12980
rect 3332 12928 3384 12980
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 6000 12928 6052 12980
rect 6736 12928 6788 12980
rect 8484 12928 8536 12980
rect 10324 12928 10376 12980
rect 10784 12971 10836 12980
rect 10784 12937 10793 12971
rect 10793 12937 10827 12971
rect 10827 12937 10836 12971
rect 10784 12928 10836 12937
rect 12348 12928 12400 12980
rect 15384 12928 15436 12980
rect 15660 12928 15712 12980
rect 17776 12971 17828 12980
rect 17776 12937 17785 12971
rect 17785 12937 17819 12971
rect 17819 12937 17828 12971
rect 17776 12928 17828 12937
rect 18144 12971 18196 12980
rect 18144 12937 18153 12971
rect 18153 12937 18187 12971
rect 18187 12937 18196 12971
rect 18144 12928 18196 12937
rect 20812 12971 20864 12980
rect 20812 12937 20821 12971
rect 20821 12937 20855 12971
rect 20855 12937 20864 12971
rect 20812 12928 20864 12937
rect 21272 12971 21324 12980
rect 21272 12937 21281 12971
rect 21281 12937 21315 12971
rect 21315 12937 21324 12971
rect 21272 12928 21324 12937
rect 22744 12971 22796 12980
rect 22744 12937 22753 12971
rect 22753 12937 22787 12971
rect 22787 12937 22796 12971
rect 22744 12928 22796 12937
rect 23388 12928 23440 12980
rect 2412 12860 2464 12912
rect 2780 12792 2832 12844
rect 3056 12792 3108 12844
rect 3332 12792 3384 12844
rect 3976 12792 4028 12844
rect 4252 12835 4304 12844
rect 2504 12724 2556 12776
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 4620 12792 4672 12844
rect 5264 12792 5316 12844
rect 8392 12860 8444 12912
rect 12900 12860 12952 12912
rect 18972 12860 19024 12912
rect 19432 12860 19484 12912
rect 20628 12860 20680 12912
rect 25596 12928 25648 12980
rect 2228 12656 2280 12708
rect 2872 12656 2924 12708
rect 3700 12656 3752 12708
rect 4344 12656 4396 12708
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 9036 12792 9088 12844
rect 11336 12792 11388 12844
rect 11612 12792 11664 12844
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 13544 12792 13596 12844
rect 14004 12792 14056 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 19064 12792 19116 12844
rect 22008 12792 22060 12844
rect 23112 12792 23164 12844
rect 9404 12724 9456 12776
rect 12256 12724 12308 12776
rect 12440 12724 12492 12776
rect 13084 12724 13136 12776
rect 13360 12724 13412 12776
rect 17868 12724 17920 12776
rect 18420 12724 18472 12776
rect 19432 12724 19484 12776
rect 20168 12767 20220 12776
rect 20168 12733 20177 12767
rect 20177 12733 20211 12767
rect 20211 12733 20220 12767
rect 20168 12724 20220 12733
rect 23848 12767 23900 12776
rect 23848 12733 23857 12767
rect 23857 12733 23891 12767
rect 23891 12733 23900 12767
rect 23848 12724 23900 12733
rect 2412 12588 2464 12640
rect 5172 12588 5224 12640
rect 6368 12588 6420 12640
rect 7932 12588 7984 12640
rect 10140 12588 10192 12640
rect 10784 12588 10836 12640
rect 11060 12588 11112 12640
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 12992 12656 13044 12708
rect 14372 12656 14424 12708
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 15476 12588 15528 12640
rect 16580 12631 16632 12640
rect 16580 12597 16589 12631
rect 16589 12597 16623 12631
rect 16623 12597 16632 12631
rect 16580 12588 16632 12597
rect 19432 12588 19484 12640
rect 21824 12656 21876 12708
rect 22008 12656 22060 12708
rect 24216 12656 24268 12708
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 21364 12588 21416 12640
rect 23572 12588 23624 12640
rect 24768 12588 24820 12640
rect 24860 12588 24912 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 2320 12384 2372 12436
rect 2688 12384 2740 12436
rect 3240 12384 3292 12436
rect 3700 12427 3752 12436
rect 3700 12393 3709 12427
rect 3709 12393 3743 12427
rect 3743 12393 3752 12427
rect 3700 12384 3752 12393
rect 3884 12384 3936 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 7380 12427 7432 12436
rect 7380 12393 7389 12427
rect 7389 12393 7423 12427
rect 7423 12393 7432 12427
rect 7380 12384 7432 12393
rect 8576 12384 8628 12436
rect 9404 12427 9456 12436
rect 9404 12393 9413 12427
rect 9413 12393 9447 12427
rect 9447 12393 9456 12427
rect 9404 12384 9456 12393
rect 10692 12384 10744 12436
rect 11796 12384 11848 12436
rect 12900 12384 12952 12436
rect 13820 12384 13872 12436
rect 2964 12316 3016 12368
rect 5448 12316 5500 12368
rect 6828 12359 6880 12368
rect 6828 12325 6837 12359
rect 6837 12325 6871 12359
rect 6871 12325 6880 12359
rect 6828 12316 6880 12325
rect 7840 12359 7892 12368
rect 7840 12325 7849 12359
rect 7849 12325 7883 12359
rect 7883 12325 7892 12359
rect 7840 12316 7892 12325
rect 8852 12316 8904 12368
rect 10876 12316 10928 12368
rect 2320 12248 2372 12300
rect 2596 12248 2648 12300
rect 3056 12248 3108 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 11336 12316 11388 12368
rect 12992 12359 13044 12368
rect 12992 12325 13001 12359
rect 13001 12325 13035 12359
rect 13035 12325 13044 12359
rect 12992 12316 13044 12325
rect 14280 12384 14332 12436
rect 14556 12384 14608 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 15476 12384 15528 12436
rect 16764 12384 16816 12436
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 18788 12384 18840 12436
rect 21272 12384 21324 12436
rect 21732 12384 21784 12436
rect 22744 12427 22796 12436
rect 22744 12393 22753 12427
rect 22753 12393 22787 12427
rect 22787 12393 22796 12427
rect 22744 12384 22796 12393
rect 23756 12384 23808 12436
rect 24768 12384 24820 12436
rect 15568 12316 15620 12368
rect 11060 12248 11112 12300
rect 13084 12248 13136 12300
rect 13728 12248 13780 12300
rect 14556 12248 14608 12300
rect 16580 12316 16632 12368
rect 19064 12316 19116 12368
rect 24860 12316 24912 12368
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 17040 12248 17092 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 17592 12248 17644 12300
rect 18420 12248 18472 12300
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 21824 12248 21876 12300
rect 22928 12248 22980 12300
rect 4712 12223 4764 12232
rect 2780 12112 2832 12164
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 7932 12180 7984 12232
rect 8116 12180 8168 12232
rect 10784 12180 10836 12232
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14004 12223 14056 12232
rect 14004 12189 14013 12223
rect 14013 12189 14047 12223
rect 14047 12189 14056 12223
rect 14004 12180 14056 12189
rect 15844 12223 15896 12232
rect 15844 12189 15853 12223
rect 15853 12189 15887 12223
rect 15887 12189 15896 12223
rect 15844 12180 15896 12189
rect 16304 12180 16356 12232
rect 16764 12180 16816 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 4252 12112 4304 12164
rect 14832 12112 14884 12164
rect 2412 12044 2464 12096
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 14372 12044 14424 12096
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 20076 12044 20128 12096
rect 20904 12044 20956 12096
rect 21364 12044 21416 12096
rect 23848 12044 23900 12096
rect 24032 12044 24084 12096
rect 25044 12087 25096 12096
rect 25044 12053 25053 12087
rect 25053 12053 25087 12087
rect 25087 12053 25096 12087
rect 25044 12044 25096 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 2228 11840 2280 11892
rect 1676 11636 1728 11688
rect 2964 11840 3016 11892
rect 4712 11840 4764 11892
rect 7748 11840 7800 11892
rect 7840 11883 7892 11892
rect 7840 11849 7849 11883
rect 7849 11849 7883 11883
rect 7883 11849 7892 11883
rect 8116 11883 8168 11892
rect 7840 11840 7892 11849
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 11060 11840 11112 11892
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 12808 11840 12860 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 2596 11772 2648 11824
rect 4620 11772 4672 11824
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 12716 11772 12768 11824
rect 3148 11704 3200 11713
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11704 11704 11756 11756
rect 13084 11747 13136 11756
rect 13084 11713 13093 11747
rect 13093 11713 13127 11747
rect 13127 11713 13136 11747
rect 13084 11704 13136 11713
rect 14004 11704 14056 11756
rect 14556 11704 14608 11756
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 4436 11636 4488 11688
rect 2596 11568 2648 11620
rect 4528 11611 4580 11620
rect 4528 11577 4537 11611
rect 4537 11577 4571 11611
rect 4571 11577 4580 11611
rect 4528 11568 4580 11577
rect 12072 11636 12124 11688
rect 16304 11840 16356 11892
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 21272 11883 21324 11892
rect 18420 11840 18472 11849
rect 15200 11747 15252 11756
rect 15200 11713 15209 11747
rect 15209 11713 15243 11747
rect 15243 11713 15252 11747
rect 15200 11704 15252 11713
rect 16028 11704 16080 11756
rect 16488 11704 16540 11756
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 21548 11883 21600 11892
rect 21548 11849 21557 11883
rect 21557 11849 21591 11883
rect 21591 11849 21600 11883
rect 21548 11840 21600 11849
rect 21824 11840 21876 11892
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 23020 11840 23072 11892
rect 19524 11747 19576 11756
rect 19524 11713 19533 11747
rect 19533 11713 19567 11747
rect 19567 11713 19576 11747
rect 19524 11704 19576 11713
rect 24952 11840 25004 11892
rect 25136 11840 25188 11892
rect 24032 11772 24084 11824
rect 24860 11704 24912 11756
rect 2136 11500 2188 11552
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 3424 11500 3476 11552
rect 4988 11500 5040 11552
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11704 11500 11756 11552
rect 13728 11568 13780 11620
rect 12348 11500 12400 11552
rect 14832 11568 14884 11620
rect 21272 11636 21324 11688
rect 22284 11636 22336 11688
rect 25504 11679 25556 11688
rect 25504 11645 25513 11679
rect 25513 11645 25547 11679
rect 25547 11645 25556 11679
rect 25504 11636 25556 11645
rect 15292 11500 15344 11552
rect 17960 11568 18012 11620
rect 24032 11568 24084 11620
rect 17040 11500 17092 11552
rect 17592 11543 17644 11552
rect 17592 11509 17601 11543
rect 17601 11509 17635 11543
rect 17635 11509 17644 11543
rect 17592 11500 17644 11509
rect 18788 11500 18840 11552
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23940 11500 23992 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2412 11339 2464 11348
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 2596 11296 2648 11348
rect 2872 11296 2924 11348
rect 3608 11296 3660 11348
rect 4528 11296 4580 11348
rect 11704 11296 11756 11348
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 12440 11296 12492 11348
rect 13176 11296 13228 11348
rect 13820 11296 13872 11348
rect 14280 11296 14332 11348
rect 15200 11296 15252 11348
rect 15752 11296 15804 11348
rect 16856 11339 16908 11348
rect 16856 11305 16865 11339
rect 16865 11305 16899 11339
rect 16899 11305 16908 11339
rect 16856 11296 16908 11305
rect 18880 11296 18932 11348
rect 20904 11339 20956 11348
rect 20904 11305 20913 11339
rect 20913 11305 20947 11339
rect 20947 11305 20956 11339
rect 20904 11296 20956 11305
rect 22100 11339 22152 11348
rect 22100 11305 22109 11339
rect 22109 11305 22143 11339
rect 22143 11305 22152 11339
rect 22100 11296 22152 11305
rect 23572 11296 23624 11348
rect 24124 11296 24176 11348
rect 3148 11228 3200 11280
rect 11152 11228 11204 11280
rect 13084 11271 13136 11280
rect 13084 11237 13093 11271
rect 13093 11237 13127 11271
rect 13127 11237 13136 11271
rect 13084 11228 13136 11237
rect 15844 11228 15896 11280
rect 16212 11228 16264 11280
rect 16764 11271 16816 11280
rect 16764 11237 16773 11271
rect 16773 11237 16807 11271
rect 16807 11237 16816 11271
rect 16764 11228 16816 11237
rect 18972 11228 19024 11280
rect 24492 11228 24544 11280
rect 3056 11160 3108 11212
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 12808 11160 12860 11212
rect 15660 11203 15712 11212
rect 2872 11092 2924 11144
rect 3240 11092 3292 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 13820 11092 13872 11144
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 16856 11160 16908 11212
rect 18788 11160 18840 11212
rect 21916 11203 21968 11212
rect 21916 11169 21925 11203
rect 21925 11169 21959 11203
rect 21959 11169 21968 11203
rect 21916 11160 21968 11169
rect 22560 11160 22612 11212
rect 23112 11160 23164 11212
rect 24124 11160 24176 11212
rect 24584 11203 24636 11212
rect 24584 11169 24593 11203
rect 24593 11169 24627 11203
rect 24627 11169 24636 11203
rect 24584 11160 24636 11169
rect 24860 11160 24912 11212
rect 15476 11092 15528 11144
rect 10968 11024 11020 11076
rect 11980 11024 12032 11076
rect 16028 11092 16080 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17684 11092 17736 11144
rect 24952 11092 25004 11144
rect 16120 11024 16172 11076
rect 16304 11024 16356 11076
rect 16488 11024 16540 11076
rect 17960 11067 18012 11076
rect 17960 11033 17969 11067
rect 17969 11033 18003 11067
rect 18003 11033 18012 11067
rect 17960 11024 18012 11033
rect 11336 10956 11388 11008
rect 14280 10956 14332 11008
rect 22560 10956 22612 11008
rect 23940 10999 23992 11008
rect 23940 10965 23949 10999
rect 23949 10965 23983 10999
rect 23983 10965 23992 10999
rect 23940 10956 23992 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 2136 10795 2188 10804
rect 2136 10761 2145 10795
rect 2145 10761 2179 10795
rect 2179 10761 2188 10795
rect 2136 10752 2188 10761
rect 2320 10752 2372 10804
rect 2780 10795 2832 10804
rect 2780 10761 2789 10795
rect 2789 10761 2823 10795
rect 2823 10761 2832 10795
rect 2780 10752 2832 10761
rect 12808 10752 12860 10804
rect 13728 10752 13780 10804
rect 14740 10752 14792 10804
rect 1952 10684 2004 10736
rect 572 10616 624 10668
rect 6000 10616 6052 10668
rect 11888 10616 11940 10668
rect 12716 10616 12768 10668
rect 14648 10684 14700 10736
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 15660 10752 15712 10804
rect 16028 10752 16080 10804
rect 17684 10795 17736 10804
rect 17684 10761 17693 10795
rect 17693 10761 17727 10795
rect 17727 10761 17736 10795
rect 17684 10752 17736 10761
rect 21916 10795 21968 10804
rect 21916 10761 21925 10795
rect 21925 10761 21959 10795
rect 21959 10761 21968 10795
rect 21916 10752 21968 10761
rect 23112 10795 23164 10804
rect 23112 10761 23121 10795
rect 23121 10761 23155 10795
rect 23155 10761 23164 10795
rect 23112 10752 23164 10761
rect 23664 10752 23716 10804
rect 24860 10752 24912 10804
rect 23940 10684 23992 10736
rect 26148 10684 26200 10736
rect 16212 10616 16264 10668
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 13912 10480 13964 10532
rect 14004 10480 14056 10532
rect 15384 10480 15436 10532
rect 12348 10412 12400 10464
rect 13820 10455 13872 10464
rect 13820 10421 13829 10455
rect 13829 10421 13863 10455
rect 13863 10421 13872 10455
rect 13820 10412 13872 10421
rect 15752 10455 15804 10464
rect 15752 10421 15761 10455
rect 15761 10421 15795 10455
rect 15795 10421 15804 10455
rect 15752 10412 15804 10421
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17316 10455 17368 10464
rect 17316 10421 17325 10455
rect 17325 10421 17359 10455
rect 17359 10421 17368 10455
rect 17316 10412 17368 10421
rect 24400 10455 24452 10464
rect 24400 10421 24409 10455
rect 24409 10421 24443 10455
rect 24443 10421 24452 10455
rect 24400 10412 24452 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 12624 10208 12676 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 13176 10251 13228 10260
rect 13176 10217 13185 10251
rect 13185 10217 13219 10251
rect 13219 10217 13228 10251
rect 13176 10208 13228 10217
rect 13820 10208 13872 10260
rect 15292 10251 15344 10260
rect 15292 10217 15301 10251
rect 15301 10217 15335 10251
rect 15335 10217 15344 10251
rect 15292 10208 15344 10217
rect 16120 10251 16172 10260
rect 16120 10217 16129 10251
rect 16129 10217 16163 10251
rect 16163 10217 16172 10251
rect 16120 10208 16172 10217
rect 22836 10208 22888 10260
rect 24676 10208 24728 10260
rect 14004 10140 14056 10192
rect 16212 10140 16264 10192
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 17684 10072 17736 10124
rect 23480 10115 23532 10124
rect 23480 10081 23489 10115
rect 23489 10081 23523 10115
rect 23523 10081 23532 10115
rect 23480 10072 23532 10081
rect 23756 10072 23808 10124
rect 24952 10072 25004 10124
rect 13636 10004 13688 10056
rect 14004 9936 14056 9988
rect 14372 9936 14424 9988
rect 25780 9936 25832 9988
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 13084 9664 13136 9716
rect 15660 9664 15712 9716
rect 23756 9664 23808 9716
rect 13636 9596 13688 9648
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 14280 9596 14332 9648
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 16488 9596 16540 9648
rect 24952 9664 25004 9716
rect 14096 9528 14148 9537
rect 22744 9528 22796 9580
rect 23756 9528 23808 9580
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 13912 9460 13964 9512
rect 23940 9324 23992 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 13912 9120 13964 9172
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 24952 8984 25004 9036
rect 25412 8984 25464 9036
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 24124 8619 24176 8628
rect 24124 8585 24133 8619
rect 24133 8585 24167 8619
rect 24167 8585 24176 8619
rect 24124 8576 24176 8585
rect 24952 8619 25004 8628
rect 24952 8585 24961 8619
rect 24961 8585 24995 8619
rect 24995 8585 25004 8619
rect 24952 8576 25004 8585
rect 19984 8508 20036 8560
rect 24676 8508 24728 8560
rect 23940 8415 23992 8424
rect 23940 8381 23949 8415
rect 23949 8381 23983 8415
rect 23983 8381 23992 8415
rect 23940 8372 23992 8381
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 24676 5899 24728 5908
rect 24676 5865 24685 5899
rect 24685 5865 24719 5899
rect 24719 5865 24728 5899
rect 24676 5856 24728 5865
rect 24492 5763 24544 5772
rect 24492 5729 24501 5763
rect 24501 5729 24535 5763
rect 24535 5729 24544 5763
rect 24492 5720 24544 5729
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 24676 5312 24728 5364
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 24032 4768 24084 4820
rect 24676 4700 24728 4752
rect 24492 4675 24544 4684
rect 24492 4641 24501 4675
rect 24501 4641 24535 4675
rect 24535 4641 24544 4675
rect 24492 4632 24544 4641
rect 24216 4564 24268 4616
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 24124 4267 24176 4276
rect 24124 4233 24133 4267
rect 24133 4233 24167 4267
rect 24167 4233 24176 4267
rect 24124 4224 24176 4233
rect 24216 4156 24268 4208
rect 24584 3927 24636 3936
rect 24584 3893 24593 3927
rect 24593 3893 24627 3927
rect 24627 3893 24636 3927
rect 24584 3884 24636 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 11980 2635 12032 2644
rect 11980 2601 11989 2635
rect 11989 2601 12023 2635
rect 12023 2601 12032 2635
rect 11980 2592 12032 2601
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 14004 2635 14056 2644
rect 12440 2592 12492 2601
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 18512 2363 18564 2372
rect 18512 2329 18521 2363
rect 18521 2329 18555 2363
rect 18555 2329 18564 2363
rect 18512 2320 18564 2329
rect 19524 2252 19576 2304
rect 25136 2252 25188 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 1950 27520 2006 28000
rect 2502 27520 2558 28000
rect 3054 27520 3110 28000
rect 3606 27520 3662 28000
rect 4066 27704 4122 27713
rect 4066 27639 4122 27648
rect 308 24410 336 27520
rect 860 27418 888 27520
rect 768 27390 888 27418
rect 296 24404 348 24410
rect 296 24346 348 24352
rect 570 23488 626 23497
rect 570 23423 626 23432
rect 584 22778 612 23423
rect 572 22772 624 22778
rect 572 22714 624 22720
rect 768 15065 796 27390
rect 1412 25242 1440 27520
rect 1412 25214 1900 25242
rect 1584 25152 1636 25158
rect 1584 25094 1636 25100
rect 1676 25152 1728 25158
rect 1676 25094 1728 25100
rect 1400 24608 1452 24614
rect 1400 24550 1452 24556
rect 1308 24404 1360 24410
rect 1308 24346 1360 24352
rect 754 15056 810 15065
rect 754 14991 810 15000
rect 570 10704 626 10713
rect 570 10639 572 10648
rect 624 10639 626 10648
rect 572 10610 624 10616
rect 570 7304 626 7313
rect 570 7239 626 7248
rect 584 7041 612 7239
rect 570 7032 626 7041
rect 570 6967 626 6976
rect 1320 2417 1348 24346
rect 1412 22273 1440 24550
rect 1492 24064 1544 24070
rect 1596 24041 1624 25094
rect 1688 24614 1716 25094
rect 1676 24608 1728 24614
rect 1676 24550 1728 24556
rect 1492 24006 1544 24012
rect 1582 24032 1638 24041
rect 1398 22264 1454 22273
rect 1398 22199 1454 22208
rect 1400 22160 1452 22166
rect 1398 22128 1400 22137
rect 1452 22128 1454 22137
rect 1398 22063 1454 22072
rect 1504 21593 1532 24006
rect 1582 23967 1638 23976
rect 1490 21584 1546 21593
rect 1490 21519 1546 21528
rect 1492 21344 1544 21350
rect 1398 21312 1454 21321
rect 1492 21286 1544 21292
rect 1398 21247 1454 21256
rect 1412 21146 1440 21247
rect 1504 21185 1532 21286
rect 1490 21176 1546 21185
rect 1400 21140 1452 21146
rect 1490 21111 1546 21120
rect 1400 21082 1452 21088
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1596 19825 1624 20198
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 1688 19360 1716 24550
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1780 22681 1808 23054
rect 1766 22672 1822 22681
rect 1766 22607 1822 22616
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 1780 21729 1808 22442
rect 1766 21720 1822 21729
rect 1766 21655 1822 21664
rect 1596 19332 1716 19360
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1412 17882 1440 19246
rect 1400 17876 1452 17882
rect 1400 17818 1452 17824
rect 1490 16552 1546 16561
rect 1490 16487 1546 16496
rect 1504 14498 1532 16487
rect 1596 15609 1624 19332
rect 1676 19236 1728 19242
rect 1676 19178 1728 19184
rect 1688 17785 1716 19178
rect 1872 18873 1900 25214
rect 1964 25129 1992 27520
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 1950 25120 2006 25129
rect 1950 25055 2006 25064
rect 2044 24744 2096 24750
rect 2044 24686 2096 24692
rect 1952 24268 2004 24274
rect 1952 24210 2004 24216
rect 1964 23526 1992 24210
rect 2056 24206 2084 24686
rect 2240 24614 2268 25298
rect 2516 24698 2544 27520
rect 3068 25702 3096 27520
rect 3330 27160 3386 27169
rect 3330 27095 3386 27104
rect 3344 26314 3372 27095
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 3620 25809 3648 27520
rect 4080 27146 4108 27639
rect 4158 27520 4214 28000
rect 4710 27520 4766 28000
rect 5262 27520 5318 28000
rect 5814 27520 5870 28000
rect 6366 27520 6422 28000
rect 6918 27520 6974 28000
rect 7562 27520 7618 28000
rect 8114 27520 8170 28000
rect 8666 27520 8722 28000
rect 9218 27520 9274 28000
rect 9770 27520 9826 28000
rect 10322 27520 10378 28000
rect 10874 27520 10930 28000
rect 11426 27520 11482 28000
rect 11978 27520 12034 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 15934 27520 15990 28000
rect 16486 27520 16542 28000
rect 17038 27520 17094 28000
rect 17590 27520 17646 28000
rect 18142 27520 18198 28000
rect 18694 27520 18750 28000
rect 19246 27520 19302 28000
rect 19798 27520 19854 28000
rect 20350 27520 20406 28000
rect 20902 27520 20958 28000
rect 21546 27520 21602 28000
rect 22098 27520 22154 28000
rect 22650 27520 22706 28000
rect 23202 27520 23258 28000
rect 23754 27520 23810 28000
rect 24306 27520 24362 28000
rect 24858 27520 24914 28000
rect 25410 27520 25466 28000
rect 25686 27704 25742 27713
rect 25686 27639 25742 27648
rect 4172 27418 4200 27520
rect 4172 27390 4292 27418
rect 4080 27118 4200 27146
rect 3790 26480 3846 26489
rect 3790 26415 3846 26424
rect 3606 25800 3662 25809
rect 3606 25735 3662 25744
rect 3056 25696 3108 25702
rect 3056 25638 3108 25644
rect 3516 25356 3568 25362
rect 3516 25298 3568 25304
rect 2778 25256 2834 25265
rect 2778 25191 2780 25200
rect 2832 25191 2834 25200
rect 2780 25162 2832 25168
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 2424 24670 2544 24698
rect 2686 24712 2742 24721
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2044 24200 2096 24206
rect 2042 24168 2044 24177
rect 2096 24168 2098 24177
rect 2042 24103 2098 24112
rect 1952 23520 2004 23526
rect 1952 23462 2004 23468
rect 1964 21298 1992 23462
rect 2042 22536 2098 22545
rect 2042 22471 2098 22480
rect 2056 22098 2084 22471
rect 2044 22092 2096 22098
rect 2044 22034 2096 22040
rect 2056 21418 2084 22034
rect 2044 21412 2096 21418
rect 2044 21354 2096 21360
rect 2136 21344 2188 21350
rect 1964 21292 2136 21298
rect 1964 21286 2188 21292
rect 1964 21270 2176 21286
rect 2148 20806 2176 21270
rect 2136 20800 2188 20806
rect 2240 20777 2268 24550
rect 2424 23066 2452 24670
rect 2686 24647 2742 24656
rect 2700 24614 2728 24647
rect 2688 24608 2740 24614
rect 2502 24576 2558 24585
rect 2688 24550 2740 24556
rect 2502 24511 2558 24520
rect 2516 24274 2544 24511
rect 2504 24268 2556 24274
rect 2504 24210 2556 24216
rect 2516 23866 2544 24210
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2504 23860 2556 23866
rect 2504 23802 2556 23808
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 2608 23089 2636 23122
rect 2594 23080 2650 23089
rect 2424 23038 2544 23066
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2424 22574 2452 22918
rect 2412 22568 2464 22574
rect 2412 22510 2464 22516
rect 2424 22234 2452 22510
rect 2412 22228 2464 22234
rect 2412 22170 2464 22176
rect 2516 22114 2544 23038
rect 2594 23015 2650 23024
rect 2792 22817 2820 24006
rect 2976 23866 3004 25094
rect 3424 24744 3476 24750
rect 3424 24686 3476 24692
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2976 23662 3004 23802
rect 2964 23656 3016 23662
rect 2964 23598 3016 23604
rect 3332 23180 3384 23186
rect 3332 23122 3384 23128
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2778 22808 2834 22817
rect 2778 22743 2834 22752
rect 2780 22568 2832 22574
rect 2780 22510 2832 22516
rect 2424 22086 2544 22114
rect 2320 21616 2372 21622
rect 2320 21558 2372 21564
rect 2332 21146 2360 21558
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2136 20742 2188 20748
rect 2226 20768 2282 20777
rect 2044 20256 2096 20262
rect 2042 20224 2044 20233
rect 2096 20224 2098 20233
rect 2042 20159 2098 20168
rect 2148 19514 2176 20742
rect 2226 20703 2282 20712
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2136 19508 2188 19514
rect 2136 19450 2188 19456
rect 1858 18864 1914 18873
rect 1768 18828 1820 18834
rect 1858 18799 1914 18808
rect 1768 18770 1820 18776
rect 1780 18426 1808 18770
rect 1952 18692 2004 18698
rect 1952 18634 2004 18640
rect 1768 18420 1820 18426
rect 1768 18362 1820 18368
rect 1780 18086 1808 18362
rect 1964 18154 1992 18634
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1952 18148 2004 18154
rect 1952 18090 2004 18096
rect 1768 18080 1820 18086
rect 1768 18022 1820 18028
rect 1674 17776 1730 17785
rect 1674 17711 1730 17720
rect 1964 16776 1992 18090
rect 2056 17882 2084 18566
rect 2136 18216 2188 18222
rect 2136 18158 2188 18164
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 1872 16748 1992 16776
rect 1872 16658 1900 16748
rect 2056 16726 2084 17818
rect 2148 17134 2176 18158
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 17649 2268 17682
rect 2226 17640 2282 17649
rect 2226 17575 2282 17584
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2240 16794 2268 17575
rect 2332 17218 2360 20266
rect 2424 18737 2452 22086
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2502 20768 2558 20777
rect 2502 20703 2558 20712
rect 2516 19666 2544 20703
rect 2608 19786 2636 20878
rect 2700 20602 2728 20946
rect 2792 20874 2820 22510
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 2688 20596 2740 20602
rect 2688 20538 2740 20544
rect 2792 20482 2820 20810
rect 2700 20454 2820 20482
rect 2700 19990 2728 20454
rect 2884 20369 2912 22918
rect 2976 22642 3004 23054
rect 2964 22636 3016 22642
rect 3016 22596 3280 22624
rect 2964 22578 3016 22584
rect 2964 22432 3016 22438
rect 2962 22400 2964 22409
rect 3016 22400 3018 22409
rect 2962 22335 3018 22344
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3068 21690 3096 21966
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 3056 21480 3108 21486
rect 3056 21422 3108 21428
rect 3068 20806 3096 21422
rect 3160 21146 3188 22170
rect 3252 21894 3280 22596
rect 3344 22409 3372 23122
rect 3330 22400 3386 22409
rect 3330 22335 3386 22344
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3056 20800 3108 20806
rect 3056 20742 3108 20748
rect 2870 20360 2926 20369
rect 2870 20295 2926 20304
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2976 20058 3004 20198
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 2688 19984 2740 19990
rect 2688 19926 2740 19932
rect 2780 19916 2832 19922
rect 2780 19858 2832 19864
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 2516 19638 2728 19666
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2502 19000 2558 19009
rect 2502 18935 2504 18944
rect 2556 18935 2558 18944
rect 2504 18906 2556 18912
rect 2410 18728 2466 18737
rect 2410 18663 2466 18672
rect 2516 18426 2544 18906
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2424 17338 2452 17614
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2332 17190 2452 17218
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 1582 15600 1638 15609
rect 1582 15535 1638 15544
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1596 14657 1624 14758
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1504 14470 1624 14498
rect 1492 14408 1544 14414
rect 1492 14350 1544 14356
rect 1504 13802 1532 14350
rect 1492 13796 1544 13802
rect 1492 13738 1544 13744
rect 1596 11898 1624 14470
rect 1584 11892 1636 11898
rect 1584 11834 1636 11840
rect 1688 11694 1716 15914
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1780 13190 1808 14418
rect 1872 13530 1900 15982
rect 1964 15706 1992 16594
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1964 15434 1992 15642
rect 1952 15428 2004 15434
rect 1952 15370 2004 15376
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 1952 15088 2004 15094
rect 1952 15030 2004 15036
rect 1964 14090 1992 15030
rect 2056 14822 2084 15302
rect 2240 15026 2268 15914
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2056 14249 2084 14758
rect 2042 14240 2098 14249
rect 2042 14175 2098 14184
rect 1964 14062 2084 14090
rect 2332 14074 2360 15506
rect 2424 15502 2452 17190
rect 2504 17060 2556 17066
rect 2504 17002 2556 17008
rect 2516 16726 2544 17002
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2516 16250 2544 16662
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2516 15502 2544 16186
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2424 15094 2452 15438
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2608 14521 2636 19450
rect 2594 14512 2650 14521
rect 2594 14447 2650 14456
rect 2410 14104 2466 14113
rect 1952 13796 2004 13802
rect 1952 13738 2004 13744
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 11688 1728 11694
rect 1676 11630 1728 11636
rect 1688 11354 1716 11630
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1964 10742 1992 13738
rect 2056 12594 2084 14062
rect 2320 14068 2372 14074
rect 2410 14039 2466 14048
rect 2320 14010 2372 14016
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2240 12714 2268 13330
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2056 12566 2268 12594
rect 2240 11898 2268 12566
rect 2332 12442 2360 14010
rect 2424 13308 2452 14039
rect 2596 14000 2648 14006
rect 2594 13968 2596 13977
rect 2648 13968 2650 13977
rect 2594 13903 2650 13912
rect 2700 13920 2728 19638
rect 2792 18970 2820 19858
rect 2872 19848 2924 19854
rect 2870 19816 2872 19825
rect 2924 19816 2926 19825
rect 2870 19751 2926 19760
rect 2884 19446 2912 19751
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2792 16250 2820 17682
rect 2884 16726 2912 19110
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3238 18048 3294 18057
rect 3238 17983 3294 17992
rect 2964 17536 3016 17542
rect 2964 17478 3016 17484
rect 2976 16794 3004 17478
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 3146 16688 3202 16697
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2884 16046 2912 16662
rect 3146 16623 3202 16632
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 3056 14952 3108 14958
rect 3160 14929 3188 16623
rect 3252 16114 3280 17983
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 3252 15706 3280 16050
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3056 14894 3108 14900
rect 3146 14920 3202 14929
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2792 14278 2820 14826
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 14113 2820 14214
rect 2778 14104 2834 14113
rect 3068 14074 3096 14894
rect 3252 14890 3280 15302
rect 3146 14855 3202 14864
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 2778 14039 2834 14048
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 2962 13968 3018 13977
rect 2700 13892 2820 13920
rect 2962 13903 3018 13912
rect 3146 13968 3202 13977
rect 3146 13903 3202 13912
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2608 13462 2636 13806
rect 2792 13716 2820 13892
rect 2976 13870 3004 13903
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 3056 13728 3108 13734
rect 2792 13688 3004 13716
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 2596 13320 2648 13326
rect 2424 13280 2596 13308
rect 2596 13262 2648 13268
rect 2608 12986 2636 13262
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2412 12912 2464 12918
rect 2412 12854 2464 12860
rect 2424 12646 2452 12854
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2516 12458 2544 12718
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2424 12430 2544 12458
rect 2700 12442 2728 13330
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2688 12436 2740 12442
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 10810 2176 11494
rect 2332 10810 2360 12242
rect 2424 12186 2452 12430
rect 2688 12378 2740 12384
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2424 12158 2544 12186
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2424 11354 2452 12038
rect 2516 11558 2544 12158
rect 2608 11830 2636 12242
rect 2700 12050 2728 12378
rect 2792 12170 2820 12786
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2700 12022 2820 12050
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2596 11620 2648 11626
rect 2596 11562 2648 11568
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2608 11354 2636 11562
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2596 11348 2648 11354
rect 2596 11290 2648 11296
rect 2792 10810 2820 12022
rect 2884 11354 2912 12650
rect 2976 12374 3004 13688
rect 3056 13670 3108 13676
rect 3068 13190 3096 13670
rect 3056 13184 3108 13190
rect 3056 13126 3108 13132
rect 3068 12850 3096 13126
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 3054 12336 3110 12345
rect 2976 11898 3004 12310
rect 3054 12271 3056 12280
rect 3108 12271 3110 12280
rect 3056 12242 3108 12248
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 2778 3496 2834 3505
rect 2778 3431 2834 3440
rect 1306 2408 1362 2417
rect 1306 2343 1362 2352
rect 2792 480 2820 3431
rect 2884 1465 2912 11086
rect 2976 3369 3004 11630
rect 3068 11218 3096 12242
rect 3160 11762 3188 13903
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3252 13530 3280 13738
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3344 12986 3372 18906
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3344 12850 3372 12922
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 3160 11286 3188 11698
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3252 11150 3280 12378
rect 3436 11558 3464 24686
rect 3528 24614 3556 25298
rect 3804 24954 3832 26415
rect 4066 25936 4122 25945
rect 4066 25871 4122 25880
rect 4080 25378 4108 25871
rect 4172 25498 4200 27118
rect 4264 26081 4292 27390
rect 4250 26072 4306 26081
rect 4250 26007 4306 26016
rect 4724 25809 4752 27520
rect 4896 26308 4948 26314
rect 4896 26250 4948 26256
rect 4710 25800 4766 25809
rect 4710 25735 4766 25744
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 4080 25350 4200 25378
rect 3792 24948 3844 24954
rect 3792 24890 3844 24896
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3528 23594 3556 24550
rect 4172 24410 4200 25350
rect 4908 24954 4936 26250
rect 5080 25356 5132 25362
rect 5080 25298 5132 25304
rect 4896 24948 4948 24954
rect 4896 24890 4948 24896
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 3792 24268 3844 24274
rect 3792 24210 3844 24216
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 3620 21486 3648 24006
rect 3804 23730 3832 24210
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 3976 23860 4028 23866
rect 3976 23802 4028 23808
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3988 23662 4016 23802
rect 4172 23730 4200 24006
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 3976 23656 4028 23662
rect 3976 23598 4028 23604
rect 3700 23520 3752 23526
rect 3988 23497 4016 23598
rect 3700 23462 3752 23468
rect 3974 23488 4030 23497
rect 3712 23254 3740 23462
rect 3974 23423 4030 23432
rect 3700 23248 3752 23254
rect 3698 23216 3700 23225
rect 4252 23248 4304 23254
rect 3752 23216 3754 23225
rect 4252 23190 4304 23196
rect 3698 23151 3754 23160
rect 4264 22438 4292 23190
rect 4252 22432 4304 22438
rect 4252 22374 4304 22380
rect 4264 22098 4292 22374
rect 4540 22234 4568 23734
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 3792 21888 3844 21894
rect 3792 21830 3844 21836
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3620 21078 3648 21422
rect 3608 21072 3660 21078
rect 3608 21014 3660 21020
rect 3620 20466 3648 21014
rect 3804 20806 3832 21830
rect 4448 21350 4476 21898
rect 4540 21690 4568 22170
rect 4620 22160 4672 22166
rect 4620 22102 4672 22108
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4448 20942 4476 21286
rect 4632 21185 4660 22102
rect 4618 21176 4674 21185
rect 4618 21111 4620 21120
rect 4672 21111 4674 21120
rect 4620 21082 4672 21088
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 3792 20800 3844 20806
rect 3792 20742 3844 20748
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4264 20534 4292 20742
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3620 20058 3648 20402
rect 3698 20088 3754 20097
rect 3608 20052 3660 20058
rect 3698 20023 3754 20032
rect 3608 19994 3660 20000
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3528 19514 3556 19790
rect 3608 19712 3660 19718
rect 3608 19654 3660 19660
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 18630 3556 19314
rect 3620 19174 3648 19654
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3528 17542 3556 18566
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 3528 17105 3556 17478
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3516 16992 3568 16998
rect 3516 16934 3568 16940
rect 3528 16794 3556 16934
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3528 16590 3556 16730
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 16114 3556 16526
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3514 15872 3570 15881
rect 3514 15807 3570 15816
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 2962 3360 3018 3369
rect 2962 3295 3018 3304
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 2778 0 2834 480
rect 3436 377 3464 11047
rect 3528 2689 3556 15807
rect 3620 12986 3648 19110
rect 3712 15473 3740 20023
rect 4264 19854 4292 20470
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 4618 20224 4674 20233
rect 4252 19848 4304 19854
rect 4252 19790 4304 19796
rect 4264 19310 4292 19790
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 3896 18630 3924 19178
rect 3974 19136 4030 19145
rect 3974 19071 4030 19080
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3790 17912 3846 17921
rect 3790 17847 3846 17856
rect 3698 15464 3754 15473
rect 3698 15399 3754 15408
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3712 12866 3740 15302
rect 3804 14929 3832 17847
rect 3790 14920 3846 14929
rect 3790 14855 3846 14864
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3804 13326 3832 14010
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3620 12838 3740 12866
rect 3620 11354 3648 12838
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3712 12442 3740 12650
rect 3896 12442 3924 18566
rect 3988 15706 4016 19071
rect 4172 18426 4200 19178
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 4080 17898 4108 18022
rect 4080 17870 4200 17898
rect 4172 17746 4200 17870
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 4080 17134 4108 17614
rect 4172 17338 4200 17682
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4068 17128 4120 17134
rect 4264 17116 4292 19246
rect 4356 18902 4384 19654
rect 4344 18896 4396 18902
rect 4344 18838 4396 18844
rect 4120 17088 4292 17116
rect 4068 17070 4120 17076
rect 4080 17005 4108 17070
rect 4066 16144 4122 16153
rect 4066 16079 4122 16088
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3988 15473 4016 15506
rect 3974 15464 4030 15473
rect 3974 15399 4030 15408
rect 3976 14000 4028 14006
rect 3976 13942 4028 13948
rect 3988 13530 4016 13942
rect 4080 13530 4108 16079
rect 4172 15366 4200 17088
rect 4448 16590 4476 20198
rect 4618 20159 4674 20168
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4540 18766 4568 19178
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4632 18408 4660 20159
rect 4724 19825 4752 24550
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 4710 19816 4766 19825
rect 4710 19751 4766 19760
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4724 18970 4752 19654
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4816 18698 4844 20334
rect 4908 19417 4936 24754
rect 5092 24614 5120 25298
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 5092 20097 5120 24550
rect 5276 24426 5304 27520
rect 5828 25242 5856 27520
rect 6276 25288 6328 25294
rect 5828 25214 6224 25242
rect 6276 25230 6328 25236
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 5276 24398 5488 24426
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 5276 23526 5304 24006
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 5184 22030 5212 23462
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5172 21004 5224 21010
rect 5172 20946 5224 20952
rect 5184 20466 5212 20946
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5078 20088 5134 20097
rect 5078 20023 5134 20032
rect 5080 19916 5132 19922
rect 5080 19858 5132 19864
rect 4894 19408 4950 19417
rect 4894 19343 4950 19352
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4632 18380 4844 18408
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 4632 17338 4660 18226
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4448 15706 4476 16526
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13870 4200 14214
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4068 13252 4120 13258
rect 4264 13240 4292 15030
rect 4120 13212 4292 13240
rect 4068 13194 4120 13200
rect 4264 12850 4292 13212
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3698 11656 3754 11665
rect 3698 11591 3754 11600
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 5137 3740 11591
rect 3882 10024 3938 10033
rect 3882 9959 3938 9968
rect 3896 6361 3924 9959
rect 3882 6352 3938 6361
rect 3882 6287 3938 6296
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3988 2938 4016 12786
rect 4264 12170 4292 12786
rect 4356 12714 4384 15098
rect 4540 15042 4568 16730
rect 4618 15464 4674 15473
rect 4618 15399 4674 15408
rect 4448 15014 4568 15042
rect 4448 14249 4476 15014
rect 4632 14770 4660 15399
rect 4540 14742 4660 14770
rect 4434 14240 4490 14249
rect 4434 14175 4490 14184
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4448 12306 4476 14175
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4448 11694 4476 12242
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4066 11248 4122 11257
rect 4066 11183 4122 11192
rect 4080 10577 4108 11183
rect 4448 11121 4476 11630
rect 4540 11626 4568 14742
rect 4618 14648 4674 14657
rect 4618 14583 4674 14592
rect 4632 14550 4660 14583
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4632 13530 4660 14486
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4724 14074 4752 14350
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4816 13705 4844 18380
rect 4908 17338 4936 19343
rect 5092 19310 5120 19858
rect 5080 19304 5132 19310
rect 5080 19246 5132 19252
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4908 17134 4936 17274
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 5000 16046 5028 18022
rect 5092 17338 5120 18906
rect 5172 18896 5224 18902
rect 5172 18838 5224 18844
rect 5184 18426 5212 18838
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16794 5212 16934
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 4988 16040 5040 16046
rect 5276 15994 5304 23462
rect 5354 22672 5410 22681
rect 5354 22607 5410 22616
rect 5368 22574 5396 22607
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5354 21720 5410 21729
rect 5354 21655 5356 21664
rect 5408 21655 5410 21664
rect 5356 21626 5408 21632
rect 5368 21486 5396 21626
rect 5356 21480 5408 21486
rect 5356 21422 5408 21428
rect 5460 19802 5488 24398
rect 6092 24064 6144 24070
rect 6092 24006 6144 24012
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5644 23322 5672 23666
rect 6104 23662 6132 24006
rect 6092 23656 6144 23662
rect 6092 23598 6144 23604
rect 6104 23322 6132 23598
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 6092 23316 6144 23322
rect 6092 23258 6144 23264
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22432 5592 22438
rect 5540 22374 5592 22380
rect 5552 21894 5580 22374
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 6104 21350 6132 22034
rect 5724 21344 5776 21350
rect 6092 21344 6144 21350
rect 5724 21286 5776 21292
rect 6090 21312 6092 21321
rect 6144 21312 6146 21321
rect 5736 21049 5764 21286
rect 6090 21247 6146 21256
rect 5722 21040 5778 21049
rect 5722 20975 5778 20984
rect 6196 20913 6224 25214
rect 6288 24614 6316 25230
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6182 20904 6238 20913
rect 6182 20839 6238 20848
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20262 5580 20402
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5368 19774 5488 19802
rect 5368 16833 5396 19774
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 5460 18766 5488 19654
rect 5552 19514 5580 20198
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 6012 19514 6040 20198
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 6000 19508 6052 19514
rect 6000 19450 6052 19456
rect 6288 18970 6316 24550
rect 6380 24410 6408 27520
rect 6368 24404 6420 24410
rect 6368 24346 6420 24352
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 23905 6408 24210
rect 6828 24064 6880 24070
rect 6828 24006 6880 24012
rect 6366 23896 6422 23905
rect 6366 23831 6368 23840
rect 6420 23831 6422 23840
rect 6368 23802 6420 23808
rect 6368 23588 6420 23594
rect 6368 23530 6420 23536
rect 6380 19961 6408 23530
rect 6840 23526 6868 24006
rect 6828 23520 6880 23526
rect 6828 23462 6880 23468
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6564 22982 6592 23122
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6734 23080 6790 23089
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6564 22234 6592 22918
rect 6656 22438 6684 23054
rect 6734 23015 6736 23024
rect 6788 23015 6790 23024
rect 6736 22986 6788 22992
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 6656 22234 6684 22374
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6840 22030 6868 23462
rect 6932 23225 6960 27520
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7484 24614 7512 25366
rect 7472 24608 7524 24614
rect 7472 24550 7524 24556
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 6918 23216 6974 23225
rect 6918 23151 6974 23160
rect 7300 22574 7328 23258
rect 7392 23118 7420 23462
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 22778 7420 23054
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6828 22024 6880 22030
rect 6828 21966 6880 21972
rect 6472 21146 6500 21966
rect 6840 21690 6868 21966
rect 7300 21894 7328 22510
rect 7392 22166 7420 22714
rect 7484 22522 7512 24550
rect 7576 22624 7604 27520
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7656 25492 7708 25498
rect 7656 25434 7708 25440
rect 7668 24886 7696 25434
rect 7852 25430 7880 25638
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 7656 24880 7708 24886
rect 8128 24834 8156 27520
rect 7656 24822 7708 24828
rect 7668 24721 7696 24822
rect 7944 24806 8156 24834
rect 8680 24834 8708 27520
rect 9128 25152 9180 25158
rect 9128 25094 9180 25100
rect 9140 24886 9168 25094
rect 9128 24880 9180 24886
rect 8680 24806 8892 24834
rect 9128 24822 9180 24828
rect 9232 24834 9260 27520
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 7654 24712 7710 24721
rect 7654 24647 7710 24656
rect 7656 24608 7708 24614
rect 7656 24550 7708 24556
rect 7668 23662 7696 24550
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7576 22596 7788 22624
rect 7484 22494 7604 22522
rect 7472 22432 7524 22438
rect 7472 22374 7524 22380
rect 7380 22160 7432 22166
rect 7380 22102 7432 22108
rect 7288 21888 7340 21894
rect 7288 21830 7340 21836
rect 6828 21684 6880 21690
rect 6828 21626 6880 21632
rect 7300 21554 7328 21830
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 7288 20800 7340 20806
rect 6734 20768 6790 20777
rect 7288 20742 7340 20748
rect 6734 20703 6790 20712
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 20233 6684 20334
rect 6642 20224 6698 20233
rect 6642 20159 6698 20168
rect 6366 19952 6422 19961
rect 6366 19887 6422 19896
rect 6366 19000 6422 19009
rect 6276 18964 6328 18970
rect 6748 18970 6776 20703
rect 7102 20496 7158 20505
rect 7102 20431 7104 20440
rect 7156 20431 7158 20440
rect 7104 20402 7156 20408
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 6840 19378 6868 19654
rect 6918 19544 6974 19553
rect 6918 19479 6974 19488
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 6932 19009 6960 19479
rect 7208 19174 7236 19654
rect 7300 19310 7328 20742
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6918 19000 6974 19009
rect 6366 18935 6422 18944
rect 6736 18964 6788 18970
rect 6276 18906 6328 18912
rect 5448 18760 5500 18766
rect 5448 18702 5500 18708
rect 5446 18592 5502 18601
rect 5502 18550 5580 18578
rect 5446 18527 5502 18536
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 17882 5488 18226
rect 5552 17882 5580 18550
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5722 18184 5778 18193
rect 5722 18119 5724 18128
rect 5776 18119 5778 18128
rect 5724 18090 5776 18096
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5460 17202 5488 17818
rect 6182 17776 6238 17785
rect 6182 17711 6238 17720
rect 6090 17640 6146 17649
rect 6090 17575 6146 17584
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 6104 17338 6132 17575
rect 6196 17338 6224 17711
rect 6274 17640 6330 17649
rect 6274 17575 6330 17584
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5538 16960 5594 16969
rect 5538 16895 5594 16904
rect 5354 16824 5410 16833
rect 5354 16759 5410 16768
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4988 15982 5040 15988
rect 5000 15910 5028 15982
rect 5092 15966 5304 15994
rect 4988 15904 5040 15910
rect 4986 15872 4988 15881
rect 5040 15872 5042 15881
rect 4986 15807 5042 15816
rect 5092 15162 5120 15966
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5184 14618 5212 15846
rect 5262 15464 5318 15473
rect 5262 15399 5318 15408
rect 5276 15162 5304 15399
rect 5368 15366 5396 16526
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5368 14396 5396 15302
rect 5460 14618 5488 15642
rect 5552 15570 5580 16895
rect 6184 16652 6236 16658
rect 6288 16640 6316 17575
rect 6236 16612 6316 16640
rect 6184 16594 6236 16600
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6288 16250 6316 16612
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 6104 15502 6132 16050
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 6104 15026 6132 15438
rect 6288 15094 6316 16186
rect 6276 15088 6328 15094
rect 6276 15030 6328 15036
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 5814 14920 5870 14929
rect 5814 14855 5870 14864
rect 5828 14822 5856 14855
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 6104 14618 6132 14962
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5448 14408 5500 14414
rect 5368 14368 5448 14396
rect 5448 14350 5500 14356
rect 4802 13696 4858 13705
rect 4802 13631 4858 13640
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12986 4660 13330
rect 5460 13326 5488 14350
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 5276 12850 5304 13126
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 4632 11830 4660 12786
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11898 4752 12174
rect 5184 12102 5212 12582
rect 5460 12374 5488 13262
rect 5552 12442 5580 13670
rect 6012 13462 6040 14010
rect 6104 13870 6132 14554
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6288 13569 6316 15030
rect 6274 13560 6330 13569
rect 6274 13495 6330 13504
rect 6000 13456 6052 13462
rect 6000 13398 6052 13404
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 6012 12986 6040 13398
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6380 12646 6408 18935
rect 6918 18935 6974 18944
rect 6736 18906 6788 18912
rect 6748 18834 6776 18906
rect 7208 18902 7236 19110
rect 7196 18896 7248 18902
rect 7196 18838 7248 18844
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6564 18426 6592 18566
rect 6840 18465 6868 18634
rect 6826 18456 6882 18465
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6748 18414 6826 18442
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6564 16726 6592 17682
rect 6748 17678 6776 18414
rect 6826 18391 6882 18400
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 6828 18080 6880 18086
rect 6826 18048 6828 18057
rect 6880 18048 6882 18057
rect 6826 17983 6882 17992
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 7392 17542 7420 18226
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 6748 17105 6776 17478
rect 7012 17264 7064 17270
rect 7010 17232 7012 17241
rect 7064 17232 7066 17241
rect 7010 17167 7066 17176
rect 6734 17096 6790 17105
rect 6734 17031 6790 17040
rect 6748 16794 6776 17031
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6552 16720 6604 16726
rect 6552 16662 6604 16668
rect 6642 16280 6698 16289
rect 6564 16224 6642 16232
rect 6564 16204 6644 16224
rect 6564 15638 6592 16204
rect 6696 16215 6698 16224
rect 6644 16186 6696 16192
rect 6932 16130 6960 16730
rect 6748 16102 6960 16130
rect 7484 16114 7512 22374
rect 7576 20369 7604 22494
rect 7654 22400 7710 22409
rect 7654 22335 7710 22344
rect 7562 20360 7618 20369
rect 7562 20295 7618 20304
rect 7668 19922 7696 22335
rect 7760 22001 7788 22596
rect 7852 22438 7880 23530
rect 7840 22432 7892 22438
rect 7840 22374 7892 22380
rect 7838 22264 7894 22273
rect 7838 22199 7894 22208
rect 7746 21992 7802 22001
rect 7746 21927 7802 21936
rect 7760 21298 7788 21927
rect 7852 21865 7880 22199
rect 7838 21856 7894 21865
rect 7838 21791 7894 21800
rect 7760 21270 7880 21298
rect 7746 21176 7802 21185
rect 7852 21146 7880 21270
rect 7746 21111 7748 21120
rect 7800 21111 7802 21120
rect 7840 21140 7892 21146
rect 7748 21082 7800 21088
rect 7840 21082 7892 21088
rect 7760 20602 7788 21082
rect 7852 20602 7880 21082
rect 7944 21026 7972 24806
rect 8208 24676 8260 24682
rect 8208 24618 8260 24624
rect 8116 24608 8168 24614
rect 8116 24550 8168 24556
rect 8128 24410 8156 24550
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 8036 22098 8064 23598
rect 8128 22273 8156 24346
rect 8220 24070 8248 24618
rect 8760 24608 8812 24614
rect 8760 24550 8812 24556
rect 8484 24268 8536 24274
rect 8484 24210 8536 24216
rect 8208 24064 8260 24070
rect 8208 24006 8260 24012
rect 8220 23633 8248 24006
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8206 23624 8262 23633
rect 8206 23559 8262 23568
rect 8208 23112 8260 23118
rect 8206 23080 8208 23089
rect 8260 23080 8262 23089
rect 8206 23015 8262 23024
rect 8114 22264 8170 22273
rect 8114 22199 8170 22208
rect 8208 22228 8260 22234
rect 8312 22216 8340 23734
rect 8496 23089 8524 24210
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8680 23769 8708 24006
rect 8772 23905 8800 24550
rect 8758 23896 8814 23905
rect 8758 23831 8814 23840
rect 8666 23760 8722 23769
rect 8772 23730 8800 23831
rect 8666 23695 8722 23704
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8576 23248 8628 23254
rect 8574 23216 8576 23225
rect 8628 23216 8630 23225
rect 8574 23151 8630 23160
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8482 23080 8538 23089
rect 8482 23015 8538 23024
rect 8260 22188 8340 22216
rect 8208 22170 8260 22176
rect 8024 22092 8076 22098
rect 8024 22034 8076 22040
rect 8036 21146 8064 22034
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8128 21690 8156 21966
rect 8680 21894 8708 23122
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8668 21888 8720 21894
rect 8668 21830 8720 21836
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8114 21584 8170 21593
rect 8114 21519 8170 21528
rect 8128 21418 8156 21519
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8680 21049 8708 21830
rect 8772 21593 8800 22374
rect 8758 21584 8814 21593
rect 8758 21519 8814 21528
rect 8666 21040 8722 21049
rect 7944 20998 8064 21026
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 7840 19916 7892 19922
rect 7840 19858 7892 19864
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7760 18970 7788 19790
rect 7852 19174 7880 19858
rect 7944 19854 7972 20878
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7944 19446 7972 19790
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7760 18737 7788 18906
rect 7746 18728 7802 18737
rect 7746 18663 7802 18672
rect 7656 18148 7708 18154
rect 7656 18090 7708 18096
rect 7564 18080 7616 18086
rect 7564 18022 7616 18028
rect 7576 17542 7604 18022
rect 7668 17610 7696 18090
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 7576 17377 7604 17478
rect 7562 17368 7618 17377
rect 7562 17303 7618 17312
rect 7472 16108 7524 16114
rect 6748 15706 6776 16102
rect 7472 16050 7524 16056
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6840 15858 6868 15914
rect 6840 15830 7144 15858
rect 6736 15700 6788 15706
rect 6736 15642 6788 15648
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6642 15600 6698 15609
rect 6642 15535 6698 15544
rect 6656 14958 6684 15535
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6748 13258 6776 13874
rect 6932 13802 6960 14758
rect 7024 13938 7052 15370
rect 7116 14618 7144 15830
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7196 14952 7248 14958
rect 7194 14920 7196 14929
rect 7248 14920 7250 14929
rect 7194 14855 7250 14864
rect 7300 14822 7328 15302
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7104 14272 7156 14278
rect 7300 14249 7328 14758
rect 7576 14550 7604 14962
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7104 14214 7156 14220
rect 7286 14240 7342 14249
rect 7116 14074 7144 14214
rect 7286 14175 7342 14184
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7116 13870 7144 14010
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6932 13530 6960 13738
rect 7668 13530 7696 17546
rect 7748 16584 7800 16590
rect 7852 16561 7880 19110
rect 8036 18902 8064 20998
rect 8666 20975 8722 20984
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 8128 19990 8156 20402
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8404 20058 8432 20334
rect 8392 20052 8444 20058
rect 8392 19994 8444 20000
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 8404 19394 8432 19994
rect 8576 19712 8628 19718
rect 8576 19654 8628 19660
rect 8312 19366 8432 19394
rect 8024 18896 8076 18902
rect 8024 18838 8076 18844
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 8128 18426 8156 18770
rect 8312 18766 8340 19366
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8588 18630 8616 19654
rect 8666 19272 8722 19281
rect 8666 19207 8722 19216
rect 8680 19174 8708 19207
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8312 17882 8340 18566
rect 8588 18222 8616 18566
rect 8576 18216 8628 18222
rect 8482 18184 8538 18193
rect 8576 18158 8628 18164
rect 8482 18119 8538 18128
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8036 17785 8064 17818
rect 8022 17776 8078 17785
rect 8022 17711 8078 17720
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7944 17241 7972 17478
rect 7930 17232 7986 17241
rect 7930 17167 7986 17176
rect 8116 17060 8168 17066
rect 8116 17002 8168 17008
rect 8022 16824 8078 16833
rect 8022 16759 8078 16768
rect 7748 16526 7800 16532
rect 7838 16552 7894 16561
rect 7760 16182 7788 16526
rect 7838 16487 7894 16496
rect 7932 16516 7984 16522
rect 7932 16458 7984 16464
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7944 15638 7972 16458
rect 8036 16182 8064 16759
rect 8024 16176 8076 16182
rect 8024 16118 8076 16124
rect 8128 16114 8156 17002
rect 8312 16794 8340 17818
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8404 17610 8432 17682
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 8404 16674 8432 17546
rect 8220 16646 8432 16674
rect 8220 16250 8248 16646
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7944 15162 7972 15574
rect 8128 15570 8156 16050
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8128 15162 8156 15506
rect 8300 15360 8352 15366
rect 8220 15308 8300 15314
rect 8220 15302 8352 15308
rect 8220 15286 8340 15302
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 8220 15026 8248 15286
rect 8496 15026 8524 18119
rect 8588 18034 8616 18158
rect 8680 18154 8708 18634
rect 8668 18148 8720 18154
rect 8668 18090 8720 18096
rect 8588 18006 8708 18034
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8588 17134 8616 17614
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8574 16824 8630 16833
rect 8574 16759 8630 16768
rect 8588 16726 8616 16759
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8574 15328 8630 15337
rect 8574 15263 8630 15272
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14482 8248 14758
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 14074 8248 14418
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8390 13696 8446 13705
rect 8390 13631 8446 13640
rect 8404 13530 8432 13631
rect 8482 13560 8538 13569
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 8392 13524 8444 13530
rect 8588 13530 8616 15263
rect 8482 13495 8538 13504
rect 8576 13524 8628 13530
rect 8392 13466 8444 13472
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12986 6776 13194
rect 7562 13016 7618 13025
rect 6736 12980 6788 12986
rect 7562 12951 7618 12960
rect 6736 12922 6788 12928
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 6840 12374 6868 12718
rect 7576 12481 7604 12951
rect 8404 12918 8432 13466
rect 8496 13326 8524 13495
rect 8576 13466 8628 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12986 8524 13262
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 7932 12640 7984 12646
rect 8404 12617 8432 12854
rect 7932 12582 7984 12588
rect 8390 12608 8446 12617
rect 7562 12472 7618 12481
rect 7380 12436 7432 12442
rect 7562 12407 7618 12416
rect 7380 12378 7432 12384
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 6828 12368 6880 12374
rect 7392 12345 7420 12378
rect 7840 12368 7892 12374
rect 6828 12310 6880 12316
rect 7378 12336 7434 12345
rect 7840 12310 7892 12316
rect 7378 12271 7434 12280
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7760 12209 7788 12242
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4986 11928 5042 11937
rect 4712 11892 4764 11898
rect 4986 11863 5042 11872
rect 4712 11834 4764 11840
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4540 11354 4568 11562
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4632 11218 4660 11766
rect 5000 11558 5028 11863
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4434 11112 4490 11121
rect 4434 11047 4490 11056
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4080 8809 4108 9415
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 4080 7857 4108 8191
rect 4066 7848 4122 7857
rect 4066 7783 4122 7792
rect 3988 2910 4108 2938
rect 3514 2680 3570 2689
rect 3514 2615 3570 2624
rect 4080 921 4108 2910
rect 5184 2145 5212 12038
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 7760 11898 7788 12135
rect 7852 11898 7880 12310
rect 7944 12238 7972 12582
rect 8390 12543 8446 12552
rect 8588 12442 8616 13466
rect 8680 13462 8708 18006
rect 8772 17241 8800 18838
rect 8758 17232 8814 17241
rect 8758 17167 8814 17176
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8772 14618 8800 14894
rect 8760 14612 8812 14618
rect 8760 14554 8812 14560
rect 8772 13802 8800 14554
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8772 13530 8800 13738
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8668 13456 8720 13462
rect 8668 13398 8720 13404
rect 8680 12889 8708 13398
rect 8666 12880 8722 12889
rect 8666 12815 8722 12824
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8864 12374 8892 24806
rect 9036 24608 9088 24614
rect 9034 24576 9036 24585
rect 9088 24576 9090 24585
rect 9034 24511 9090 24520
rect 9034 24168 9090 24177
rect 9034 24103 9090 24112
rect 9048 23866 9076 24103
rect 9036 23860 9088 23866
rect 9036 23802 9088 23808
rect 9048 23526 9076 23802
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 9140 22438 9168 24822
rect 9232 24806 9352 24834
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 19990 9076 20742
rect 9140 20398 9168 21626
rect 9232 20777 9260 24550
rect 9218 20768 9274 20777
rect 9218 20703 9274 20712
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9036 19984 9088 19990
rect 9036 19926 9088 19932
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 8944 19236 8996 19242
rect 8944 19178 8996 19184
rect 8956 16425 8984 19178
rect 9048 19174 9076 19790
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 8942 16416 8998 16425
rect 8942 16351 8998 16360
rect 8852 12368 8904 12374
rect 8850 12336 8852 12345
rect 8904 12336 8906 12345
rect 8850 12271 8906 12280
rect 8864 12245 8892 12271
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8128 11898 8156 12174
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5998 10840 6054 10849
rect 5998 10775 6054 10784
rect 6012 10674 6040 10775
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 8956 10169 8984 16351
rect 9048 12850 9076 19110
rect 9232 18970 9260 19314
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9232 18426 9260 18906
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9140 17814 9168 18090
rect 9128 17808 9180 17814
rect 9128 17750 9180 17756
rect 9232 17678 9260 18362
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 16289 9260 17478
rect 9324 16658 9352 24806
rect 9508 24682 9536 25638
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9678 24712 9734 24721
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 9600 24342 9628 24686
rect 9678 24647 9734 24656
rect 9692 24410 9720 24647
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9588 24336 9640 24342
rect 9586 24304 9588 24313
rect 9640 24304 9642 24313
rect 9586 24239 9642 24248
rect 9600 24213 9628 24239
rect 9680 23656 9732 23662
rect 9680 23598 9732 23604
rect 9586 23488 9642 23497
rect 9586 23423 9642 23432
rect 9600 23322 9628 23423
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9404 22976 9456 22982
rect 9402 22944 9404 22953
rect 9692 22953 9720 23598
rect 9456 22944 9458 22953
rect 9402 22879 9458 22888
rect 9678 22944 9734 22953
rect 9678 22879 9734 22888
rect 9680 22772 9732 22778
rect 9680 22714 9732 22720
rect 9588 21684 9640 21690
rect 9692 21672 9720 22714
rect 9784 22114 9812 27520
rect 10336 25786 10364 27520
rect 10060 25758 10364 25786
rect 10060 24290 10088 25758
rect 10888 25650 10916 27520
rect 10888 25622 11008 25650
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10874 25528 10930 25537
rect 10874 25463 10930 25472
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10336 24682 10364 25298
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9864 24268 9916 24274
rect 10060 24262 10272 24290
rect 9864 24210 9916 24216
rect 9876 23594 9904 24210
rect 9956 24200 10008 24206
rect 9956 24142 10008 24148
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9968 23526 9996 24142
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 9862 23352 9918 23361
rect 9862 23287 9918 23296
rect 9876 23118 9904 23287
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9876 22681 9904 22918
rect 9862 22672 9918 22681
rect 9862 22607 9918 22616
rect 9784 22086 9904 22114
rect 9640 21644 9720 21672
rect 9588 21626 9640 21632
rect 9876 21457 9904 22086
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9402 20360 9458 20369
rect 9402 20295 9458 20304
rect 9416 20262 9444 20295
rect 9404 20256 9456 20262
rect 9508 20233 9536 20810
rect 9772 20256 9824 20262
rect 9404 20198 9456 20204
rect 9494 20224 9550 20233
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9218 16280 9274 16289
rect 9218 16215 9274 16224
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9232 12764 9260 16215
rect 9416 15450 9444 20198
rect 9772 20198 9824 20204
rect 9494 20159 9550 20168
rect 9508 19922 9536 20159
rect 9496 19916 9548 19922
rect 9496 19858 9548 19864
rect 9508 18630 9536 19858
rect 9586 19680 9642 19689
rect 9586 19615 9642 19624
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9508 17542 9536 18566
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9496 17332 9548 17338
rect 9496 17274 9548 17280
rect 9508 16046 9536 17274
rect 9600 16697 9628 19615
rect 9678 17504 9734 17513
rect 9678 17439 9734 17448
rect 9692 17338 9720 17439
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9692 16794 9720 17070
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9586 16688 9642 16697
rect 9586 16623 9642 16632
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9600 16250 9628 16526
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 15706 9536 15982
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9494 15600 9550 15609
rect 9494 15535 9496 15544
rect 9548 15535 9550 15544
rect 9496 15506 9548 15512
rect 9680 15496 9732 15502
rect 9600 15456 9680 15484
rect 9416 15422 9536 15450
rect 9404 12776 9456 12782
rect 9232 12736 9404 12764
rect 9404 12718 9456 12724
rect 9416 12442 9444 12718
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 8942 10160 8998 10169
rect 8942 10095 8998 10104
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 9508 3641 9536 15422
rect 9600 14958 9628 15456
rect 9680 15438 9732 15444
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9600 13161 9628 13806
rect 9784 13530 9812 20198
rect 9876 19310 9904 21383
rect 9968 19553 9996 23462
rect 10060 22778 10088 24074
rect 10138 23896 10194 23905
rect 10138 23831 10194 23840
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 10152 22234 10180 23831
rect 10244 23633 10272 24262
rect 10704 24177 10732 24550
rect 10690 24168 10746 24177
rect 10690 24103 10746 24112
rect 10796 23730 10824 24618
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10230 23624 10286 23633
rect 10230 23559 10286 23568
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10232 23248 10284 23254
rect 10324 23248 10376 23254
rect 10284 23208 10324 23236
rect 10232 23190 10284 23196
rect 10324 23190 10376 23196
rect 10244 22710 10272 23190
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 10336 22778 10364 23054
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10232 22704 10284 22710
rect 10232 22646 10284 22652
rect 10600 22568 10652 22574
rect 10598 22536 10600 22545
rect 10652 22536 10654 22545
rect 10598 22471 10654 22480
rect 10782 22536 10838 22545
rect 10782 22471 10838 22480
rect 10796 22438 10824 22471
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21060 10088 21966
rect 10152 21690 10180 22170
rect 10508 22024 10560 22030
rect 10506 21992 10508 22001
rect 10692 22024 10744 22030
rect 10560 21992 10562 22001
rect 10692 21966 10744 21972
rect 10506 21927 10562 21936
rect 10520 21690 10548 21927
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10152 21185 10180 21626
rect 10704 21418 10732 21966
rect 10692 21412 10744 21418
rect 10692 21354 10744 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10138 21176 10194 21185
rect 10289 21168 10585 21188
rect 10138 21111 10194 21120
rect 10060 21032 10180 21060
rect 10152 20942 10180 21032
rect 10704 21010 10732 21354
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10796 21185 10824 21286
rect 10782 21176 10838 21185
rect 10782 21111 10838 21120
rect 10692 21004 10744 21010
rect 10692 20946 10744 20952
rect 10140 20936 10192 20942
rect 10046 20904 10102 20913
rect 10140 20878 10192 20884
rect 10046 20839 10102 20848
rect 9954 19544 10010 19553
rect 9954 19479 10010 19488
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 18970 9904 19246
rect 10060 19242 10088 20839
rect 10152 19854 10180 20878
rect 10782 20632 10838 20641
rect 10782 20567 10784 20576
rect 10836 20567 10838 20576
rect 10784 20538 10836 20544
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10048 19236 10100 19242
rect 10048 19178 10100 19184
rect 10690 19136 10746 19145
rect 10289 19068 10585 19088
rect 10690 19071 10746 19080
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 17066 9904 18566
rect 10428 18358 10456 18702
rect 10520 18426 10548 18838
rect 10704 18578 10732 19071
rect 10796 19009 10824 19382
rect 10782 19000 10838 19009
rect 10782 18935 10838 18944
rect 10612 18550 10732 18578
rect 10612 18465 10640 18550
rect 10598 18456 10654 18465
rect 10508 18420 10560 18426
rect 10598 18391 10654 18400
rect 10508 18362 10560 18368
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9968 16726 9996 17682
rect 10152 17338 10180 17818
rect 10140 17332 10192 17338
rect 10060 17292 10140 17320
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9862 16008 9918 16017
rect 9862 15943 9918 15952
rect 9876 15706 9904 15943
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 10060 15337 10088 17292
rect 10140 17274 10192 17280
rect 10796 17134 10824 18022
rect 10888 17882 10916 25463
rect 10980 23322 11008 25622
rect 11440 25514 11468 27520
rect 11702 26072 11758 26081
rect 11702 26007 11758 26016
rect 11612 25764 11664 25770
rect 11612 25706 11664 25712
rect 11256 25486 11468 25514
rect 11624 25498 11652 25706
rect 11612 25492 11664 25498
rect 11152 24608 11204 24614
rect 11150 24576 11152 24585
rect 11204 24576 11206 24585
rect 11150 24511 11206 24520
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11072 23662 11100 24006
rect 11256 23905 11284 25486
rect 11612 25434 11664 25440
rect 11336 25356 11388 25362
rect 11336 25298 11388 25304
rect 11348 24177 11376 25298
rect 11428 24608 11480 24614
rect 11426 24576 11428 24585
rect 11480 24576 11482 24585
rect 11426 24511 11482 24520
rect 11520 24200 11572 24206
rect 11334 24168 11390 24177
rect 11520 24142 11572 24148
rect 11334 24103 11390 24112
rect 11242 23896 11298 23905
rect 11242 23831 11298 23840
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11060 23656 11112 23662
rect 11058 23624 11060 23633
rect 11112 23624 11114 23633
rect 11058 23559 11114 23568
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10968 22976 11020 22982
rect 10968 22918 11020 22924
rect 11152 22976 11204 22982
rect 11152 22918 11204 22924
rect 10980 22574 11008 22918
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 11164 22098 11192 22918
rect 11242 22808 11298 22817
rect 11242 22743 11298 22752
rect 11256 22506 11284 22743
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21554 11284 21830
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11152 21412 11204 21418
rect 11152 21354 11204 21360
rect 11164 21146 11192 21354
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 11164 20602 11192 20946
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11256 20262 11284 20470
rect 11348 20369 11376 23802
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11440 22234 11468 22578
rect 11428 22228 11480 22234
rect 11428 22170 11480 22176
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11334 20360 11390 20369
rect 11334 20295 11390 20304
rect 11244 20256 11296 20262
rect 11058 20224 11114 20233
rect 11244 20198 11296 20204
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 11058 20159 11114 20168
rect 10968 18896 11020 18902
rect 11072 18850 11100 20159
rect 11256 20058 11284 20198
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11348 19689 11376 20198
rect 11440 19990 11468 20402
rect 11428 19984 11480 19990
rect 11428 19926 11480 19932
rect 11334 19680 11390 19689
rect 11334 19615 11390 19624
rect 11440 19514 11468 19926
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11020 18844 11100 18850
rect 10968 18838 11100 18844
rect 10980 18822 11100 18838
rect 11060 18624 11112 18630
rect 10980 18584 11060 18612
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10980 17678 11008 18584
rect 11060 18566 11112 18572
rect 11164 17814 11192 19314
rect 11244 18352 11296 18358
rect 11244 18294 11296 18300
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11256 17746 11284 18294
rect 11426 18184 11482 18193
rect 11426 18119 11482 18128
rect 11440 18086 11468 18119
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17202 10916 17478
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10140 16992 10192 16998
rect 10138 16960 10140 16969
rect 10192 16960 10194 16969
rect 10138 16895 10194 16904
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10138 16824 10194 16833
rect 10289 16816 10585 16836
rect 10888 16794 10916 17002
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10138 16759 10140 16768
rect 10192 16759 10194 16768
rect 10876 16788 10928 16794
rect 10140 16730 10192 16736
rect 10876 16730 10928 16736
rect 10152 16250 10180 16730
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10244 15994 10272 16526
rect 10520 16250 10548 16594
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10152 15966 10272 15994
rect 10152 15706 10180 15966
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10046 15328 10102 15337
rect 10046 15263 10102 15272
rect 10152 14958 10180 15642
rect 10140 14952 10192 14958
rect 10060 14912 10140 14940
rect 10060 14074 10088 14912
rect 10140 14894 10192 14900
rect 10704 14793 10732 16662
rect 10782 16280 10838 16289
rect 10782 16215 10784 16224
rect 10836 16215 10838 16224
rect 10784 16186 10836 16192
rect 10980 16153 11008 16934
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 10796 15706 10824 15914
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 11072 15638 11100 17138
rect 11164 17105 11192 17274
rect 11150 17096 11206 17105
rect 11150 17031 11206 17040
rect 11164 16998 11192 17031
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11256 16658 11284 17682
rect 11428 17060 11480 17066
rect 11428 17002 11480 17008
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11440 16114 11468 17002
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11060 15632 11112 15638
rect 11164 15609 11192 15846
rect 11060 15574 11112 15580
rect 11150 15600 11206 15609
rect 11072 15162 11100 15574
rect 11150 15535 11206 15544
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10690 14784 10746 14793
rect 10289 14716 10585 14736
rect 10690 14719 10746 14728
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 11072 14618 11100 15098
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10140 14544 10192 14550
rect 10138 14512 10140 14521
rect 10192 14512 10194 14521
rect 10138 14447 10194 14456
rect 11336 14272 11388 14278
rect 11242 14240 11298 14249
rect 11336 14214 11388 14220
rect 11242 14175 11298 14184
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 10152 12646 10180 13330
rect 10336 12986 10364 13330
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10690 13152 10746 13161
rect 10690 13087 10746 13096
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10704 12442 10732 13087
rect 10796 12986 10824 13223
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11150 12880 11206 12889
rect 11150 12815 11206 12824
rect 10784 12640 10836 12646
rect 11060 12640 11112 12646
rect 10784 12582 10836 12588
rect 10888 12588 11060 12594
rect 10888 12582 11112 12588
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10796 12238 10824 12582
rect 10888 12566 11100 12582
rect 10888 12374 10916 12566
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10796 10305 10824 11494
rect 10980 11082 11008 12174
rect 11072 11898 11100 12242
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 11164 11286 11192 12815
rect 11256 12481 11284 14175
rect 11348 12850 11376 14214
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11242 12472 11298 12481
rect 11242 12407 11298 12416
rect 11348 12374 11376 12786
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 11348 11014 11376 11698
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 11532 10169 11560 24142
rect 11716 20874 11744 26007
rect 11992 24426 12020 27520
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12072 24676 12124 24682
rect 12072 24618 12124 24624
rect 11808 24398 12020 24426
rect 11704 20868 11756 20874
rect 11704 20810 11756 20816
rect 11808 18834 11836 24398
rect 11888 23248 11940 23254
rect 11888 23190 11940 23196
rect 11900 22778 11928 23190
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11900 22114 11928 22714
rect 11900 22086 12020 22114
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11900 21350 11928 21490
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 21146 11928 21286
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11900 20466 11928 21082
rect 11992 20942 12020 22086
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11978 20224 12034 20233
rect 11978 20159 12034 20168
rect 11992 20058 12020 20159
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11796 18828 11848 18834
rect 11796 18770 11848 18776
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11624 13433 11652 18294
rect 11808 17921 11836 18770
rect 11992 18737 12020 19110
rect 11978 18728 12034 18737
rect 11978 18663 12034 18672
rect 11886 18320 11942 18329
rect 11886 18255 11888 18264
rect 11940 18255 11942 18264
rect 11888 18226 11940 18232
rect 11794 17912 11850 17921
rect 11704 17876 11756 17882
rect 11794 17847 11850 17856
rect 11704 17818 11756 17824
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11612 13184 11664 13190
rect 11610 13152 11612 13161
rect 11664 13152 11666 13161
rect 11610 13087 11666 13096
rect 11624 12850 11652 13087
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11716 11762 11744 17818
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11900 16998 11928 17750
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11808 16250 11836 16594
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 13734 11836 14350
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13394 11836 13670
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11808 12889 11836 13330
rect 11794 12880 11850 12889
rect 11794 12815 11796 12824
rect 11848 12815 11850 12824
rect 11796 12786 11848 12792
rect 11808 12442 11836 12786
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11900 10674 11928 16934
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 11801 12020 14826
rect 12084 13802 12112 24618
rect 12268 23254 12296 24890
rect 12544 24818 12572 27520
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12728 24614 12756 25298
rect 13004 25226 13032 25774
rect 12992 25220 13044 25226
rect 12992 25162 13044 25168
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12348 24064 12400 24070
rect 12348 24006 12400 24012
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 18426 12204 22510
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12268 21690 12296 22442
rect 12360 22234 12388 24006
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12452 22982 12480 23598
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22642 12480 22918
rect 12440 22636 12492 22642
rect 12492 22596 12572 22624
rect 12440 22578 12492 22584
rect 12348 22228 12400 22234
rect 12348 22170 12400 22176
rect 12544 22166 12572 22596
rect 12636 22234 12664 24006
rect 12728 23254 12756 24550
rect 12808 24132 12860 24138
rect 12808 24074 12860 24080
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 12820 23594 12848 24074
rect 12808 23588 12860 23594
rect 12808 23530 12860 23536
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12820 22982 12848 23530
rect 13004 23526 13032 24074
rect 12992 23520 13044 23526
rect 12992 23462 13044 23468
rect 13096 23474 13124 27520
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24750 13400 25094
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13372 24274 13400 24550
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13266 23488 13322 23497
rect 13004 23338 13032 23462
rect 13096 23446 13216 23474
rect 13004 23310 13124 23338
rect 12808 22976 12860 22982
rect 12808 22918 12860 22924
rect 12714 22536 12770 22545
rect 12714 22471 12770 22480
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12532 22160 12584 22166
rect 12532 22102 12584 22108
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21690 12480 21966
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12728 21486 12756 22471
rect 12820 21622 12848 22918
rect 12898 22672 12954 22681
rect 12898 22607 12954 22616
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12912 21554 12940 22607
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 13004 22030 13032 22442
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12360 21298 12388 21354
rect 12360 21270 12480 21298
rect 12452 19514 12480 21270
rect 12912 21146 12940 21490
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 13004 21078 13032 21490
rect 13096 21146 13124 23310
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12992 21072 13044 21078
rect 12992 21014 13044 21020
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12820 20534 12848 20946
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12624 19440 12676 19446
rect 12622 19408 12624 19417
rect 12676 19408 12678 19417
rect 12728 19378 12756 20402
rect 12622 19343 12678 19352
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18834 12480 19110
rect 12820 18970 12848 20470
rect 12990 20360 13046 20369
rect 12990 20295 12992 20304
rect 13044 20295 13046 20304
rect 12992 20266 13044 20272
rect 12900 20256 12952 20262
rect 12900 20198 12952 20204
rect 12912 20058 12940 20198
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12360 17746 12388 18634
rect 12452 18630 12480 18770
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18222 12480 18566
rect 12544 18426 12572 18702
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12544 18086 12572 18362
rect 12532 18080 12584 18086
rect 12532 18022 12584 18028
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12360 17202 12388 17682
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12452 16017 12480 16186
rect 12438 16008 12494 16017
rect 12438 15943 12494 15952
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 14618 12296 15846
rect 12544 14958 12572 18022
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16794 12664 17002
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12636 14770 12664 16594
rect 12544 14742 12664 14770
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12360 13870 12388 14486
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12452 14074 12480 14418
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 12646 12204 13330
rect 12256 13252 12308 13258
rect 12256 13194 12308 13200
rect 12268 12782 12296 13194
rect 12360 12986 12388 13806
rect 12544 13734 12572 14742
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13190 12572 13670
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 12084 11354 12112 11630
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11518 10160 11574 10169
rect 11518 10095 11574 10104
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 9494 3632 9550 3641
rect 9494 3567 9550 3576
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5170 2136 5226 2145
rect 5622 2128 5918 2148
rect 5170 2071 5226 2080
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 8312 480 8340 2887
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 11992 2650 12020 11018
rect 12176 3505 12204 12582
rect 12452 11898 12480 12718
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 10577 12388 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12346 10568 12402 10577
rect 12346 10503 12402 10512
rect 12348 10464 12400 10470
rect 12452 10452 12480 11290
rect 12400 10424 12480 10452
rect 12348 10406 12400 10412
rect 12360 10033 12388 10406
rect 12346 10024 12402 10033
rect 12346 9959 12402 9968
rect 12544 8401 12572 13126
rect 12636 10266 12664 14486
rect 12728 11830 12756 18566
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12820 16658 12848 18158
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12806 16144 12862 16153
rect 12806 16079 12808 16088
rect 12860 16079 12862 16088
rect 12912 16096 12940 19994
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13004 16250 13032 19858
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13096 19417 13124 19654
rect 13082 19408 13138 19417
rect 13082 19343 13138 19352
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13096 17218 13124 18906
rect 13188 17338 13216 23446
rect 13266 23423 13322 23432
rect 13280 19922 13308 23423
rect 13372 23322 13400 24210
rect 13360 23316 13412 23322
rect 13360 23258 13412 23264
rect 13358 22672 13414 22681
rect 13358 22607 13414 22616
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 18698 13308 19722
rect 13372 19310 13400 22607
rect 13464 22273 13492 24550
rect 13450 22264 13506 22273
rect 13450 22199 13506 22208
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13280 17814 13308 18634
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13096 17190 13216 17218
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13084 16108 13136 16114
rect 12912 16068 13032 16096
rect 12808 16050 12860 16056
rect 12820 15994 12848 16050
rect 12820 15966 12940 15994
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15162 12848 15846
rect 12912 15706 12940 15966
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13004 15609 13032 16068
rect 13084 16050 13136 16056
rect 12990 15600 13046 15609
rect 12990 15535 13046 15544
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14816 12860 14822
rect 12806 14784 12808 14793
rect 12860 14784 12862 14793
rect 12806 14719 12862 14728
rect 12820 14278 12848 14719
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12912 14090 12940 14894
rect 12820 14062 12940 14090
rect 13004 14074 13032 15535
rect 13096 15434 13124 16050
rect 13188 15745 13216 17190
rect 13266 16688 13322 16697
rect 13266 16623 13322 16632
rect 13174 15736 13230 15745
rect 13174 15671 13230 15680
rect 13084 15428 13136 15434
rect 13084 15370 13136 15376
rect 13096 14414 13124 15370
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15094 13216 15302
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13188 14618 13216 15030
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13280 14550 13308 16623
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13372 14482 13400 15302
rect 13464 14657 13492 22199
rect 13450 14648 13506 14657
rect 13450 14583 13506 14592
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13268 14272 13320 14278
rect 13556 14226 13584 24754
rect 13648 24313 13676 27520
rect 14292 25514 14320 27520
rect 13924 25486 14320 25514
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13634 24304 13690 24313
rect 13634 24239 13690 24248
rect 13648 20058 13676 24239
rect 13832 23866 13860 25094
rect 13924 24290 13952 25486
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 14280 25356 14332 25362
rect 14280 25298 14332 25304
rect 14004 25288 14056 25294
rect 14004 25230 14056 25236
rect 14016 24410 14044 25230
rect 14108 24614 14136 25298
rect 14292 24614 14320 25298
rect 14844 25242 14872 27520
rect 14384 25214 14872 25242
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14108 24449 14136 24550
rect 14094 24440 14150 24449
rect 14004 24404 14056 24410
rect 14094 24375 14150 24384
rect 14004 24346 14056 24352
rect 13924 24262 14136 24290
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13728 22568 13780 22574
rect 13832 22556 13860 23462
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13780 22528 13860 22556
rect 13728 22510 13780 22516
rect 13924 22522 13952 23122
rect 14016 22710 14044 24006
rect 14108 22930 14136 24262
rect 14186 23760 14242 23769
rect 14186 23695 14242 23704
rect 14200 23594 14228 23695
rect 14188 23588 14240 23594
rect 14188 23530 14240 23536
rect 14186 22944 14242 22953
rect 14108 22902 14186 22930
rect 14186 22879 14242 22888
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 14200 22545 14228 22879
rect 14292 22692 14320 24550
rect 14384 22817 14412 25214
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14476 24070 14504 24754
rect 14844 24682 14872 25094
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15198 24848 15254 24857
rect 15198 24783 15254 24792
rect 14832 24676 14884 24682
rect 14832 24618 14884 24624
rect 14556 24608 14608 24614
rect 14556 24550 14608 24556
rect 14740 24608 14792 24614
rect 14740 24550 14792 24556
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14370 22808 14426 22817
rect 14370 22743 14426 22752
rect 14292 22664 14412 22692
rect 14186 22536 14242 22545
rect 13924 22494 14044 22522
rect 14016 22438 14044 22494
rect 14186 22471 14242 22480
rect 13912 22432 13964 22438
rect 13912 22374 13964 22380
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13728 21004 13780 21010
rect 13728 20946 13780 20952
rect 13740 20890 13768 20946
rect 13740 20862 13860 20890
rect 13832 20244 13860 20862
rect 13924 20466 13952 22374
rect 14292 22137 14320 22374
rect 14278 22128 14334 22137
rect 14004 22092 14056 22098
rect 14278 22063 14334 22072
rect 14004 22034 14056 22040
rect 14016 21690 14044 22034
rect 14188 22024 14240 22030
rect 14186 21992 14188 22001
rect 14240 21992 14242 22001
rect 14186 21927 14242 21936
rect 14384 21690 14412 22664
rect 14476 21690 14504 24006
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14016 21350 14044 21490
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 13912 20256 13964 20262
rect 13832 20216 13912 20244
rect 14016 20233 14044 21286
rect 14108 21185 14136 21354
rect 14094 21176 14150 21185
rect 14094 21111 14096 21120
rect 14148 21111 14150 21120
rect 14096 21082 14148 21088
rect 14094 21040 14150 21049
rect 14094 20975 14150 20984
rect 13912 20198 13964 20204
rect 14002 20224 14058 20233
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13648 19514 13676 19994
rect 13728 19916 13780 19922
rect 13728 19858 13780 19864
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13740 19258 13768 19858
rect 13740 19230 13860 19258
rect 13832 19174 13860 19230
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13740 17882 13768 18090
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13832 17610 13860 19110
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13818 17368 13874 17377
rect 13818 17303 13820 17312
rect 13872 17303 13874 17312
rect 13820 17274 13872 17280
rect 13924 16674 13952 20198
rect 14002 20159 14058 20168
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14016 18630 14044 19314
rect 14108 19174 14136 20975
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14016 17513 14044 18566
rect 14108 18465 14136 18566
rect 14094 18456 14150 18465
rect 14094 18391 14150 18400
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14002 17504 14058 17513
rect 14002 17439 14058 17448
rect 13832 16646 13952 16674
rect 14004 16652 14056 16658
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13268 14214 13320 14220
rect 12992 14068 13044 14074
rect 12820 12050 12848 14062
rect 12992 14010 13044 14016
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12912 13870 12940 13942
rect 12900 13864 12952 13870
rect 12898 13832 12900 13841
rect 12952 13832 12954 13841
rect 12898 13767 12954 13776
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12900 12912 12952 12918
rect 12900 12854 12952 12860
rect 12990 12880 13046 12889
rect 12912 12646 12940 12854
rect 12990 12815 12992 12824
rect 13044 12815 13046 12824
rect 12992 12786 13044 12792
rect 13096 12782 13124 13738
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12912 12442 12940 12582
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 13004 12374 13032 12650
rect 12992 12368 13044 12374
rect 12990 12336 12992 12345
rect 13044 12336 13046 12345
rect 12990 12271 13046 12280
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 12820 12022 12940 12050
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12820 11218 12848 11834
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10674 12756 11086
rect 12820 10810 12848 11154
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12530 8392 12586 8401
rect 12530 8327 12586 8336
rect 12912 3505 12940 12022
rect 13096 11762 13124 12242
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13096 11286 13124 11698
rect 13188 11354 13216 14214
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13174 10432 13230 10441
rect 13174 10367 13230 10376
rect 13082 10296 13138 10305
rect 13188 10266 13216 10367
rect 13082 10231 13084 10240
rect 13136 10231 13138 10240
rect 13176 10260 13228 10266
rect 13084 10202 13136 10208
rect 13176 10202 13228 10208
rect 13096 9722 13124 10202
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13188 9586 13216 10202
rect 13280 9897 13308 14214
rect 13372 14198 13584 14226
rect 13372 12782 13400 14198
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13464 12730 13492 14010
rect 13544 13932 13596 13938
rect 13544 13874 13596 13880
rect 13556 13734 13584 13874
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 12850 13584 13670
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13372 12238 13400 12718
rect 13464 12702 13584 12730
rect 13450 12336 13506 12345
rect 13450 12271 13506 12280
rect 13360 12232 13412 12238
rect 13358 12200 13360 12209
rect 13412 12200 13414 12209
rect 13358 12135 13414 12144
rect 13372 12109 13400 12135
rect 13266 9888 13322 9897
rect 13266 9823 13322 9832
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13464 9489 13492 12271
rect 13556 9625 13584 12702
rect 13648 10062 13676 15846
rect 13728 15564 13780 15570
rect 13728 15506 13780 15512
rect 13740 15162 13768 15506
rect 13832 15502 13860 16646
rect 14004 16594 14056 16600
rect 13910 16416 13966 16425
rect 13910 16351 13966 16360
rect 13924 16017 13952 16351
rect 14016 16289 14044 16594
rect 14002 16280 14058 16289
rect 14002 16215 14058 16224
rect 13910 16008 13966 16017
rect 13910 15943 13966 15952
rect 14016 15706 14044 16215
rect 14108 16114 14136 18022
rect 14200 16674 14228 21626
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14278 21040 14334 21049
rect 14278 20975 14334 20984
rect 14292 20942 14320 20975
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14292 20602 14320 20878
rect 14384 20788 14412 21286
rect 14568 21185 14596 24550
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14660 23769 14688 24142
rect 14752 24070 14780 24550
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14646 23760 14702 23769
rect 14646 23695 14702 23704
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14660 21865 14688 21898
rect 14646 21856 14702 21865
rect 14646 21791 14702 21800
rect 14660 21690 14688 21791
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14554 21176 14610 21185
rect 14554 21111 14610 21120
rect 14464 20800 14516 20806
rect 14384 20760 14464 20788
rect 14464 20742 14516 20748
rect 14476 20641 14504 20742
rect 14462 20632 14518 20641
rect 14280 20596 14332 20602
rect 14660 20602 14688 21490
rect 14462 20567 14518 20576
rect 14648 20596 14700 20602
rect 14280 20538 14332 20544
rect 14648 20538 14700 20544
rect 14278 20224 14334 20233
rect 14278 20159 14334 20168
rect 14292 17626 14320 20159
rect 14646 19952 14702 19961
rect 14646 19887 14702 19896
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14370 19272 14426 19281
rect 14370 19207 14372 19216
rect 14424 19207 14426 19216
rect 14372 19178 14424 19184
rect 14384 18970 14412 19178
rect 14476 19174 14504 19654
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14476 17785 14504 19110
rect 14462 17776 14518 17785
rect 14568 17746 14596 19722
rect 14660 18034 14688 19887
rect 14752 19174 14780 24006
rect 14844 22098 14872 24618
rect 15212 24449 15240 24783
rect 15198 24440 15254 24449
rect 15198 24375 15254 24384
rect 15290 24304 15346 24313
rect 15290 24239 15292 24248
rect 15344 24239 15346 24248
rect 15292 24210 15344 24216
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23866 15332 24210
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15290 23352 15346 23361
rect 15290 23287 15346 23296
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15120 22234 15148 22510
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 15304 22098 15332 23287
rect 15396 22681 15424 27520
rect 15948 25537 15976 27520
rect 15934 25528 15990 25537
rect 16500 25498 16528 27520
rect 17052 25498 17080 27520
rect 17498 25936 17554 25945
rect 17498 25871 17554 25880
rect 15934 25463 15990 25472
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 16396 25356 16448 25362
rect 16396 25298 16448 25304
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 15936 25220 15988 25226
rect 15936 25162 15988 25168
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15764 24886 15792 25094
rect 15752 24880 15804 24886
rect 15752 24822 15804 24828
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15856 24614 15884 24686
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15476 24200 15528 24206
rect 15474 24168 15476 24177
rect 15528 24168 15530 24177
rect 15474 24103 15530 24112
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15474 23624 15530 23633
rect 15474 23559 15530 23568
rect 15488 23526 15516 23559
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15382 22672 15438 22681
rect 15382 22607 15438 22616
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15212 21962 15240 22034
rect 15200 21956 15252 21962
rect 15200 21898 15252 21904
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21434 15424 22170
rect 15304 21406 15424 21434
rect 15304 21146 15332 21406
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15292 21140 15344 21146
rect 15292 21082 15344 21088
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14740 18760 14792 18766
rect 14740 18702 14792 18708
rect 14752 18154 14780 18702
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14660 18006 14780 18034
rect 14646 17912 14702 17921
rect 14752 17882 14780 18006
rect 14646 17847 14702 17856
rect 14740 17876 14792 17882
rect 14462 17711 14518 17720
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14292 17598 14504 17626
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14200 16646 14320 16674
rect 14384 16658 14412 16934
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14096 16108 14148 16114
rect 14096 16050 14148 16056
rect 14200 15910 14228 16458
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13740 15065 13768 15098
rect 13726 15056 13782 15065
rect 13726 14991 13782 15000
rect 13740 14278 13768 14991
rect 13832 14906 13860 15438
rect 13924 15026 13952 15438
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13832 14878 13952 14906
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13832 14074 13860 14350
rect 13924 14278 13952 14878
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 14108 14550 14136 14758
rect 14096 14544 14148 14550
rect 14094 14512 14096 14521
rect 14148 14512 14150 14521
rect 14094 14447 14150 14456
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11665 13768 12242
rect 13832 11898 13860 12378
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13726 11656 13782 11665
rect 13726 11591 13728 11600
rect 13780 11591 13782 11600
rect 13728 11562 13780 11568
rect 13740 11531 13768 11562
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13832 11234 13860 11290
rect 13924 11257 13952 14214
rect 14094 13696 14150 13705
rect 14094 13631 14150 13640
rect 14108 13025 14136 13631
rect 14094 13016 14150 13025
rect 14094 12951 14150 12960
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14016 12238 14044 12786
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 14016 11762 14044 12174
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13740 11206 13860 11234
rect 13910 11248 13966 11257
rect 13740 10810 13768 11206
rect 13910 11183 13966 11192
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13832 10470 13860 11086
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10266 13860 10406
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 9654 13676 9998
rect 13636 9648 13688 9654
rect 13542 9616 13598 9625
rect 13636 9590 13688 9596
rect 13542 9551 13598 9560
rect 13924 9518 13952 10474
rect 14016 10198 14044 10474
rect 14004 10192 14056 10198
rect 14004 10134 14056 10140
rect 14004 9988 14056 9994
rect 14004 9930 14056 9936
rect 13912 9512 13964 9518
rect 13450 9480 13506 9489
rect 13912 9454 13964 9460
rect 13450 9415 13506 9424
rect 13924 9178 13952 9454
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13910 3632 13966 3641
rect 13910 3567 13966 3576
rect 12162 3496 12218 3505
rect 12162 3431 12218 3440
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 12438 2952 12494 2961
rect 12438 2887 12494 2896
rect 12452 2650 12480 2887
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 13924 480 13952 3567
rect 14016 2650 14044 9930
rect 14108 9586 14136 12951
rect 14200 9654 14228 15846
rect 14292 14074 14320 16646
rect 14372 16652 14424 16658
rect 14372 16594 14424 16600
rect 14384 16250 14412 16594
rect 14476 16561 14504 17598
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14476 15910 14504 16390
rect 14464 15904 14516 15910
rect 14462 15872 14464 15881
rect 14516 15872 14518 15881
rect 14462 15807 14518 15816
rect 14568 15722 14596 17546
rect 14660 17270 14688 17847
rect 14740 17818 14792 17824
rect 14844 17728 14872 20810
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15304 20398 15332 21082
rect 15396 20913 15424 21286
rect 15382 20904 15438 20913
rect 15382 20839 15438 20848
rect 15292 20392 15344 20398
rect 15344 20352 15424 20380
rect 15292 20334 15344 20340
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 14936 20058 14964 20266
rect 15290 20224 15346 20233
rect 15290 20159 15346 20168
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 15014 19000 15070 19009
rect 15014 18935 15016 18944
rect 15068 18935 15070 18944
rect 15016 18906 15068 18912
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15108 18080 15160 18086
rect 15108 18022 15160 18028
rect 15120 17898 15148 18022
rect 15120 17870 15240 17898
rect 15212 17814 15240 17870
rect 15200 17808 15252 17814
rect 15200 17750 15252 17756
rect 14752 17700 14872 17728
rect 15108 17740 15160 17746
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14476 15694 14596 15722
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14476 13841 14504 15694
rect 14646 15192 14702 15201
rect 14646 15127 14648 15136
rect 14700 15127 14702 15136
rect 14648 15098 14700 15104
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14462 13832 14518 13841
rect 14462 13767 14518 13776
rect 14280 13388 14332 13394
rect 14280 13330 14332 13336
rect 14292 12850 14320 13330
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14372 12708 14424 12714
rect 14372 12650 14424 12656
rect 14280 12436 14332 12442
rect 14280 12378 14332 12384
rect 14292 11354 14320 12378
rect 14384 12102 14412 12650
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10130 14320 10950
rect 14384 10674 14412 12038
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14292 9654 14320 10066
rect 14384 9994 14412 10610
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 3422 368 3478 377
rect 3422 303 3478 312
rect 8298 0 8354 480
rect 13910 0 13966 480
rect 14476 105 14504 13767
rect 14568 12442 14596 14010
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14568 11898 14596 12242
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14554 11792 14610 11801
rect 14554 11727 14556 11736
rect 14608 11727 14610 11736
rect 14556 11698 14608 11704
rect 14660 10742 14688 15098
rect 14752 13734 14780 17700
rect 15108 17682 15160 17688
rect 15120 17649 15148 17682
rect 14922 17640 14978 17649
rect 14844 17598 14922 17626
rect 14844 17202 14872 17598
rect 14922 17575 14924 17584
rect 14976 17575 14978 17584
rect 15106 17640 15162 17649
rect 15106 17575 15162 17584
rect 14924 17546 14976 17552
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14922 17232 14978 17241
rect 14832 17196 14884 17202
rect 14922 17167 14978 17176
rect 14832 17138 14884 17144
rect 14936 17066 14964 17167
rect 14924 17060 14976 17066
rect 14924 17002 14976 17008
rect 14936 16794 14964 17002
rect 14924 16788 14976 16794
rect 14924 16730 14976 16736
rect 14832 16720 14884 16726
rect 14832 16662 14884 16668
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13530 14780 13670
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14752 10810 14780 13466
rect 14844 13433 14872 16662
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 14890 15332 20159
rect 15396 19922 15424 20352
rect 15384 19916 15436 19922
rect 15384 19858 15436 19864
rect 15396 18222 15424 19858
rect 15488 19145 15516 21286
rect 15474 19136 15530 19145
rect 15474 19071 15530 19080
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15396 17746 15424 18158
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15476 16720 15528 16726
rect 15474 16688 15476 16697
rect 15528 16688 15530 16697
rect 15474 16623 15530 16632
rect 15382 16552 15438 16561
rect 15382 16487 15438 16496
rect 15292 14884 15344 14890
rect 15292 14826 15344 14832
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14830 13424 14886 13433
rect 15304 13394 15332 14350
rect 14830 13359 14886 13368
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15396 13274 15424 16487
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13938 15516 14214
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15304 13246 15424 13274
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12442 15332 13246
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 14844 11626 14872 12106
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 15212 11354 15240 11698
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 15304 10266 15332 11494
rect 15396 10538 15424 12922
rect 15488 12646 15516 13398
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12442 15516 12582
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15488 11150 15516 12378
rect 15580 12374 15608 24006
rect 15658 23896 15714 23905
rect 15658 23831 15714 23840
rect 15672 23594 15700 23831
rect 15660 23588 15712 23594
rect 15660 23530 15712 23536
rect 15660 23180 15712 23186
rect 15660 23122 15712 23128
rect 15672 22778 15700 23122
rect 15660 22772 15712 22778
rect 15660 22714 15712 22720
rect 15752 22500 15804 22506
rect 15752 22442 15804 22448
rect 15764 22137 15792 22442
rect 15750 22128 15806 22137
rect 15660 22092 15712 22098
rect 15750 22063 15806 22072
rect 15660 22034 15712 22040
rect 15672 21146 15700 22034
rect 15660 21140 15712 21146
rect 15660 21082 15712 21088
rect 15750 20632 15806 20641
rect 15660 20596 15712 20602
rect 15750 20567 15806 20576
rect 15660 20538 15712 20544
rect 15672 19990 15700 20538
rect 15660 19984 15712 19990
rect 15660 19926 15712 19932
rect 15672 19514 15700 19926
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15764 19446 15792 20567
rect 15752 19440 15804 19446
rect 15658 19408 15714 19417
rect 15752 19382 15804 19388
rect 15658 19343 15714 19352
rect 15672 18902 15700 19343
rect 15660 18896 15712 18902
rect 15660 18838 15712 18844
rect 15856 18426 15884 24550
rect 15948 22030 15976 25162
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 22953 16160 24550
rect 16224 24070 16252 25230
rect 16408 24682 16436 25298
rect 16764 25220 16816 25226
rect 16764 25162 16816 25168
rect 16776 24818 16804 25162
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 16764 24812 16816 24818
rect 16764 24754 16816 24760
rect 16396 24676 16448 24682
rect 16396 24618 16448 24624
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 16316 24070 16344 24550
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16316 23497 16344 24006
rect 16302 23488 16358 23497
rect 16302 23423 16358 23432
rect 16118 22944 16174 22953
rect 16118 22879 16174 22888
rect 16302 22672 16358 22681
rect 16302 22607 16358 22616
rect 16026 22536 16082 22545
rect 16026 22471 16082 22480
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 15948 21690 15976 21966
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15934 21448 15990 21457
rect 15934 21383 15936 21392
rect 15988 21383 15990 21392
rect 15936 21354 15988 21360
rect 16040 19310 16068 22471
rect 16120 21888 16172 21894
rect 16120 21830 16172 21836
rect 16132 21593 16160 21830
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16118 21584 16174 21593
rect 16118 21519 16120 21528
rect 16172 21519 16174 21528
rect 16120 21490 16172 21496
rect 16224 20330 16252 21626
rect 16316 20806 16344 22607
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16212 20324 16264 20330
rect 16212 20266 16264 20272
rect 16224 19378 16252 20266
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15856 16590 15884 18022
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15948 17338 15976 17750
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16316 16794 16344 16934
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15856 16250 15884 16526
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15672 12986 15700 14962
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15844 14476 15896 14482
rect 15844 14418 15896 14424
rect 15856 14074 15884 14418
rect 15844 14068 15896 14074
rect 15844 14010 15896 14016
rect 15948 13190 15976 14894
rect 16132 14822 16160 15302
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15580 12073 15608 12310
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15566 12064 15622 12073
rect 15566 11999 15622 12008
rect 15764 11354 15792 12242
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15856 11286 15884 12174
rect 16040 11762 16068 13942
rect 16132 13394 16160 14758
rect 16316 14278 16344 15506
rect 16304 14272 16356 14278
rect 16304 14214 16356 14220
rect 16120 13388 16172 13394
rect 16172 13348 16252 13376
rect 16120 13330 16172 13336
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15672 10810 15700 11154
rect 16040 11150 16068 11698
rect 16224 11370 16252 13348
rect 16316 12238 16344 14214
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11898 16344 12038
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16224 11342 16344 11370
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 10810 16068 11086
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15672 9722 15700 10746
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15764 8945 15792 10406
rect 16132 10266 16160 11018
rect 16224 10674 16252 11222
rect 16316 11082 16344 11342
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16408 10849 16436 24618
rect 16762 24440 16818 24449
rect 16762 24375 16818 24384
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16592 23254 16620 24142
rect 16684 23866 16712 24210
rect 16672 23860 16724 23866
rect 16672 23802 16724 23808
rect 16684 23730 16712 23802
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 16684 23322 16712 23666
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 16592 22574 16620 23190
rect 16580 22568 16632 22574
rect 16580 22510 16632 22516
rect 16592 22234 16620 22510
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16500 20890 16528 20946
rect 16500 20862 16712 20890
rect 16684 20602 16712 20862
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16486 20088 16542 20097
rect 16684 20058 16712 20538
rect 16486 20023 16542 20032
rect 16672 20052 16724 20058
rect 16500 18873 16528 20023
rect 16672 19994 16724 20000
rect 16486 18864 16542 18873
rect 16486 18799 16542 18808
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17898 16528 18022
rect 16500 17882 16620 17898
rect 16500 17876 16632 17882
rect 16500 17870 16580 17876
rect 16580 17818 16632 17824
rect 16486 16552 16542 16561
rect 16486 16487 16542 16496
rect 16500 16250 16528 16487
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16670 16416 16726 16425
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16592 16046 16620 16390
rect 16670 16351 16726 16360
rect 16580 16040 16632 16046
rect 16684 16017 16712 16351
rect 16580 15982 16632 15988
rect 16670 16008 16726 16017
rect 16592 15473 16620 15982
rect 16670 15943 16726 15952
rect 16578 15464 16634 15473
rect 16578 15399 16634 15408
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 14958 16528 15302
rect 16776 14958 16804 24375
rect 17052 23866 17080 25094
rect 17512 24154 17540 25871
rect 17604 24857 17632 27520
rect 17868 25356 17920 25362
rect 17788 25316 17868 25344
rect 17590 24848 17646 24857
rect 17590 24783 17646 24792
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17696 24342 17724 24686
rect 17788 24614 17816 25316
rect 17868 25298 17920 25304
rect 18156 24834 18184 27520
rect 18604 25220 18656 25226
rect 18604 25162 18656 25168
rect 18156 24806 18276 24834
rect 18616 24818 18644 25162
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24336 17736 24342
rect 17684 24278 17736 24284
rect 17512 24126 17724 24154
rect 17498 24032 17554 24041
rect 17498 23967 17554 23976
rect 17512 23866 17540 23967
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17052 23594 17080 23802
rect 17040 23588 17092 23594
rect 17040 23530 17092 23536
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16868 22710 16896 23122
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17408 22500 17460 22506
rect 17408 22442 17460 22448
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17144 21146 17172 22034
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17132 21140 17184 21146
rect 17132 21082 17184 21088
rect 17052 21049 17080 21082
rect 17038 21040 17094 21049
rect 17038 20975 17094 20984
rect 16854 19952 16910 19961
rect 16854 19887 16910 19896
rect 16868 19514 16896 19887
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16868 18426 16896 19314
rect 17132 19168 17184 19174
rect 17132 19110 17184 19116
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 17144 18057 17172 19110
rect 17328 18057 17356 21966
rect 17420 21321 17448 22442
rect 17406 21312 17462 21321
rect 17406 21247 17462 21256
rect 17498 21176 17554 21185
rect 17498 21111 17554 21120
rect 17512 20534 17540 21111
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17604 20346 17632 22578
rect 17696 22030 17724 24126
rect 17788 22409 17816 24550
rect 17774 22400 17830 22409
rect 17774 22335 17830 22344
rect 17880 22098 17908 24550
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17972 23594 18000 24006
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 23588 18012 23594
rect 17960 23530 18012 23536
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17972 22234 18000 23122
rect 18064 22982 18092 23598
rect 18144 23112 18196 23118
rect 18142 23080 18144 23089
rect 18196 23080 18198 23089
rect 18142 23015 18198 23024
rect 18052 22976 18104 22982
rect 18052 22918 18104 22924
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17696 21622 17724 21966
rect 17684 21616 17736 21622
rect 17684 21558 17736 21564
rect 18064 21486 18092 22918
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17604 20318 17724 20346
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 19922 17632 20198
rect 17592 19916 17644 19922
rect 17592 19858 17644 19864
rect 17604 19718 17632 19858
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17512 18426 17540 18770
rect 17500 18420 17552 18426
rect 17500 18362 17552 18368
rect 17130 18048 17186 18057
rect 17130 17983 17186 17992
rect 17314 18048 17370 18057
rect 17314 17983 17370 17992
rect 17038 17776 17094 17785
rect 17038 17711 17040 17720
rect 17092 17711 17094 17720
rect 17040 17682 17092 17688
rect 17052 16658 17080 17682
rect 17132 17060 17184 17066
rect 17132 17002 17184 17008
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16854 16008 16910 16017
rect 16854 15943 16856 15952
rect 16908 15943 16910 15952
rect 16856 15914 16908 15920
rect 16854 15872 16910 15881
rect 16854 15807 16910 15816
rect 16488 14952 16540 14958
rect 16488 14894 16540 14900
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16500 13512 16528 13942
rect 16684 13938 16712 14758
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16580 13524 16632 13530
rect 16500 13484 16580 13512
rect 16580 13466 16632 13472
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12374 16620 12582
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16776 12238 16804 12378
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 11762 16804 12174
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16500 11665 16528 11698
rect 16486 11656 16542 11665
rect 16486 11591 16542 11600
rect 16776 11286 16804 11698
rect 16868 11354 16896 15807
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 12850 16988 14758
rect 17052 14346 17080 14962
rect 17040 14340 17092 14346
rect 17040 14282 17092 14288
rect 17052 13462 17080 14282
rect 17040 13456 17092 13462
rect 17040 13398 17092 13404
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11558 17080 12242
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16394 10840 16450 10849
rect 16394 10775 16450 10784
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16224 10198 16252 10610
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 15750 8936 15806 8945
rect 15750 8871 15806 8880
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 16408 7993 16436 10775
rect 16500 9654 16528 11018
rect 16868 10470 16896 11154
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16394 7984 16450 7993
rect 16394 7919 16450 7928
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 16868 7449 16896 10406
rect 16854 7440 16910 7449
rect 16854 7375 16910 7384
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 17052 4049 17080 11494
rect 17144 9625 17172 17002
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17512 16114 17540 16662
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17328 14929 17356 15030
rect 17314 14920 17370 14929
rect 17314 14855 17370 14864
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17236 13530 17264 13738
rect 17224 13524 17276 13530
rect 17224 13466 17276 13472
rect 17314 12472 17370 12481
rect 17314 12407 17370 12416
rect 17328 12306 17356 12407
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17314 11248 17370 11257
rect 17420 11234 17448 15982
rect 17512 15910 17540 16050
rect 17500 15904 17552 15910
rect 17500 15846 17552 15852
rect 17512 15434 17540 15846
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17604 15366 17632 19654
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17696 13705 17724 20318
rect 17868 19780 17920 19786
rect 17868 19722 17920 19728
rect 17880 19258 17908 19722
rect 17880 19230 18000 19258
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17788 19009 17816 19110
rect 17774 19000 17830 19009
rect 17774 18935 17830 18944
rect 17972 18902 18000 19230
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18064 18290 18092 19110
rect 18156 18970 18184 21558
rect 18248 19417 18276 24806
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18510 24712 18566 24721
rect 18510 24647 18566 24656
rect 18420 24404 18472 24410
rect 18420 24346 18472 24352
rect 18326 24032 18382 24041
rect 18326 23967 18382 23976
rect 18340 21962 18368 23967
rect 18432 22710 18460 24346
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18328 21956 18380 21962
rect 18328 21898 18380 21904
rect 18328 21480 18380 21486
rect 18328 21422 18380 21428
rect 18418 21448 18474 21457
rect 18340 20874 18368 21422
rect 18418 21383 18474 21392
rect 18432 21350 18460 21383
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18418 21176 18474 21185
rect 18418 21111 18474 21120
rect 18432 21010 18460 21111
rect 18420 21004 18472 21010
rect 18420 20946 18472 20952
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18340 20262 18368 20810
rect 18328 20256 18380 20262
rect 18524 20233 18552 24647
rect 18616 21146 18644 24754
rect 18708 22522 18736 27520
rect 19156 25356 19208 25362
rect 19156 25298 19208 25304
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18788 24948 18840 24954
rect 18788 24890 18840 24896
rect 18800 23168 18828 24890
rect 18892 24410 18920 25230
rect 18972 25220 19024 25226
rect 18972 25162 19024 25168
rect 18984 24750 19012 25162
rect 18972 24744 19024 24750
rect 19168 24721 19196 25298
rect 18972 24686 19024 24692
rect 19154 24712 19210 24721
rect 19154 24647 19156 24656
rect 19208 24647 19210 24656
rect 19156 24618 19208 24624
rect 18972 24608 19024 24614
rect 19260 24585 19288 27520
rect 19812 25786 19840 27520
rect 19812 25758 20024 25786
rect 20364 25770 20392 27520
rect 20916 25838 20944 27520
rect 20904 25832 20956 25838
rect 20534 25800 20590 25809
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19338 24848 19394 24857
rect 19522 24848 19578 24857
rect 19338 24783 19394 24792
rect 19444 24806 19522 24834
rect 18972 24550 19024 24556
rect 19246 24576 19302 24585
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18984 24206 19012 24550
rect 19246 24511 19302 24520
rect 18972 24200 19024 24206
rect 18970 24168 18972 24177
rect 19024 24168 19026 24177
rect 18970 24103 19026 24112
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 18800 23140 18920 23168
rect 18786 23080 18842 23089
rect 18786 23015 18842 23024
rect 18800 22642 18828 23015
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18708 22494 18828 22522
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18708 20602 18736 20878
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18328 20198 18380 20204
rect 18510 20224 18566 20233
rect 18340 19922 18368 20198
rect 18510 20159 18566 20168
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 18234 19408 18290 19417
rect 18234 19343 18290 19352
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 18156 18426 18184 18906
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18340 18306 18368 19858
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18510 19272 18566 19281
rect 18432 18737 18460 19246
rect 18510 19207 18512 19216
rect 18564 19207 18566 19216
rect 18512 19178 18564 19184
rect 18616 18766 18644 19314
rect 18604 18760 18656 18766
rect 18418 18728 18474 18737
rect 18604 18702 18656 18708
rect 18418 18663 18474 18672
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18052 18284 18104 18290
rect 18052 18226 18104 18232
rect 18156 18278 18368 18306
rect 18064 18170 18092 18226
rect 17880 18142 18092 18170
rect 17880 17814 17908 18142
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17882 18092 18022
rect 18052 17876 18104 17882
rect 18052 17818 18104 17824
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17774 17640 17830 17649
rect 17774 17575 17776 17584
rect 17828 17575 17830 17584
rect 17776 17546 17828 17552
rect 18064 16998 18092 17682
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16794 18092 16934
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18052 16040 18104 16046
rect 18156 16028 18184 18278
rect 18432 18222 18460 18566
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18524 17814 18552 18634
rect 18800 18465 18828 22494
rect 18786 18456 18842 18465
rect 18786 18391 18842 18400
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18708 17882 18736 18226
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18340 17338 18368 17614
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18236 17060 18288 17066
rect 18236 17002 18288 17008
rect 18104 16000 18184 16028
rect 18052 15982 18104 15988
rect 18248 15706 18276 17002
rect 18340 16250 18368 17274
rect 18708 17202 18736 17818
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18524 16561 18552 16934
rect 18510 16552 18566 16561
rect 18708 16522 18736 17138
rect 18510 16487 18566 16496
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18340 15638 18368 16186
rect 18708 16046 18736 16458
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17788 15366 17816 15399
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17866 15192 17922 15201
rect 17866 15127 17868 15136
rect 17920 15127 17922 15136
rect 17868 15098 17920 15104
rect 17972 14890 18000 15506
rect 18340 14958 18368 15574
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18708 15201 18736 15438
rect 18694 15192 18750 15201
rect 18694 15127 18750 15136
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 18064 14226 18092 14894
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 17972 14198 18092 14226
rect 17972 13870 18000 14198
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17682 13696 17738 13705
rect 17682 13631 17738 13640
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 12986 17816 13398
rect 17972 13326 18000 13806
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17880 12782 17908 13126
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17604 11558 17632 12242
rect 17972 11626 18000 13262
rect 18156 12986 18184 14418
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18248 14074 18276 14350
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18432 14006 18460 14350
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18800 13870 18828 14214
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 12442 18460 12718
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18432 11898 18460 12242
rect 18800 11937 18828 12378
rect 18786 11928 18842 11937
rect 18420 11892 18472 11898
rect 18786 11863 18842 11872
rect 18420 11834 18472 11840
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17420 11206 17540 11234
rect 17314 11183 17370 11192
rect 17328 11150 17356 11183
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10470 17356 11086
rect 17316 10464 17368 10470
rect 17316 10406 17368 10412
rect 17130 9616 17186 9625
rect 17130 9551 17186 9560
rect 17038 4040 17094 4049
rect 17038 3975 17094 3984
rect 17328 3641 17356 10406
rect 17512 6361 17540 11206
rect 17604 11121 17632 11494
rect 17684 11144 17736 11150
rect 17590 11112 17646 11121
rect 17684 11086 17736 11092
rect 17590 11047 17646 11056
rect 17696 10810 17724 11086
rect 17972 11082 18000 11562
rect 18800 11558 18828 11863
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11218 18828 11494
rect 18892 11354 18920 23140
rect 18984 22982 19012 23530
rect 19076 23186 19104 24006
rect 19246 23624 19302 23633
rect 19246 23559 19302 23568
rect 19064 23180 19116 23186
rect 19064 23122 19116 23128
rect 19156 23044 19208 23050
rect 19156 22986 19208 22992
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18984 22642 19012 22918
rect 19168 22778 19196 22986
rect 19260 22982 19288 23559
rect 19248 22976 19300 22982
rect 19248 22918 19300 22924
rect 19156 22772 19208 22778
rect 19156 22714 19208 22720
rect 18972 22636 19024 22642
rect 18972 22578 19024 22584
rect 18984 22030 19012 22578
rect 19154 22128 19210 22137
rect 19064 22092 19116 22098
rect 19154 22063 19210 22072
rect 19064 22034 19116 22040
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18984 21690 19012 21966
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 19076 21350 19104 22034
rect 19168 21690 19196 22063
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 18984 20398 19012 21082
rect 18972 20392 19024 20398
rect 18972 20334 19024 20340
rect 18984 20058 19012 20334
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18984 18086 19012 18566
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 15502 19012 18022
rect 19076 16946 19104 21286
rect 19352 21146 19380 24783
rect 19444 24449 19472 24806
rect 19522 24783 19578 24792
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19430 24440 19486 24449
rect 19430 24375 19486 24384
rect 19536 24313 19564 24550
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19522 24304 19578 24313
rect 19432 24268 19484 24274
rect 19522 24239 19578 24248
rect 19432 24210 19484 24216
rect 19444 23050 19472 24210
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19536 24041 19564 24142
rect 19522 24032 19578 24041
rect 19522 23967 19578 23976
rect 19628 23866 19656 24142
rect 19616 23860 19668 23866
rect 19536 23820 19616 23848
rect 19536 23322 19564 23820
rect 19616 23802 19668 23808
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19432 23044 19484 23050
rect 19432 22986 19484 22992
rect 19430 22672 19486 22681
rect 19536 22642 19564 23258
rect 19616 23180 19668 23186
rect 19616 23122 19668 23128
rect 19628 22778 19656 23122
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19430 22607 19486 22616
rect 19524 22636 19576 22642
rect 19444 22574 19472 22607
rect 19524 22578 19576 22584
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 19628 22488 19656 22714
rect 19720 22681 19748 23054
rect 19706 22672 19762 22681
rect 19706 22607 19762 22616
rect 19800 22568 19852 22574
rect 19904 22556 19932 23054
rect 19852 22528 19932 22556
rect 19800 22510 19852 22516
rect 19536 22460 19656 22488
rect 19432 21888 19484 21894
rect 19430 21856 19432 21865
rect 19484 21856 19486 21865
rect 19430 21791 19486 21800
rect 19444 21486 19472 21791
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19168 19825 19196 19926
rect 19154 19816 19210 19825
rect 19154 19751 19210 19760
rect 19168 19514 19196 19751
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19260 19258 19288 20742
rect 19444 20602 19472 21422
rect 19536 20641 19564 22460
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19522 20632 19578 20641
rect 19432 20596 19484 20602
rect 19522 20567 19578 20576
rect 19432 20538 19484 20544
rect 19338 20360 19394 20369
rect 19338 20295 19394 20304
rect 19352 19514 19380 20295
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19706 19408 19762 19417
rect 19706 19343 19762 19352
rect 19260 19230 19380 19258
rect 19720 19242 19748 19343
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19156 18828 19208 18834
rect 19156 18770 19208 18776
rect 19168 18086 19196 18770
rect 19260 18630 19288 18838
rect 19352 18834 19380 19230
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19260 17785 19288 18566
rect 19444 18329 19472 18702
rect 19430 18320 19486 18329
rect 19430 18255 19486 18264
rect 19338 18048 19394 18057
rect 19338 17983 19394 17992
rect 19246 17776 19302 17785
rect 19246 17711 19302 17720
rect 19076 16918 19196 16946
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18984 14618 19012 15438
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19076 13258 19104 13806
rect 19064 13252 19116 13258
rect 19064 13194 19116 13200
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18984 12238 19012 12854
rect 19076 12850 19104 13194
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19076 12374 19104 12786
rect 19168 12753 19196 16918
rect 19352 16658 19380 17983
rect 19536 17814 19564 19110
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19524 17808 19576 17814
rect 19524 17750 19576 17756
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19444 16794 19472 17682
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16794 20024 25758
rect 20352 25764 20404 25770
rect 20904 25774 20956 25780
rect 20534 25735 20590 25744
rect 20352 25706 20404 25712
rect 20444 25356 20496 25362
rect 20444 25298 20496 25304
rect 20076 25152 20128 25158
rect 20076 25094 20128 25100
rect 20088 24614 20116 25094
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 23497 20116 24550
rect 20180 24410 20208 24618
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20166 24304 20222 24313
rect 20166 24239 20222 24248
rect 20074 23488 20130 23497
rect 20074 23423 20130 23432
rect 20076 22568 20128 22574
rect 20076 22510 20128 22516
rect 20088 22234 20116 22510
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 20180 22114 20208 24239
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20272 22234 20300 23122
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20364 22137 20392 24754
rect 20456 24070 20484 25298
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20088 22086 20208 22114
rect 20350 22128 20406 22137
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20088 16674 20116 22086
rect 20350 22063 20406 22072
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20168 21004 20220 21010
rect 20168 20946 20220 20952
rect 20180 19718 20208 20946
rect 20272 20874 20300 21830
rect 20456 21570 20484 24006
rect 20364 21542 20484 21570
rect 20260 20868 20312 20874
rect 20260 20810 20312 20816
rect 20168 19712 20220 19718
rect 20364 19689 20392 21542
rect 20548 21457 20576 25735
rect 21560 25514 21588 27520
rect 21468 25486 21588 25514
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21088 25152 21140 25158
rect 21088 25094 21140 25100
rect 21100 24886 21128 25094
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20732 23798 20760 24210
rect 20720 23792 20772 23798
rect 20718 23760 20720 23769
rect 20772 23760 20774 23769
rect 20718 23695 20774 23704
rect 20916 23662 20944 24822
rect 20996 24812 21048 24818
rect 20996 24754 21048 24760
rect 21008 24614 21036 24754
rect 21192 24750 21220 25230
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 20996 24608 21048 24614
rect 20996 24550 21048 24556
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20904 23112 20956 23118
rect 20904 23054 20956 23060
rect 20718 22944 20774 22953
rect 20718 22879 20774 22888
rect 20534 21448 20590 21457
rect 20456 21406 20534 21434
rect 20168 19654 20220 19660
rect 20350 19680 20406 19689
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19536 16646 20116 16674
rect 19352 16182 19380 16594
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19352 14464 19380 15302
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19260 14436 19380 14464
rect 19260 14278 19288 14436
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19352 13530 19380 14282
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19444 12918 19472 14758
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19432 12776 19484 12782
rect 19154 12744 19210 12753
rect 19432 12718 19484 12724
rect 19154 12679 19210 12688
rect 19444 12646 19472 12718
rect 19432 12640 19484 12646
rect 19430 12608 19432 12617
rect 19484 12608 19486 12617
rect 19430 12543 19486 12552
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18984 11286 19012 12174
rect 19536 11762 19564 16646
rect 19982 16008 20038 16017
rect 19982 15943 20038 15952
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17696 10130 17724 10746
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19996 8566 20024 15943
rect 20180 14550 20208 19654
rect 20350 19615 20406 19624
rect 20456 18086 20484 21406
rect 20534 21383 20590 21392
rect 20732 21146 20760 22879
rect 20916 21894 20944 23054
rect 21008 22098 21036 24550
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 21008 21350 21036 22034
rect 20996 21344 21048 21350
rect 20996 21286 21048 21292
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20732 21010 20760 21082
rect 20720 21004 20772 21010
rect 20720 20946 20772 20952
rect 21100 20942 21128 23598
rect 21192 21434 21220 24686
rect 21364 24608 21416 24614
rect 21364 24550 21416 24556
rect 21376 24313 21404 24550
rect 21362 24304 21418 24313
rect 21362 24239 21418 24248
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21284 23662 21312 24074
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21272 23656 21324 23662
rect 21376 23633 21404 24006
rect 21468 23905 21496 25486
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21560 24954 21588 25298
rect 21548 24948 21600 24954
rect 21548 24890 21600 24896
rect 21916 24880 21968 24886
rect 21916 24822 21968 24828
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 21454 23896 21510 23905
rect 21454 23831 21510 23840
rect 21272 23598 21324 23604
rect 21362 23624 21418 23633
rect 21362 23559 21364 23568
rect 21416 23559 21418 23568
rect 21364 23530 21416 23536
rect 21652 23254 21680 24142
rect 21836 24041 21864 24278
rect 21822 24032 21878 24041
rect 21822 23967 21878 23976
rect 21836 23866 21864 23967
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21928 23254 21956 24822
rect 22112 24818 22140 27520
rect 22664 24857 22692 27520
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 22282 24848 22338 24857
rect 22100 24812 22152 24818
rect 22282 24783 22338 24792
rect 22650 24848 22706 24857
rect 22650 24783 22706 24792
rect 22744 24812 22796 24818
rect 22100 24754 22152 24760
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22020 23338 22048 23666
rect 22020 23322 22140 23338
rect 22020 23316 22152 23322
rect 22020 23310 22100 23316
rect 22100 23258 22152 23264
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21916 23248 21968 23254
rect 21916 23190 21968 23196
rect 21652 22778 21680 23190
rect 21640 22772 21692 22778
rect 21640 22714 21692 22720
rect 21270 22128 21326 22137
rect 21270 22063 21326 22072
rect 21284 21962 21312 22063
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21928 21865 21956 23190
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 22112 22114 22140 22374
rect 22020 22086 22140 22114
rect 21914 21856 21970 21865
rect 21914 21791 21970 21800
rect 22020 21690 22048 22086
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 21192 21406 21312 21434
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20904 20868 20956 20874
rect 20904 20810 20956 20816
rect 20718 20496 20774 20505
rect 20718 20431 20774 20440
rect 20732 20398 20760 20431
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 20824 19922 20852 20810
rect 20916 20262 20944 20810
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20916 19961 20944 20198
rect 20902 19952 20958 19961
rect 20812 19916 20864 19922
rect 20902 19887 20958 19896
rect 20812 19858 20864 19864
rect 20824 19378 20852 19858
rect 20812 19372 20864 19378
rect 20812 19314 20864 19320
rect 20824 18970 20852 19314
rect 20812 18964 20864 18970
rect 20812 18906 20864 18912
rect 21008 18850 21036 20198
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 20824 18822 21036 18850
rect 20732 18426 20760 18770
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20548 17542 20576 18226
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16590 20484 17070
rect 20548 17066 20576 17478
rect 20536 17060 20588 17066
rect 20536 17002 20588 17008
rect 20548 16658 20576 17002
rect 20720 16720 20772 16726
rect 20824 16697 20852 18822
rect 20994 18728 21050 18737
rect 20994 18663 21050 18672
rect 21008 18426 21036 18663
rect 20996 18420 21048 18426
rect 20996 18362 21048 18368
rect 21008 18222 21036 18362
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 20996 17672 21048 17678
rect 20916 17620 20996 17626
rect 20916 17614 21048 17620
rect 20916 17598 21036 17614
rect 20916 16998 20944 17598
rect 21100 17338 21128 17682
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20916 16794 20944 16934
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20720 16662 20772 16668
rect 20810 16688 20866 16697
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20444 16584 20496 16590
rect 20444 16526 20496 16532
rect 20258 16008 20314 16017
rect 20258 15943 20314 15952
rect 20272 15609 20300 15943
rect 20258 15600 20314 15609
rect 20258 15535 20314 15544
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15162 20392 15438
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20364 14958 20392 15098
rect 20548 15026 20576 16594
rect 20732 16250 20760 16662
rect 20810 16623 20866 16632
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20720 16040 20772 16046
rect 20824 16028 20852 16526
rect 20916 16250 20944 16730
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20902 16144 20958 16153
rect 20902 16079 20958 16088
rect 20772 16000 20852 16028
rect 20720 15982 20772 15988
rect 20732 15366 20760 15982
rect 20916 15688 20944 16079
rect 21100 15706 21128 17274
rect 20824 15660 20944 15688
rect 21088 15700 21140 15706
rect 20720 15360 20772 15366
rect 20626 15328 20682 15337
rect 20720 15302 20772 15308
rect 20626 15263 20682 15272
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 14074 20300 14418
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20640 12918 20668 15263
rect 20732 14414 20760 15302
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 13530 20760 14350
rect 20824 14074 20852 15660
rect 21088 15642 21140 15648
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20916 15162 20944 15506
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20824 12986 20852 13262
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12102 20116 12582
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20088 8265 20116 12038
rect 20074 8256 20130 8265
rect 19622 8188 19918 8208
rect 20074 8191 20130 8200
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 20180 7041 20208 12718
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20916 11354 20944 12038
rect 20904 11348 20956 11354
rect 20904 11290 20956 11296
rect 21008 10849 21036 14758
rect 20994 10840 21050 10849
rect 20994 10775 21050 10784
rect 21192 10577 21220 21286
rect 21284 20262 21312 21406
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21376 20058 21404 20878
rect 21638 20632 21694 20641
rect 21638 20567 21694 20576
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21284 19174 21312 19858
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 13954 21312 19110
rect 21560 19009 21588 19178
rect 21546 19000 21602 19009
rect 21546 18935 21602 18944
rect 21548 18828 21600 18834
rect 21548 18770 21600 18776
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21376 17814 21404 18566
rect 21468 18426 21496 18702
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21560 18086 21588 18770
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21560 17882 21588 18022
rect 21548 17876 21600 17882
rect 21548 17818 21600 17824
rect 21364 17808 21416 17814
rect 21364 17750 21416 17756
rect 21376 17338 21404 17750
rect 21652 17649 21680 20567
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 21730 19136 21786 19145
rect 21730 19071 21786 19080
rect 21638 17640 21694 17649
rect 21638 17575 21694 17584
rect 21364 17332 21416 17338
rect 21364 17274 21416 17280
rect 21364 15496 21416 15502
rect 21364 15438 21416 15444
rect 21376 14550 21404 15438
rect 21454 15192 21510 15201
rect 21454 15127 21510 15136
rect 21364 14544 21416 14550
rect 21364 14486 21416 14492
rect 21376 14074 21404 14486
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21284 13926 21404 13954
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21284 12986 21312 13330
rect 21376 13326 21404 13926
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21284 12442 21312 12922
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 21284 11898 21312 12135
rect 21376 12102 21404 12582
rect 21468 12306 21496 15127
rect 21546 14512 21602 14521
rect 21546 14447 21602 14456
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21364 12096 21416 12102
rect 21364 12038 21416 12044
rect 21560 11898 21588 14447
rect 21640 13728 21692 13734
rect 21640 13670 21692 13676
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21284 11694 21312 11834
rect 21272 11688 21324 11694
rect 21272 11630 21324 11636
rect 21652 10713 21680 13670
rect 21744 12442 21772 19071
rect 21914 19000 21970 19009
rect 21914 18935 21970 18944
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 21836 17270 21864 18362
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21836 16726 21864 17206
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21836 15502 21864 16662
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15162 21864 15438
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21928 14770 21956 18935
rect 22020 15337 22048 20198
rect 22098 18592 22154 18601
rect 22098 18527 22154 18536
rect 22006 15328 22062 15337
rect 22006 15263 22062 15272
rect 22112 15162 22140 18527
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21928 14742 22048 14770
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21928 13938 21956 14554
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 21836 12714 21864 13806
rect 21928 13530 21956 13874
rect 22020 13705 22048 14742
rect 22112 14618 22140 14962
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22006 13696 22062 13705
rect 22006 13631 22062 13640
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21914 13424 21970 13433
rect 21914 13359 21970 13368
rect 21824 12708 21876 12714
rect 21824 12650 21876 12656
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21836 11898 21864 12242
rect 21824 11892 21876 11898
rect 21824 11834 21876 11840
rect 21928 11218 21956 13359
rect 22020 12850 22048 13631
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21928 10810 21956 11154
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 21638 10704 21694 10713
rect 21638 10639 21694 10648
rect 21178 10568 21234 10577
rect 21178 10503 21234 10512
rect 20442 8392 20498 8401
rect 20442 8327 20498 8336
rect 20166 7032 20222 7041
rect 20166 6967 20222 6976
rect 17498 6352 17554 6361
rect 17498 6287 17554 6296
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 17314 3632 17370 3641
rect 17314 3567 17370 3576
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 18510 2408 18566 2417
rect 18510 2343 18512 2352
rect 18564 2343 18566 2352
rect 18512 2314 18564 2320
rect 19524 2304 19576 2310
rect 19524 2246 19576 2252
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 19536 480 19564 2246
rect 20456 1465 20484 8327
rect 22020 7449 22048 12650
rect 22112 11354 22140 14350
rect 22204 13530 22232 24686
rect 22296 24342 22324 24783
rect 22744 24754 22796 24760
rect 22466 24712 22522 24721
rect 22466 24647 22522 24656
rect 22284 24336 22336 24342
rect 22284 24278 22336 24284
rect 22296 23866 22324 24278
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22480 23662 22508 24647
rect 22650 24168 22706 24177
rect 22650 24103 22652 24112
rect 22704 24103 22706 24112
rect 22652 24074 22704 24080
rect 22468 23656 22520 23662
rect 22468 23598 22520 23604
rect 22376 23316 22428 23322
rect 22376 23258 22428 23264
rect 22388 22166 22416 23258
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21486 22324 21830
rect 22388 21622 22416 22102
rect 22376 21616 22428 21622
rect 22376 21558 22428 21564
rect 22284 21480 22336 21486
rect 22284 21422 22336 21428
rect 22284 20800 22336 20806
rect 22284 20742 22336 20748
rect 22296 20330 22324 20742
rect 22284 20324 22336 20330
rect 22284 20266 22336 20272
rect 22296 19281 22324 20266
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22282 19272 22338 19281
rect 22282 19207 22338 19216
rect 22296 18086 22324 19207
rect 22284 18080 22336 18086
rect 22282 18048 22284 18057
rect 22336 18048 22338 18057
rect 22282 17983 22338 17992
rect 22282 17776 22338 17785
rect 22282 17711 22338 17720
rect 22296 15706 22324 17711
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22296 14074 22324 14418
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22282 11928 22338 11937
rect 22282 11863 22284 11872
rect 22336 11863 22338 11872
rect 22284 11834 22336 11840
rect 22296 11694 22324 11834
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22388 9489 22416 20198
rect 22480 20058 22508 22918
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22560 22500 22612 22506
rect 22560 22442 22612 22448
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22480 19825 22508 19994
rect 22466 19816 22522 19825
rect 22466 19751 22522 19760
rect 22468 19236 22520 19242
rect 22468 19178 22520 19184
rect 22480 18970 22508 19178
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22572 18714 22600 22442
rect 22480 18686 22600 18714
rect 22480 16697 22508 18686
rect 22664 18578 22692 22714
rect 22572 18550 22692 18578
rect 22466 16688 22522 16697
rect 22466 16623 22522 16632
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22480 13394 22508 16050
rect 22572 15065 22600 18550
rect 22650 18456 22706 18465
rect 22650 18391 22706 18400
rect 22664 17882 22692 18391
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22664 15473 22692 15506
rect 22650 15464 22706 15473
rect 22650 15399 22706 15408
rect 22558 15056 22614 15065
rect 22558 14991 22614 15000
rect 22572 13818 22600 14991
rect 22664 14618 22692 15399
rect 22756 15162 22784 24754
rect 22834 24712 22890 24721
rect 22834 24647 22890 24656
rect 22848 23866 22876 24647
rect 22940 24426 22968 25638
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 23032 24614 23060 25230
rect 23216 24750 23244 27520
rect 23204 24744 23256 24750
rect 23204 24686 23256 24692
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 23204 24608 23256 24614
rect 23480 24608 23532 24614
rect 23204 24550 23256 24556
rect 23400 24556 23480 24562
rect 23400 24550 23532 24556
rect 22940 24398 23060 24426
rect 23032 24274 23060 24398
rect 23020 24268 23072 24274
rect 23020 24210 23072 24216
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 23032 23526 23060 24210
rect 23216 24206 23244 24550
rect 23400 24534 23520 24550
rect 23204 24200 23256 24206
rect 23204 24142 23256 24148
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23124 22778 23152 23122
rect 23216 22982 23244 24142
rect 23400 23225 23428 24534
rect 23768 24426 23796 27520
rect 24320 25430 24348 27520
rect 24766 26480 24822 26489
rect 24766 26415 24822 26424
rect 24674 25936 24730 25945
rect 24674 25871 24730 25880
rect 24308 25424 24360 25430
rect 24308 25366 24360 25372
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24688 24954 24716 25871
rect 24780 25378 24808 26415
rect 24872 25514 24900 27520
rect 25424 27418 25452 27520
rect 25332 27390 25452 27418
rect 25134 27160 25190 27169
rect 25134 27095 25190 27104
rect 24872 25486 24992 25514
rect 24780 25350 24900 25378
rect 24766 25256 24822 25265
rect 24766 25191 24768 25200
rect 24820 25191 24822 25200
rect 24768 25162 24820 25168
rect 24872 25106 24900 25350
rect 24780 25078 24900 25106
rect 24676 24948 24728 24954
rect 24676 24890 24728 24896
rect 23768 24398 24072 24426
rect 24780 24410 24808 25078
rect 24860 24608 24912 24614
rect 24860 24550 24912 24556
rect 23664 24064 23716 24070
rect 23664 24006 23716 24012
rect 23676 23798 23704 24006
rect 23664 23792 23716 23798
rect 23664 23734 23716 23740
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 23386 23216 23442 23225
rect 23386 23151 23442 23160
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23492 22794 23520 23530
rect 23848 23520 23900 23526
rect 23662 23488 23718 23497
rect 23900 23468 23980 23474
rect 23848 23462 23980 23468
rect 23860 23446 23980 23462
rect 23662 23423 23718 23432
rect 23676 23322 23704 23423
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23216 22766 23520 22794
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23124 20874 23152 21014
rect 23112 20868 23164 20874
rect 23112 20810 23164 20816
rect 23020 20256 23072 20262
rect 23018 20224 23020 20233
rect 23072 20224 23074 20233
rect 23018 20159 23074 20168
rect 22834 19816 22890 19825
rect 22834 19751 22890 19760
rect 22848 16114 22876 19751
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 22940 16833 22968 17682
rect 23032 17048 23060 20159
rect 23124 20058 23152 20810
rect 23112 20052 23164 20058
rect 23112 19994 23164 20000
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23124 18426 23152 18702
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23032 17020 23152 17048
rect 23018 16960 23074 16969
rect 23018 16895 23074 16904
rect 22926 16824 22982 16833
rect 22926 16759 22928 16768
rect 22980 16759 22982 16768
rect 22928 16730 22980 16736
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22836 15972 22888 15978
rect 22836 15914 22888 15920
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22652 14612 22704 14618
rect 22652 14554 22704 14560
rect 22756 13938 22784 14826
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22572 13790 22692 13818
rect 22468 13388 22520 13394
rect 22468 13330 22520 13336
rect 22558 12336 22614 12345
rect 22558 12271 22614 12280
rect 22572 11218 22600 12271
rect 22664 11393 22692 13790
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22756 12986 22784 13398
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22744 12436 22796 12442
rect 22744 12378 22796 12384
rect 22756 12345 22784 12378
rect 22742 12336 22798 12345
rect 22742 12271 22798 12280
rect 22742 12064 22798 12073
rect 22742 11999 22798 12008
rect 22650 11384 22706 11393
rect 22650 11319 22706 11328
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22572 10674 22600 10950
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22756 9586 22784 11999
rect 22848 10266 22876 15914
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22940 15638 22968 15846
rect 22928 15632 22980 15638
rect 22928 15574 22980 15580
rect 22940 15162 22968 15574
rect 22928 15156 22980 15162
rect 22928 15098 22980 15104
rect 22940 14006 22968 15098
rect 23032 14618 23060 16895
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 23020 13932 23072 13938
rect 23020 13874 23072 13880
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 22940 11778 22968 12242
rect 23032 11898 23060 13874
rect 23124 13462 23152 17020
rect 23216 15094 23244 22766
rect 23480 22568 23532 22574
rect 23478 22536 23480 22545
rect 23532 22536 23534 22545
rect 23478 22471 23534 22480
rect 23572 22500 23624 22506
rect 23572 22442 23624 22448
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 22098 23428 22374
rect 23388 22092 23440 22098
rect 23388 22034 23440 22040
rect 23584 21978 23612 22442
rect 23400 21950 23612 21978
rect 23400 21146 23428 21950
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23492 21418 23520 21830
rect 23676 21554 23704 23054
rect 23846 22672 23902 22681
rect 23846 22607 23902 22616
rect 23756 21888 23808 21894
rect 23756 21830 23808 21836
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23480 21412 23532 21418
rect 23480 21354 23532 21360
rect 23676 21146 23704 21490
rect 23768 21486 23796 21830
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23388 21140 23440 21146
rect 23388 21082 23440 21088
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23768 21078 23796 21286
rect 23756 21072 23808 21078
rect 23756 21014 23808 21020
rect 23480 20800 23532 20806
rect 23480 20742 23532 20748
rect 23386 19952 23442 19961
rect 23386 19887 23442 19896
rect 23296 18624 23348 18630
rect 23400 18601 23428 19887
rect 23492 18737 23520 20742
rect 23768 20602 23796 21014
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23584 18902 23612 20402
rect 23662 20360 23718 20369
rect 23662 20295 23718 20304
rect 23756 20324 23808 20330
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23478 18728 23534 18737
rect 23478 18663 23534 18672
rect 23572 18692 23624 18698
rect 23572 18634 23624 18640
rect 23296 18566 23348 18572
rect 23386 18592 23442 18601
rect 23308 18222 23336 18566
rect 23386 18527 23442 18536
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23308 16794 23336 18158
rect 23296 16788 23348 16794
rect 23296 16730 23348 16736
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23308 15366 23336 16526
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 13530 23244 14282
rect 23308 14278 23336 15302
rect 23400 14929 23428 18362
rect 23584 17882 23612 18634
rect 23572 17876 23624 17882
rect 23572 17818 23624 17824
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 16658 23520 17614
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23478 16008 23534 16017
rect 23478 15943 23534 15952
rect 23492 15910 23520 15943
rect 23480 15904 23532 15910
rect 23480 15846 23532 15852
rect 23386 14920 23442 14929
rect 23386 14855 23442 14864
rect 23400 14600 23428 14855
rect 23400 14572 23520 14600
rect 23492 14414 23520 14572
rect 23572 14476 23624 14482
rect 23572 14418 23624 14424
rect 23480 14408 23532 14414
rect 23584 14385 23612 14418
rect 23480 14350 23532 14356
rect 23570 14376 23626 14385
rect 23570 14311 23626 14320
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23124 12850 23152 13398
rect 23308 13326 23336 14214
rect 23480 13932 23532 13938
rect 23400 13892 23480 13920
rect 23400 13705 23428 13892
rect 23480 13874 23532 13880
rect 23584 13870 23612 14311
rect 23676 14006 23704 20295
rect 23756 20266 23808 20272
rect 23768 19514 23796 20266
rect 23756 19508 23808 19514
rect 23756 19450 23808 19456
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23768 18222 23796 18838
rect 23860 18630 23888 22607
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23756 18216 23808 18222
rect 23756 18158 23808 18164
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23952 18034 23980 23446
rect 24044 19417 24072 24398
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24872 24290 24900 24550
rect 24964 24410 24992 25486
rect 25044 25356 25096 25362
rect 25044 25298 25096 25304
rect 25056 24614 25084 25298
rect 25044 24608 25096 24614
rect 25044 24550 25096 24556
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 24780 24262 24900 24290
rect 24136 24041 24164 24210
rect 24122 24032 24178 24041
rect 24674 24032 24730 24041
rect 24122 23967 24178 23976
rect 24136 23866 24164 23967
rect 24289 23964 24585 23984
rect 24674 23967 24730 23976
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24124 23860 24176 23866
rect 24124 23802 24176 23808
rect 24124 23112 24176 23118
rect 24124 23054 24176 23060
rect 24216 23112 24268 23118
rect 24216 23054 24268 23060
rect 24136 22234 24164 23054
rect 24124 22228 24176 22234
rect 24124 22170 24176 22176
rect 24228 22166 24256 23054
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24216 22160 24268 22166
rect 24216 22102 24268 22108
rect 24596 21978 24624 22170
rect 24688 22137 24716 23967
rect 24780 23089 24808 24262
rect 25148 23866 25176 27095
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24766 23080 24822 23089
rect 24766 23015 24822 23024
rect 24872 22574 24900 23598
rect 24860 22568 24912 22574
rect 24860 22510 24912 22516
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 24766 22264 24822 22273
rect 24766 22199 24822 22208
rect 24674 22128 24730 22137
rect 24674 22063 24730 22072
rect 24596 21950 24716 21978
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24688 21672 24716 21950
rect 24596 21644 24716 21672
rect 24596 20874 24624 21644
rect 24674 21584 24730 21593
rect 24674 21519 24730 21528
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24124 20256 24176 20262
rect 24228 20233 24256 20402
rect 24124 20198 24176 20204
rect 24214 20224 24270 20233
rect 24030 19408 24086 19417
rect 24030 19343 24086 19352
rect 24136 18970 24164 20198
rect 24270 20182 24348 20210
rect 24214 20159 24270 20168
rect 24320 20058 24348 20182
rect 24308 20052 24360 20058
rect 24308 19994 24360 20000
rect 24216 19984 24268 19990
rect 24216 19926 24268 19932
rect 24228 19394 24256 19926
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24228 19378 24348 19394
rect 24228 19372 24360 19378
rect 24228 19366 24308 19372
rect 24308 19314 24360 19320
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24122 18864 24178 18873
rect 24122 18799 24124 18808
rect 24176 18799 24178 18808
rect 24124 18770 24176 18776
rect 24136 18086 24164 18770
rect 24320 18766 24348 19314
rect 24308 18760 24360 18766
rect 24308 18702 24360 18708
rect 24216 18624 24268 18630
rect 24216 18566 24268 18572
rect 24124 18080 24176 18086
rect 23768 17218 23796 18022
rect 23952 18006 24072 18034
rect 24124 18022 24176 18028
rect 23848 17808 23900 17814
rect 23848 17750 23900 17756
rect 23860 17338 23888 17750
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 23768 17190 23888 17218
rect 23756 17060 23808 17066
rect 23756 17002 23808 17008
rect 23768 16250 23796 17002
rect 23756 16244 23808 16250
rect 23756 16186 23808 16192
rect 23754 16144 23810 16153
rect 23754 16079 23810 16088
rect 23768 14521 23796 16079
rect 23860 15473 23888 17190
rect 24044 16810 24072 18006
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 23952 16782 24072 16810
rect 23846 15464 23902 15473
rect 23846 15399 23902 15408
rect 23846 15328 23902 15337
rect 23846 15263 23902 15272
rect 23860 14550 23888 15263
rect 23848 14544 23900 14550
rect 23754 14512 23810 14521
rect 23848 14486 23900 14492
rect 23754 14447 23810 14456
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 23860 13870 23888 14486
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 23848 13864 23900 13870
rect 23848 13806 23900 13812
rect 23480 13728 23532 13734
rect 23386 13696 23442 13705
rect 23480 13670 23532 13676
rect 23386 13631 23442 13640
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23492 13002 23520 13670
rect 23662 13152 23718 13161
rect 23662 13087 23718 13096
rect 23400 12986 23520 13002
rect 23388 12980 23520 12986
rect 23440 12974 23520 12980
rect 23388 12922 23440 12928
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23020 11892 23072 11898
rect 23020 11834 23072 11840
rect 22940 11750 23060 11778
rect 23032 11558 23060 11750
rect 23478 11656 23534 11665
rect 23478 11591 23534 11600
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 10985 23060 11494
rect 23112 11212 23164 11218
rect 23112 11154 23164 11160
rect 23018 10976 23074 10985
rect 23018 10911 23074 10920
rect 23124 10810 23152 11154
rect 23202 11112 23258 11121
rect 23202 11047 23258 11056
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 23216 10010 23244 11047
rect 23492 10130 23520 11591
rect 23584 11354 23612 12582
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23676 10810 23704 13087
rect 23768 12442 23796 13806
rect 23848 13184 23900 13190
rect 23848 13126 23900 13132
rect 23860 12782 23888 13126
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23860 12102 23888 12718
rect 23952 12617 23980 16782
rect 24032 16652 24084 16658
rect 24032 16594 24084 16600
rect 24044 16114 24072 16594
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24032 15632 24084 15638
rect 24032 15574 24084 15580
rect 24044 14414 24072 15574
rect 24136 15162 24164 16934
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 24228 15042 24256 18566
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24320 16794 24348 17138
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24688 16561 24716 21519
rect 24780 19394 24808 22199
rect 25240 22030 25268 22374
rect 25044 22024 25096 22030
rect 25044 21966 25096 21972
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25056 21457 25084 21966
rect 25240 21690 25268 21966
rect 25228 21684 25280 21690
rect 25228 21626 25280 21632
rect 25240 21486 25268 21626
rect 25228 21480 25280 21486
rect 25042 21448 25098 21457
rect 25228 21422 25280 21428
rect 25042 21383 25098 21392
rect 25056 21146 25084 21383
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 19990 24900 20742
rect 25136 20324 25188 20330
rect 25136 20266 25188 20272
rect 24860 19984 24912 19990
rect 24860 19926 24912 19932
rect 25148 19825 25176 20266
rect 25134 19816 25190 19825
rect 25134 19751 25190 19760
rect 25332 19394 25360 27390
rect 25502 24848 25558 24857
rect 25502 24783 25558 24792
rect 24780 19366 24900 19394
rect 24872 18970 24900 19366
rect 25240 19366 25360 19394
rect 25410 19408 25466 19417
rect 25042 19000 25098 19009
rect 24860 18964 24912 18970
rect 25042 18935 25098 18944
rect 24860 18906 24912 18912
rect 25056 18426 25084 18935
rect 25136 18828 25188 18834
rect 25136 18770 25188 18776
rect 25148 18426 25176 18770
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 24768 18216 24820 18222
rect 24768 18158 24820 18164
rect 24780 17898 24808 18158
rect 24780 17882 24900 17898
rect 24780 17876 24912 17882
rect 24780 17870 24860 17876
rect 24860 17818 24912 17824
rect 25240 17218 25268 19366
rect 25410 19343 25466 19352
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25056 17190 25268 17218
rect 24674 16552 24730 16561
rect 24674 16487 24730 16496
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24780 15706 24808 16050
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24674 15464 24730 15473
rect 24674 15399 24730 15408
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24136 15014 24256 15042
rect 24032 14408 24084 14414
rect 24032 14350 24084 14356
rect 23938 12608 23994 12617
rect 23938 12543 23994 12552
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 24032 12096 24084 12102
rect 24032 12038 24084 12044
rect 24044 11830 24072 12038
rect 24032 11824 24084 11830
rect 24032 11766 24084 11772
rect 24032 11620 24084 11626
rect 24032 11562 24084 11568
rect 23940 11552 23992 11558
rect 23940 11494 23992 11500
rect 23952 11014 23980 11494
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23754 10840 23810 10849
rect 23664 10804 23716 10810
rect 23754 10775 23810 10784
rect 23664 10746 23716 10752
rect 23768 10130 23796 10775
rect 23940 10736 23992 10742
rect 23940 10678 23992 10684
rect 23480 10124 23532 10130
rect 23756 10124 23808 10130
rect 23532 10084 23612 10112
rect 23480 10066 23532 10072
rect 23216 9982 23520 10010
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22374 9480 22430 9489
rect 22374 9415 22430 9424
rect 22006 7440 22062 7449
rect 22006 7375 22062 7384
rect 23492 5137 23520 9982
rect 23584 9704 23612 10084
rect 23756 10066 23808 10072
rect 23846 9888 23902 9897
rect 23846 9823 23902 9832
rect 23756 9716 23808 9722
rect 23584 9676 23756 9704
rect 23756 9658 23808 9664
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23478 5128 23534 5137
rect 23478 5063 23534 5072
rect 23478 3496 23534 3505
rect 23478 3431 23534 3440
rect 20442 1456 20498 1465
rect 20442 1391 20498 1400
rect 23492 921 23520 3431
rect 23768 2689 23796 9522
rect 23754 2680 23810 2689
rect 23754 2615 23810 2624
rect 23860 2417 23888 9823
rect 23952 9382 23980 10678
rect 23940 9376 23992 9382
rect 23940 9318 23992 9324
rect 23940 8424 23992 8430
rect 23940 8366 23992 8372
rect 23952 7857 23980 8366
rect 23938 7848 23994 7857
rect 23938 7783 23994 7792
rect 24044 4826 24072 11562
rect 24136 11354 24164 15014
rect 24216 14884 24268 14890
rect 24216 14826 24268 14832
rect 24228 14618 24256 14826
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24584 14000 24636 14006
rect 24584 13942 24636 13948
rect 24596 13682 24624 13942
rect 24688 13802 24716 15399
rect 24780 15162 24808 15642
rect 24858 15192 24914 15201
rect 24768 15156 24820 15162
rect 24858 15127 24914 15136
rect 24768 15098 24820 15104
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24676 13796 24728 13802
rect 24676 13738 24728 13744
rect 24596 13654 24716 13682
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24228 12714 24256 13466
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12708 24268 12714
rect 24216 12650 24268 12656
rect 24228 11880 24256 12650
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24228 11852 24348 11880
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24136 9761 24164 11154
rect 24320 11064 24348 11852
rect 24490 11656 24546 11665
rect 24490 11591 24546 11600
rect 24504 11286 24532 11591
rect 24492 11280 24544 11286
rect 24492 11222 24544 11228
rect 24582 11248 24638 11257
rect 24582 11183 24584 11192
rect 24636 11183 24638 11192
rect 24584 11154 24636 11160
rect 24228 11036 24348 11064
rect 24122 9752 24178 9761
rect 24122 9687 24178 9696
rect 24122 9072 24178 9081
rect 24122 9007 24178 9016
rect 24136 8634 24164 9007
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24122 4720 24178 4729
rect 24122 4655 24178 4664
rect 24136 4282 24164 4655
rect 24228 4622 24256 11036
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24412 10169 24440 10406
rect 24688 10266 24716 13654
rect 24780 13161 24808 14758
rect 24766 13152 24822 13161
rect 24766 13087 24822 13096
rect 24872 13002 24900 15127
rect 25056 14793 25084 17190
rect 25136 17060 25188 17066
rect 25136 17002 25188 17008
rect 25148 16833 25176 17002
rect 25134 16824 25190 16833
rect 25134 16759 25190 16768
rect 25226 16688 25282 16697
rect 25226 16623 25282 16632
rect 25134 16552 25190 16561
rect 25134 16487 25190 16496
rect 25042 14784 25098 14793
rect 25042 14719 25098 14728
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 25056 13938 25084 14418
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 24952 13864 25004 13870
rect 25056 13841 25084 13874
rect 24952 13806 25004 13812
rect 25042 13832 25098 13841
rect 24780 12974 24900 13002
rect 24780 12646 24808 12974
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24860 12640 24912 12646
rect 24860 12582 24912 12588
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24398 10160 24454 10169
rect 24398 10095 24454 10104
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24398 9616 24454 9625
rect 24780 9602 24808 12378
rect 24872 12374 24900 12582
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24872 11762 24900 12310
rect 24964 11898 24992 13806
rect 25042 13767 25098 13776
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 24952 11892 25004 11898
rect 24952 11834 25004 11840
rect 25056 11801 25084 12038
rect 25148 11898 25176 16487
rect 25240 16046 25268 16623
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25240 12209 25268 14350
rect 25332 13394 25360 19246
rect 25424 15162 25452 19343
rect 25516 16250 25544 24783
rect 25594 23352 25650 23361
rect 25700 23322 25728 27639
rect 25962 27520 26018 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 25976 24562 26004 27520
rect 25884 24534 26004 24562
rect 25594 23287 25650 23296
rect 25688 23316 25740 23322
rect 25608 22778 25636 23287
rect 25688 23258 25740 23264
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25596 22568 25648 22574
rect 25596 22510 25648 22516
rect 25608 22030 25636 22510
rect 25792 22438 25820 23122
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25596 22024 25648 22030
rect 25594 21992 25596 22001
rect 25648 21992 25650 22001
rect 25594 21927 25650 21936
rect 25608 21901 25636 21927
rect 25792 19446 25820 22374
rect 25780 19440 25832 19446
rect 25780 19382 25832 19388
rect 25596 19236 25648 19242
rect 25596 19178 25648 19184
rect 25608 18737 25636 19178
rect 25792 19174 25820 19382
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25594 18728 25650 18737
rect 25594 18663 25650 18672
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25504 16244 25556 16250
rect 25504 16186 25556 16192
rect 25504 15904 25556 15910
rect 25504 15846 25556 15852
rect 25412 15156 25464 15162
rect 25412 15098 25464 15104
rect 25412 13932 25464 13938
rect 25412 13874 25464 13880
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25226 12200 25282 12209
rect 25226 12135 25282 12144
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25042 11792 25098 11801
rect 24860 11756 24912 11762
rect 25042 11727 25098 11736
rect 24860 11698 24912 11704
rect 24872 11370 24900 11698
rect 24872 11342 24992 11370
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24872 10810 24900 11154
rect 24964 11150 24992 11342
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 10804 24912 10810
rect 24860 10746 24912 10752
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24964 9722 24992 10066
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 24398 9551 24400 9560
rect 24452 9551 24454 9560
rect 24688 9574 24808 9602
rect 24400 9522 24452 9528
rect 24688 8809 24716 9574
rect 24766 9208 24822 9217
rect 24766 9143 24768 9152
rect 24820 9143 24822 9152
rect 24768 9114 24820 9120
rect 25424 9042 25452 13874
rect 25516 11694 25544 15846
rect 25608 12986 25636 18362
rect 25686 18048 25742 18057
rect 25686 17983 25742 17992
rect 25700 14958 25728 17983
rect 25778 17912 25834 17921
rect 25778 17847 25834 17856
rect 25688 14952 25740 14958
rect 25688 14894 25740 14900
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25504 11688 25556 11694
rect 25504 11630 25556 11636
rect 25792 9994 25820 17847
rect 25780 9988 25832 9994
rect 25780 9930 25832 9936
rect 25884 9081 25912 24534
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 25976 15201 26004 24346
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 26068 21350 26096 22034
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26068 20097 26096 21286
rect 26054 20088 26110 20097
rect 26054 20023 26110 20032
rect 25962 15192 26018 15201
rect 25962 15127 26018 15136
rect 26068 14385 26096 20023
rect 26146 17368 26202 17377
rect 26146 17303 26202 17312
rect 26054 14376 26110 14385
rect 26054 14311 26110 14320
rect 26160 10742 26188 17303
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 26148 10736 26200 10742
rect 26148 10678 26200 10684
rect 26344 9217 26372 14214
rect 26528 9704 26556 27520
rect 27080 14278 27108 27520
rect 27632 25498 27660 27520
rect 27620 25492 27672 25498
rect 27620 25434 27672 25440
rect 27068 14272 27120 14278
rect 27068 14214 27120 14220
rect 26436 9676 26556 9704
rect 26330 9208 26386 9217
rect 26330 9143 26386 9152
rect 25870 9072 25926 9081
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 25412 9036 25464 9042
rect 25870 9007 25926 9016
rect 25412 8978 25464 8984
rect 24766 8936 24822 8945
rect 24766 8871 24822 8880
rect 24674 8800 24730 8809
rect 24289 8732 24585 8752
rect 24674 8735 24730 8744
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24688 6089 24716 8502
rect 24674 6080 24730 6089
rect 24674 6015 24730 6024
rect 24674 5944 24730 5953
rect 24674 5879 24676 5888
rect 24728 5879 24730 5888
rect 24676 5850 24728 5856
rect 24490 5808 24546 5817
rect 24490 5743 24492 5752
rect 24544 5743 24546 5752
rect 24492 5714 24544 5720
rect 24504 5658 24532 5714
rect 24504 5630 24716 5658
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5630
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24676 4752 24728 4758
rect 24490 4720 24546 4729
rect 24676 4694 24728 4700
rect 24490 4655 24492 4664
rect 24544 4655 24546 4664
rect 24492 4626 24544 4632
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 24228 4214 24256 4558
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24216 4208 24268 4214
rect 24688 4162 24716 4694
rect 24780 4593 24808 8871
rect 24964 8634 24992 8978
rect 24952 8628 25004 8634
rect 24952 8570 25004 8576
rect 26436 5953 26464 9676
rect 26422 5944 26478 5953
rect 26422 5879 26478 5888
rect 24766 4584 24822 4593
rect 24766 4519 24822 4528
rect 24216 4150 24268 4156
rect 24596 4134 24716 4162
rect 24596 3942 24624 4134
rect 24584 3936 24636 3942
rect 24582 3904 24584 3913
rect 24636 3904 24638 3913
rect 24582 3839 24638 3848
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 23846 2408 23902 2417
rect 23846 2343 23902 2352
rect 25136 2304 25188 2310
rect 25136 2246 25188 2252
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 23478 912 23534 921
rect 23478 847 23534 856
rect 25148 480 25176 2246
rect 14462 96 14518 105
rect 14462 31 14518 40
rect 19522 0 19578 480
rect 25134 0 25190 480
<< via2 >>
rect 4066 27648 4122 27704
rect 570 23432 626 23488
rect 754 15000 810 15056
rect 570 10668 626 10704
rect 570 10648 572 10668
rect 572 10648 624 10668
rect 624 10648 626 10668
rect 570 7248 626 7304
rect 570 6976 626 7032
rect 1398 22208 1454 22264
rect 1398 22108 1400 22128
rect 1400 22108 1452 22128
rect 1452 22108 1454 22128
rect 1398 22072 1454 22108
rect 1582 23976 1638 24032
rect 1490 21528 1546 21584
rect 1398 21256 1454 21312
rect 1490 21120 1546 21176
rect 1582 19760 1638 19816
rect 1766 22616 1822 22672
rect 1766 21664 1822 21720
rect 1490 16496 1546 16552
rect 1950 25064 2006 25120
rect 3330 27104 3386 27160
rect 25686 27648 25742 27704
rect 3790 26424 3846 26480
rect 3606 25744 3662 25800
rect 2778 25220 2834 25256
rect 2778 25200 2780 25220
rect 2780 25200 2832 25220
rect 2832 25200 2834 25220
rect 2042 24148 2044 24168
rect 2044 24148 2096 24168
rect 2096 24148 2098 24168
rect 2042 24112 2098 24148
rect 2042 22480 2098 22536
rect 2686 24656 2742 24712
rect 2502 24520 2558 24576
rect 2594 23024 2650 23080
rect 2778 22752 2834 22808
rect 2042 20204 2044 20224
rect 2044 20204 2096 20224
rect 2096 20204 2098 20224
rect 2042 20168 2098 20204
rect 2226 20712 2282 20768
rect 1858 18808 1914 18864
rect 1674 17720 1730 17776
rect 2226 17584 2282 17640
rect 2502 20712 2558 20768
rect 2962 22380 2964 22400
rect 2964 22380 3016 22400
rect 3016 22380 3018 22400
rect 2962 22344 3018 22380
rect 3330 22344 3386 22400
rect 2870 20304 2926 20360
rect 2502 18964 2558 19000
rect 2502 18944 2504 18964
rect 2504 18944 2556 18964
rect 2556 18944 2558 18964
rect 2410 18672 2466 18728
rect 1582 15544 1638 15600
rect 1582 14592 1638 14648
rect 2042 14184 2098 14240
rect 2594 14456 2650 14512
rect 2410 14048 2466 14104
rect 2594 13948 2596 13968
rect 2596 13948 2648 13968
rect 2648 13948 2650 13968
rect 2594 13912 2650 13948
rect 2870 19796 2872 19816
rect 2872 19796 2924 19816
rect 2924 19796 2926 19816
rect 2870 19760 2926 19796
rect 3238 17992 3294 18048
rect 3146 16632 3202 16688
rect 2778 14048 2834 14104
rect 3146 14864 3202 14920
rect 2962 13912 3018 13968
rect 3146 13912 3202 13968
rect 3054 12300 3110 12336
rect 3054 12280 3056 12300
rect 3056 12280 3108 12300
rect 3108 12280 3110 12300
rect 2778 3440 2834 3496
rect 1306 2352 1362 2408
rect 4066 25880 4122 25936
rect 4250 26016 4306 26072
rect 4710 25744 4766 25800
rect 3974 23432 4030 23488
rect 3698 23196 3700 23216
rect 3700 23196 3752 23216
rect 3752 23196 3754 23216
rect 3698 23160 3754 23196
rect 4618 21140 4674 21176
rect 4618 21120 4620 21140
rect 4620 21120 4672 21140
rect 4672 21120 4674 21140
rect 3698 20032 3754 20088
rect 3514 17040 3570 17096
rect 3514 15816 3570 15872
rect 3422 11056 3478 11112
rect 2962 3304 3018 3360
rect 2870 1400 2926 1456
rect 3974 19080 4030 19136
rect 3790 17856 3846 17912
rect 3698 15408 3754 15464
rect 3790 14864 3846 14920
rect 4066 16088 4122 16144
rect 3974 15408 4030 15464
rect 4618 20168 4674 20224
rect 4710 19760 4766 19816
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5078 20032 5134 20088
rect 4894 19352 4950 19408
rect 3698 11600 3754 11656
rect 3882 9968 3938 10024
rect 3882 6296 3938 6352
rect 3698 5072 3754 5128
rect 4618 15408 4674 15464
rect 4434 14184 4490 14240
rect 4066 11192 4122 11248
rect 4618 14592 4674 14648
rect 5354 22616 5410 22672
rect 5354 21684 5410 21720
rect 5354 21664 5356 21684
rect 5356 21664 5408 21684
rect 5408 21664 5410 21684
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 6090 21292 6092 21312
rect 6092 21292 6144 21312
rect 6144 21292 6146 21312
rect 6090 21256 6146 21292
rect 5722 20984 5778 21040
rect 6182 20848 6238 20904
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 6366 23860 6422 23896
rect 6366 23840 6368 23860
rect 6368 23840 6420 23860
rect 6420 23840 6422 23860
rect 6734 23044 6790 23080
rect 6734 23024 6736 23044
rect 6736 23024 6788 23044
rect 6788 23024 6790 23044
rect 6918 23160 6974 23216
rect 7654 24656 7710 24712
rect 6734 20712 6790 20768
rect 6642 20168 6698 20224
rect 6366 19896 6422 19952
rect 6366 18944 6422 19000
rect 7102 20460 7158 20496
rect 7102 20440 7104 20460
rect 7104 20440 7156 20460
rect 7156 20440 7158 20460
rect 6918 19488 6974 19544
rect 5446 18536 5502 18592
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5722 18148 5778 18184
rect 5722 18128 5724 18148
rect 5724 18128 5776 18148
rect 5776 18128 5778 18148
rect 6182 17720 6238 17776
rect 6090 17584 6146 17640
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 6274 17584 6330 17640
rect 5538 16904 5594 16960
rect 5354 16768 5410 16824
rect 4986 15852 4988 15872
rect 4988 15852 5040 15872
rect 5040 15852 5042 15872
rect 4986 15816 5042 15852
rect 5262 15408 5318 15464
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5814 14864 5870 14920
rect 4802 13640 4858 13696
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 6274 13504 6330 13560
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 6918 18944 6974 19000
rect 6826 18400 6882 18456
rect 6826 18028 6828 18048
rect 6828 18028 6880 18048
rect 6880 18028 6882 18048
rect 6826 17992 6882 18028
rect 7010 17212 7012 17232
rect 7012 17212 7064 17232
rect 7064 17212 7066 17232
rect 7010 17176 7066 17212
rect 6734 17040 6790 17096
rect 6642 16244 6698 16280
rect 6642 16224 6644 16244
rect 6644 16224 6696 16244
rect 6696 16224 6698 16244
rect 7654 22344 7710 22400
rect 7562 20304 7618 20360
rect 7838 22208 7894 22264
rect 7746 21936 7802 21992
rect 7838 21800 7894 21856
rect 7746 21140 7802 21176
rect 7746 21120 7748 21140
rect 7748 21120 7800 21140
rect 7800 21120 7802 21140
rect 8206 23568 8262 23624
rect 8206 23060 8208 23080
rect 8208 23060 8260 23080
rect 8260 23060 8262 23080
rect 8206 23024 8262 23060
rect 8114 22208 8170 22264
rect 8758 23840 8814 23896
rect 8666 23704 8722 23760
rect 8574 23196 8576 23216
rect 8576 23196 8628 23216
rect 8628 23196 8630 23216
rect 8574 23160 8630 23196
rect 8482 23024 8538 23080
rect 8114 21528 8170 21584
rect 8758 21528 8814 21584
rect 7746 18672 7802 18728
rect 7562 17312 7618 17368
rect 6642 15544 6698 15600
rect 7194 14900 7196 14920
rect 7196 14900 7248 14920
rect 7248 14900 7250 14920
rect 7194 14864 7250 14900
rect 7286 14184 7342 14240
rect 8666 20984 8722 21040
rect 8666 19216 8722 19272
rect 8482 18128 8538 18184
rect 8022 17720 8078 17776
rect 7930 17176 7986 17232
rect 8022 16768 8078 16824
rect 7838 16496 7894 16552
rect 8574 16768 8630 16824
rect 8574 15272 8630 15328
rect 8390 13640 8446 13696
rect 8482 13504 8538 13560
rect 7562 12960 7618 13016
rect 7562 12416 7618 12472
rect 7378 12280 7434 12336
rect 7746 12144 7802 12200
rect 4986 11872 5042 11928
rect 4434 11056 4490 11112
rect 4066 10512 4122 10568
rect 4066 9424 4122 9480
rect 4066 8744 4122 8800
rect 4066 8200 4122 8256
rect 4066 7792 4122 7848
rect 3514 2624 3570 2680
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 8390 12552 8446 12608
rect 8758 17176 8814 17232
rect 8666 12824 8722 12880
rect 9034 24556 9036 24576
rect 9036 24556 9088 24576
rect 9088 24556 9090 24576
rect 9034 24520 9090 24556
rect 9034 24112 9090 24168
rect 9218 20712 9274 20768
rect 8942 16360 8998 16416
rect 8850 12316 8852 12336
rect 8852 12316 8904 12336
rect 8904 12316 8906 12336
rect 8850 12280 8906 12316
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5998 10784 6054 10840
rect 9678 24656 9734 24712
rect 9586 24284 9588 24304
rect 9588 24284 9640 24304
rect 9640 24284 9642 24304
rect 9586 24248 9642 24284
rect 9586 23432 9642 23488
rect 9402 22924 9404 22944
rect 9404 22924 9456 22944
rect 9456 22924 9458 22944
rect 9402 22888 9458 22924
rect 9678 22888 9734 22944
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10874 25472 10930 25528
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9862 23296 9918 23352
rect 9862 22616 9918 22672
rect 9862 21392 9918 21448
rect 9402 20304 9458 20360
rect 9218 16224 9274 16280
rect 9494 20168 9550 20224
rect 9586 19624 9642 19680
rect 9678 17448 9734 17504
rect 9586 16632 9642 16688
rect 9494 15564 9550 15600
rect 9494 15544 9496 15564
rect 9496 15544 9548 15564
rect 9548 15544 9550 15564
rect 8942 10104 8998 10160
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 10138 23840 10194 23896
rect 10690 24112 10746 24168
rect 10230 23568 10286 23624
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10598 22516 10600 22536
rect 10600 22516 10652 22536
rect 10652 22516 10654 22536
rect 10598 22480 10654 22516
rect 10782 22480 10838 22536
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10506 21972 10508 21992
rect 10508 21972 10560 21992
rect 10560 21972 10562 21992
rect 10506 21936 10562 21972
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10138 21120 10194 21176
rect 10782 21120 10838 21176
rect 10046 20848 10102 20904
rect 9954 19488 10010 19544
rect 10782 20596 10838 20632
rect 10782 20576 10784 20596
rect 10784 20576 10836 20596
rect 10836 20576 10838 20596
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10690 19080 10746 19136
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10782 18944 10838 19000
rect 10598 18400 10654 18456
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9862 15952 9918 16008
rect 11702 26016 11758 26072
rect 11150 24556 11152 24576
rect 11152 24556 11204 24576
rect 11204 24556 11206 24576
rect 11150 24520 11206 24556
rect 11426 24556 11428 24576
rect 11428 24556 11480 24576
rect 11480 24556 11482 24576
rect 11426 24520 11482 24556
rect 11334 24112 11390 24168
rect 11242 23840 11298 23896
rect 11058 23604 11060 23624
rect 11060 23604 11112 23624
rect 11112 23604 11114 23624
rect 11058 23568 11114 23604
rect 11242 22752 11298 22808
rect 11334 20304 11390 20360
rect 11058 20168 11114 20224
rect 11334 19624 11390 19680
rect 11426 18128 11482 18184
rect 10138 16940 10140 16960
rect 10140 16940 10192 16960
rect 10192 16940 10194 16960
rect 10138 16904 10194 16940
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10138 16788 10194 16824
rect 10138 16768 10140 16788
rect 10140 16768 10192 16788
rect 10192 16768 10194 16788
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10046 15272 10102 15328
rect 10782 16244 10838 16280
rect 10782 16224 10784 16244
rect 10784 16224 10836 16244
rect 10836 16224 10838 16244
rect 10966 16088 11022 16144
rect 11150 17040 11206 17096
rect 11150 15544 11206 15600
rect 10690 14728 10746 14784
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10138 14492 10140 14512
rect 10140 14492 10192 14512
rect 10192 14492 10194 14512
rect 10138 14456 10194 14492
rect 11242 14184 11298 14240
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 9586 13096 9642 13152
rect 10782 13232 10838 13288
rect 10690 13096 10746 13152
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11150 12824 11206 12880
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 11242 12416 11298 12472
rect 10782 10240 10838 10296
rect 11978 20168 12034 20224
rect 11978 18672 12034 18728
rect 11886 18284 11942 18320
rect 11886 18264 11888 18284
rect 11888 18264 11940 18284
rect 11940 18264 11942 18284
rect 11794 17856 11850 17912
rect 11610 13368 11666 13424
rect 11610 13132 11612 13152
rect 11612 13132 11664 13152
rect 11664 13132 11666 13152
rect 11610 13096 11666 13132
rect 11794 12844 11850 12880
rect 11794 12824 11796 12844
rect 11796 12824 11848 12844
rect 11848 12824 11850 12844
rect 12714 22480 12770 22536
rect 12898 22616 12954 22672
rect 12622 19388 12624 19408
rect 12624 19388 12676 19408
rect 12676 19388 12678 19408
rect 12622 19352 12678 19388
rect 12990 20324 13046 20360
rect 12990 20304 12992 20324
rect 12992 20304 13044 20324
rect 13044 20304 13046 20324
rect 12438 15952 12494 16008
rect 11978 11736 12034 11792
rect 11518 10104 11574 10160
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 9494 3576 9550 3632
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 8298 2896 8354 2952
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 5170 2080 5226 2136
rect 4066 856 4122 912
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12346 10512 12402 10568
rect 12346 9968 12402 10024
rect 12806 16108 12862 16144
rect 12806 16088 12808 16108
rect 12808 16088 12860 16108
rect 12860 16088 12862 16108
rect 13082 19352 13138 19408
rect 13266 23432 13322 23488
rect 13358 22616 13414 22672
rect 13450 22208 13506 22264
rect 12990 15544 13046 15600
rect 12806 14764 12808 14784
rect 12808 14764 12860 14784
rect 12860 14764 12862 14784
rect 12806 14728 12862 14764
rect 13266 16632 13322 16688
rect 13174 15680 13230 15736
rect 13450 14592 13506 14648
rect 13634 24248 13690 24304
rect 14094 24384 14150 24440
rect 14186 23704 14242 23760
rect 14186 22888 14242 22944
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15198 24792 15254 24848
rect 14370 22752 14426 22808
rect 14186 22480 14242 22536
rect 14278 22072 14334 22128
rect 14186 21972 14188 21992
rect 14188 21972 14240 21992
rect 14240 21972 14242 21992
rect 14186 21936 14242 21972
rect 14094 21140 14150 21176
rect 14094 21120 14096 21140
rect 14096 21120 14148 21140
rect 14148 21120 14150 21140
rect 14094 20984 14150 21040
rect 13818 17332 13874 17368
rect 13818 17312 13820 17332
rect 13820 17312 13872 17332
rect 13872 17312 13874 17332
rect 14002 20168 14058 20224
rect 14094 18400 14150 18456
rect 14002 17448 14058 17504
rect 12898 13812 12900 13832
rect 12900 13812 12952 13832
rect 12952 13812 12954 13832
rect 12898 13776 12954 13812
rect 12990 12844 13046 12880
rect 12990 12824 12992 12844
rect 12992 12824 13044 12844
rect 13044 12824 13046 12844
rect 12990 12316 12992 12336
rect 12992 12316 13044 12336
rect 13044 12316 13046 12336
rect 12990 12280 13046 12316
rect 12530 8336 12586 8392
rect 13174 10376 13230 10432
rect 13082 10260 13138 10296
rect 13082 10240 13084 10260
rect 13084 10240 13136 10260
rect 13136 10240 13138 10260
rect 13450 12280 13506 12336
rect 13358 12180 13360 12200
rect 13360 12180 13412 12200
rect 13412 12180 13414 12200
rect 13358 12144 13414 12180
rect 13266 9832 13322 9888
rect 13910 16360 13966 16416
rect 14002 16224 14058 16280
rect 13910 15952 13966 16008
rect 14278 20984 14334 21040
rect 14646 23704 14702 23760
rect 14646 21800 14702 21856
rect 14554 21120 14610 21176
rect 14462 20576 14518 20632
rect 14278 20168 14334 20224
rect 14646 19896 14702 19952
rect 14370 19236 14426 19272
rect 14370 19216 14372 19236
rect 14372 19216 14424 19236
rect 14424 19216 14426 19236
rect 14462 17720 14518 17776
rect 15198 24384 15254 24440
rect 15290 24268 15346 24304
rect 15290 24248 15292 24268
rect 15292 24248 15344 24268
rect 15344 24248 15346 24268
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15290 23296 15346 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15934 25472 15990 25528
rect 17498 25880 17554 25936
rect 15474 24148 15476 24168
rect 15476 24148 15528 24168
rect 15528 24148 15530 24168
rect 15474 24112 15530 24148
rect 15474 23568 15530 23624
rect 15382 22616 15438 22672
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14646 17856 14702 17912
rect 13726 15000 13782 15056
rect 14094 14492 14096 14512
rect 14096 14492 14148 14512
rect 14148 14492 14150 14512
rect 14094 14456 14150 14492
rect 13726 11620 13782 11656
rect 13726 11600 13728 11620
rect 13728 11600 13780 11620
rect 13780 11600 13782 11620
rect 14094 13640 14150 13696
rect 14094 12960 14150 13016
rect 13910 11192 13966 11248
rect 13542 9560 13598 9616
rect 13450 9424 13506 9480
rect 13910 3576 13966 3632
rect 12162 3440 12218 3496
rect 12898 3440 12954 3496
rect 12438 2896 12494 2952
rect 14462 16496 14518 16552
rect 14462 15852 14464 15872
rect 14464 15852 14516 15872
rect 14516 15852 14518 15872
rect 14462 15816 14518 15852
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15382 20848 15438 20904
rect 15290 20168 15346 20224
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 15014 18964 15070 19000
rect 15014 18944 15016 18964
rect 15016 18944 15068 18964
rect 15068 18944 15070 18964
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14646 15156 14702 15192
rect 14646 15136 14648 15156
rect 14648 15136 14700 15156
rect 14700 15136 14702 15156
rect 14462 13776 14518 13832
rect 3422 312 3478 368
rect 14554 11756 14610 11792
rect 14554 11736 14556 11756
rect 14556 11736 14608 11756
rect 14608 11736 14610 11756
rect 14922 17604 14978 17640
rect 14922 17584 14924 17604
rect 14924 17584 14976 17604
rect 14976 17584 14978 17604
rect 15106 17584 15162 17640
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14922 17176 14978 17232
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15474 19080 15530 19136
rect 15474 16668 15476 16688
rect 15476 16668 15528 16688
rect 15528 16668 15530 16688
rect 15474 16632 15530 16668
rect 15382 16496 15438 16552
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14830 13368 14886 13424
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15658 23840 15714 23896
rect 15750 22072 15806 22128
rect 15750 20576 15806 20632
rect 15658 19352 15714 19408
rect 16302 23432 16358 23488
rect 16118 22888 16174 22944
rect 16302 22616 16358 22672
rect 16026 22480 16082 22536
rect 15934 21412 15990 21448
rect 15934 21392 15936 21412
rect 15936 21392 15988 21412
rect 15988 21392 15990 21412
rect 16118 21548 16174 21584
rect 16118 21528 16120 21548
rect 16120 21528 16172 21548
rect 16172 21528 16174 21548
rect 15566 12008 15622 12064
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 16762 24384 16818 24440
rect 16486 20032 16542 20088
rect 16486 18808 16542 18864
rect 16486 16496 16542 16552
rect 16670 16360 16726 16416
rect 16670 15952 16726 16008
rect 16578 15408 16634 15464
rect 17590 24792 17646 24848
rect 17498 23976 17554 24032
rect 17038 20984 17094 21040
rect 16854 19896 16910 19952
rect 17406 21256 17462 21312
rect 17498 21120 17554 21176
rect 17774 22344 17830 22400
rect 18142 23060 18144 23080
rect 18144 23060 18196 23080
rect 18196 23060 18198 23080
rect 18142 23024 18198 23060
rect 17130 17992 17186 18048
rect 17314 17992 17370 18048
rect 17038 17740 17094 17776
rect 17038 17720 17040 17740
rect 17040 17720 17092 17740
rect 17092 17720 17094 17740
rect 16854 15972 16910 16008
rect 16854 15952 16856 15972
rect 16856 15952 16908 15972
rect 16908 15952 16910 15972
rect 16854 15816 16910 15872
rect 16486 11600 16542 11656
rect 16394 10784 16450 10840
rect 15750 8880 15806 8936
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 16394 7928 16450 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 16854 7384 16910 7440
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 17314 14864 17370 14920
rect 17314 12416 17370 12472
rect 17314 11192 17370 11248
rect 17774 18944 17830 19000
rect 18510 24656 18566 24712
rect 18326 23976 18382 24032
rect 18418 21392 18474 21448
rect 18418 21120 18474 21176
rect 19154 24676 19210 24712
rect 19154 24656 19156 24676
rect 19156 24656 19208 24676
rect 19208 24656 19210 24676
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19338 24792 19394 24848
rect 19246 24520 19302 24576
rect 18970 24148 18972 24168
rect 18972 24148 19024 24168
rect 19024 24148 19026 24168
rect 18970 24112 19026 24148
rect 18786 23024 18842 23080
rect 18510 20168 18566 20224
rect 18234 19352 18290 19408
rect 18510 19236 18566 19272
rect 18510 19216 18512 19236
rect 18512 19216 18564 19236
rect 18564 19216 18566 19236
rect 18418 18672 18474 18728
rect 17774 17604 17830 17640
rect 17774 17584 17776 17604
rect 17776 17584 17828 17604
rect 17828 17584 17830 17604
rect 18786 18400 18842 18456
rect 18510 16496 18566 16552
rect 17774 15408 17830 15464
rect 17866 15156 17922 15192
rect 17866 15136 17868 15156
rect 17868 15136 17920 15156
rect 17920 15136 17922 15156
rect 18694 15136 18750 15192
rect 17682 13640 17738 13696
rect 18786 11872 18842 11928
rect 17130 9560 17186 9616
rect 17038 3984 17094 4040
rect 17590 11056 17646 11112
rect 19246 23568 19302 23624
rect 19154 22072 19210 22128
rect 19522 24792 19578 24848
rect 19430 24384 19486 24440
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19522 24248 19578 24304
rect 19522 23976 19578 24032
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19430 22616 19486 22672
rect 19706 22616 19762 22672
rect 19430 21836 19432 21856
rect 19432 21836 19484 21856
rect 19484 21836 19486 21856
rect 19430 21800 19486 21836
rect 19154 19760 19210 19816
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19522 20576 19578 20632
rect 19338 20304 19394 20360
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19706 19352 19762 19408
rect 19430 18264 19486 18320
rect 19338 17992 19394 18048
rect 19246 17720 19302 17776
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 20534 25744 20590 25800
rect 20166 24248 20222 24304
rect 20074 23432 20130 23488
rect 20350 22072 20406 22128
rect 20718 23740 20720 23760
rect 20720 23740 20772 23760
rect 20772 23740 20774 23760
rect 20718 23704 20774 23740
rect 20718 22888 20774 22944
rect 19154 12688 19210 12744
rect 19430 12588 19432 12608
rect 19432 12588 19484 12608
rect 19484 12588 19486 12608
rect 19430 12552 19486 12588
rect 19982 15952 20038 16008
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 20350 19624 20406 19680
rect 20534 21392 20590 21448
rect 21362 24248 21418 24304
rect 21454 23840 21510 23896
rect 21362 23588 21418 23624
rect 21362 23568 21364 23588
rect 21364 23568 21416 23588
rect 21416 23568 21418 23588
rect 21822 23976 21878 24032
rect 22282 24792 22338 24848
rect 22650 24792 22706 24848
rect 21270 22072 21326 22128
rect 21914 21800 21970 21856
rect 20718 20440 20774 20496
rect 20902 19896 20958 19952
rect 20994 18672 21050 18728
rect 20258 15952 20314 16008
rect 20258 15544 20314 15600
rect 20810 16632 20866 16688
rect 20902 16088 20958 16144
rect 20626 15272 20682 15328
rect 20074 8200 20130 8256
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 20994 10784 21050 10840
rect 21638 20576 21694 20632
rect 21546 18944 21602 19000
rect 21730 19080 21786 19136
rect 21638 17584 21694 17640
rect 21454 15136 21510 15192
rect 21270 12144 21326 12200
rect 21546 14456 21602 14512
rect 21914 18944 21970 19000
rect 22098 18536 22154 18592
rect 22006 15272 22062 15328
rect 22006 13640 22062 13696
rect 21914 13368 21970 13424
rect 21638 10648 21694 10704
rect 21178 10512 21234 10568
rect 20442 8336 20498 8392
rect 20166 6976 20222 7032
rect 17498 6296 17554 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 17314 3576 17370 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 18510 2372 18566 2408
rect 18510 2352 18512 2372
rect 18512 2352 18564 2372
rect 18564 2352 18566 2372
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 22466 24656 22522 24712
rect 22650 24132 22706 24168
rect 22650 24112 22652 24132
rect 22652 24112 22704 24132
rect 22704 24112 22706 24132
rect 22282 19216 22338 19272
rect 22282 18028 22284 18048
rect 22284 18028 22336 18048
rect 22336 18028 22338 18048
rect 22282 17992 22338 18028
rect 22282 17720 22338 17776
rect 22282 11892 22338 11928
rect 22282 11872 22284 11892
rect 22284 11872 22336 11892
rect 22336 11872 22338 11892
rect 22466 19760 22522 19816
rect 22466 16632 22522 16688
rect 22650 18400 22706 18456
rect 22650 15408 22706 15464
rect 22558 15000 22614 15056
rect 22834 24656 22890 24712
rect 24766 26424 24822 26480
rect 24674 25880 24730 25936
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 25134 27104 25190 27160
rect 24766 25220 24822 25256
rect 24766 25200 24768 25220
rect 24768 25200 24820 25220
rect 24820 25200 24822 25220
rect 23386 23160 23442 23216
rect 23662 23432 23718 23488
rect 23018 20204 23020 20224
rect 23020 20204 23072 20224
rect 23072 20204 23074 20224
rect 23018 20168 23074 20204
rect 22834 19760 22890 19816
rect 23018 16904 23074 16960
rect 22926 16788 22982 16824
rect 22926 16768 22928 16788
rect 22928 16768 22980 16788
rect 22980 16768 22982 16788
rect 22558 12280 22614 12336
rect 22742 12280 22798 12336
rect 22742 12008 22798 12064
rect 22650 11328 22706 11384
rect 23478 22516 23480 22536
rect 23480 22516 23532 22536
rect 23532 22516 23534 22536
rect 23478 22480 23534 22516
rect 23846 22616 23902 22672
rect 23386 19896 23442 19952
rect 23662 20304 23718 20360
rect 23478 18672 23534 18728
rect 23386 18536 23442 18592
rect 23478 15952 23534 16008
rect 23386 14864 23442 14920
rect 23570 14320 23626 14376
rect 24122 23976 24178 24032
rect 24674 23976 24730 24032
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 24766 23024 24822 23080
rect 24766 22208 24822 22264
rect 24674 22072 24730 22128
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21528 24730 21584
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24030 19352 24086 19408
rect 24214 20168 24270 20224
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24122 18828 24178 18864
rect 24122 18808 24124 18828
rect 24124 18808 24176 18828
rect 24176 18808 24178 18828
rect 23754 16088 23810 16144
rect 23846 15408 23902 15464
rect 23846 15272 23902 15328
rect 23754 14456 23810 14512
rect 23386 13640 23442 13696
rect 23662 13096 23718 13152
rect 23478 11600 23534 11656
rect 23018 10920 23074 10976
rect 23202 11056 23258 11112
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 25042 21392 25098 21448
rect 25134 19760 25190 19816
rect 25502 24792 25558 24848
rect 25042 18944 25098 19000
rect 25410 19352 25466 19408
rect 24674 16496 24730 16552
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24674 15408 24730 15464
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 23938 12552 23994 12608
rect 23754 10784 23810 10840
rect 22374 9424 22430 9480
rect 22006 7384 22062 7440
rect 23846 9832 23902 9888
rect 23478 5072 23534 5128
rect 23478 3440 23534 3496
rect 20442 1400 20498 1456
rect 23754 2624 23810 2680
rect 23938 7792 23994 7848
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24858 15136 24914 15192
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24490 11600 24546 11656
rect 24582 11212 24638 11248
rect 24582 11192 24584 11212
rect 24584 11192 24636 11212
rect 24636 11192 24638 11212
rect 24122 9696 24178 9752
rect 24122 9016 24178 9072
rect 24122 4664 24178 4720
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24766 13096 24822 13152
rect 25134 16768 25190 16824
rect 25226 16632 25282 16688
rect 25134 16496 25190 16552
rect 25042 14728 25098 14784
rect 24398 10104 24454 10160
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24398 9580 24454 9616
rect 25042 13776 25098 13832
rect 25594 23296 25650 23352
rect 25594 21972 25596 21992
rect 25596 21972 25648 21992
rect 25648 21972 25650 21992
rect 25594 21936 25650 21972
rect 25594 18672 25650 18728
rect 25226 12144 25282 12200
rect 25042 11736 25098 11792
rect 24398 9560 24400 9580
rect 24400 9560 24452 9580
rect 24452 9560 24454 9580
rect 24766 9172 24822 9208
rect 24766 9152 24768 9172
rect 24768 9152 24820 9172
rect 24820 9152 24822 9172
rect 25686 17992 25742 18048
rect 25778 17856 25834 17912
rect 26054 20032 26110 20088
rect 25962 15136 26018 15192
rect 26146 17312 26202 17368
rect 26054 14320 26110 14376
rect 26330 9152 26386 9208
rect 25870 9016 25926 9072
rect 24766 8880 24822 8936
rect 24674 8744 24730 8800
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24674 6024 24730 6080
rect 24674 5908 24730 5944
rect 24674 5888 24676 5908
rect 24676 5888 24728 5908
rect 24728 5888 24730 5908
rect 24490 5772 24546 5808
rect 24490 5752 24492 5772
rect 24492 5752 24544 5772
rect 24544 5752 24546 5772
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24490 4684 24546 4720
rect 24490 4664 24492 4684
rect 24492 4664 24544 4684
rect 24544 4664 24546 4684
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 26422 5888 26478 5944
rect 24766 4528 24822 4584
rect 24582 3884 24584 3904
rect 24584 3884 24636 3904
rect 24636 3884 24638 3904
rect 24582 3848 24638 3884
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 23846 2352 23902 2408
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 23478 856 23534 912
rect 14462 40 14518 96
<< metal3 >>
rect 0 27706 480 27736
rect 4061 27706 4127 27709
rect 0 27704 4127 27706
rect 0 27648 4066 27704
rect 4122 27648 4127 27704
rect 0 27646 4127 27648
rect 0 27616 480 27646
rect 4061 27643 4127 27646
rect 25681 27706 25747 27709
rect 27520 27706 28000 27736
rect 25681 27704 28000 27706
rect 25681 27648 25686 27704
rect 25742 27648 28000 27704
rect 25681 27646 28000 27648
rect 25681 27643 25747 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 3325 27162 3391 27165
rect 0 27160 3391 27162
rect 0 27104 3330 27160
rect 3386 27104 3391 27160
rect 0 27102 3391 27104
rect 0 27072 480 27102
rect 3325 27099 3391 27102
rect 25129 27162 25195 27165
rect 27520 27162 28000 27192
rect 25129 27160 28000 27162
rect 25129 27104 25134 27160
rect 25190 27104 28000 27160
rect 25129 27102 28000 27104
rect 25129 27099 25195 27102
rect 27520 27072 28000 27102
rect 0 26482 480 26512
rect 3785 26482 3851 26485
rect 0 26480 3851 26482
rect 0 26424 3790 26480
rect 3846 26424 3851 26480
rect 0 26422 3851 26424
rect 0 26392 480 26422
rect 3785 26419 3851 26422
rect 24761 26482 24827 26485
rect 27520 26482 28000 26512
rect 24761 26480 28000 26482
rect 24761 26424 24766 26480
rect 24822 26424 28000 26480
rect 24761 26422 28000 26424
rect 24761 26419 24827 26422
rect 27520 26392 28000 26422
rect 4245 26074 4311 26077
rect 11697 26074 11763 26077
rect 4245 26072 11763 26074
rect 4245 26016 4250 26072
rect 4306 26016 11702 26072
rect 11758 26016 11763 26072
rect 4245 26014 11763 26016
rect 4245 26011 4311 26014
rect 11697 26011 11763 26014
rect 0 25938 480 25968
rect 4061 25938 4127 25941
rect 17493 25938 17559 25941
rect 0 25936 4127 25938
rect 0 25880 4066 25936
rect 4122 25880 4127 25936
rect 0 25878 4127 25880
rect 0 25848 480 25878
rect 4061 25875 4127 25878
rect 4478 25936 17559 25938
rect 4478 25880 17498 25936
rect 17554 25880 17559 25936
rect 4478 25878 17559 25880
rect 3601 25802 3667 25805
rect 4478 25802 4538 25878
rect 17493 25875 17559 25878
rect 24669 25938 24735 25941
rect 27520 25938 28000 25968
rect 24669 25936 28000 25938
rect 24669 25880 24674 25936
rect 24730 25880 28000 25936
rect 24669 25878 28000 25880
rect 24669 25875 24735 25878
rect 27520 25848 28000 25878
rect 3601 25800 4538 25802
rect 3601 25744 3606 25800
rect 3662 25744 4538 25800
rect 3601 25742 4538 25744
rect 4705 25802 4771 25805
rect 20529 25802 20595 25805
rect 4705 25800 20595 25802
rect 4705 25744 4710 25800
rect 4766 25744 20534 25800
rect 20590 25744 20595 25800
rect 4705 25742 20595 25744
rect 3601 25739 3667 25742
rect 4705 25739 4771 25742
rect 20529 25739 20595 25742
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 10869 25530 10935 25533
rect 15929 25530 15995 25533
rect 10869 25528 15995 25530
rect 10869 25472 10874 25528
rect 10930 25472 15934 25528
rect 15990 25472 15995 25528
rect 10869 25470 15995 25472
rect 10869 25467 10935 25470
rect 15929 25467 15995 25470
rect 0 25258 480 25288
rect 2773 25258 2839 25261
rect 0 25256 2839 25258
rect 0 25200 2778 25256
rect 2834 25200 2839 25256
rect 0 25198 2839 25200
rect 0 25168 480 25198
rect 2773 25195 2839 25198
rect 24761 25258 24827 25261
rect 27520 25258 28000 25288
rect 24761 25256 28000 25258
rect 24761 25200 24766 25256
rect 24822 25200 28000 25256
rect 24761 25198 28000 25200
rect 24761 25195 24827 25198
rect 27520 25168 28000 25198
rect 1945 25122 2011 25125
rect 1945 25120 5136 25122
rect 1945 25064 1950 25120
rect 2006 25064 5136 25120
rect 1945 25062 5136 25064
rect 1945 25059 2011 25062
rect 5076 24850 5136 25062
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 15193 24850 15259 24853
rect 5076 24848 15259 24850
rect 5076 24792 15198 24848
rect 15254 24792 15259 24848
rect 5076 24790 15259 24792
rect 15193 24787 15259 24790
rect 17585 24850 17651 24853
rect 19333 24850 19399 24853
rect 17585 24848 19399 24850
rect 17585 24792 17590 24848
rect 17646 24792 19338 24848
rect 19394 24792 19399 24848
rect 17585 24790 19399 24792
rect 17585 24787 17651 24790
rect 19333 24787 19399 24790
rect 19517 24850 19583 24853
rect 22277 24850 22343 24853
rect 19517 24848 22343 24850
rect 19517 24792 19522 24848
rect 19578 24792 22282 24848
rect 22338 24792 22343 24848
rect 19517 24790 22343 24792
rect 19517 24787 19583 24790
rect 22277 24787 22343 24790
rect 22645 24850 22711 24853
rect 25497 24850 25563 24853
rect 22645 24848 25563 24850
rect 22645 24792 22650 24848
rect 22706 24792 25502 24848
rect 25558 24792 25563 24848
rect 22645 24790 25563 24792
rect 22645 24787 22711 24790
rect 25497 24787 25563 24790
rect 0 24714 480 24744
rect 2681 24714 2747 24717
rect 0 24712 2747 24714
rect 0 24656 2686 24712
rect 2742 24656 2747 24712
rect 0 24654 2747 24656
rect 0 24624 480 24654
rect 2681 24651 2747 24654
rect 7649 24714 7715 24717
rect 9673 24714 9739 24717
rect 7649 24712 9739 24714
rect 7649 24656 7654 24712
rect 7710 24656 9678 24712
rect 9734 24656 9739 24712
rect 7649 24654 9739 24656
rect 7649 24651 7715 24654
rect 9673 24651 9739 24654
rect 18505 24714 18571 24717
rect 19149 24714 19215 24717
rect 22461 24714 22527 24717
rect 18505 24712 22527 24714
rect 18505 24656 18510 24712
rect 18566 24656 19154 24712
rect 19210 24656 22466 24712
rect 22522 24656 22527 24712
rect 18505 24654 22527 24656
rect 18505 24651 18571 24654
rect 19149 24651 19215 24654
rect 22461 24651 22527 24654
rect 22829 24714 22895 24717
rect 27520 24714 28000 24744
rect 22829 24712 28000 24714
rect 22829 24656 22834 24712
rect 22890 24656 28000 24712
rect 22829 24654 28000 24656
rect 22829 24651 22895 24654
rect 27520 24624 28000 24654
rect 2497 24578 2563 24581
rect 9029 24578 9095 24581
rect 2497 24576 9095 24578
rect 2497 24520 2502 24576
rect 2558 24520 9034 24576
rect 9090 24520 9095 24576
rect 2497 24518 9095 24520
rect 2497 24515 2563 24518
rect 9029 24515 9095 24518
rect 11145 24578 11211 24581
rect 11278 24578 11284 24580
rect 11145 24576 11284 24578
rect 11145 24520 11150 24576
rect 11206 24520 11284 24576
rect 11145 24518 11284 24520
rect 11145 24515 11211 24518
rect 11278 24516 11284 24518
rect 11348 24516 11354 24580
rect 11421 24578 11487 24581
rect 19241 24578 19307 24581
rect 11421 24576 19307 24578
rect 11421 24520 11426 24576
rect 11482 24520 19246 24576
rect 19302 24520 19307 24576
rect 11421 24518 19307 24520
rect 11421 24515 11487 24518
rect 19241 24515 19307 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 13854 24380 13860 24444
rect 13924 24442 13930 24444
rect 14089 24442 14155 24445
rect 13924 24440 14155 24442
rect 13924 24384 14094 24440
rect 14150 24384 14155 24440
rect 13924 24382 14155 24384
rect 13924 24380 13930 24382
rect 14089 24379 14155 24382
rect 15193 24442 15259 24445
rect 16757 24442 16823 24445
rect 19425 24442 19491 24445
rect 15193 24440 19491 24442
rect 15193 24384 15198 24440
rect 15254 24384 16762 24440
rect 16818 24384 19430 24440
rect 19486 24384 19491 24440
rect 15193 24382 19491 24384
rect 15193 24379 15259 24382
rect 16757 24379 16823 24382
rect 19425 24379 19491 24382
rect 9581 24306 9647 24309
rect 13629 24306 13695 24309
rect 9581 24304 13695 24306
rect 9581 24248 9586 24304
rect 9642 24248 13634 24304
rect 13690 24248 13695 24304
rect 9581 24246 13695 24248
rect 9581 24243 9647 24246
rect 13629 24243 13695 24246
rect 15285 24306 15351 24309
rect 19517 24306 19583 24309
rect 15285 24304 19583 24306
rect 15285 24248 15290 24304
rect 15346 24248 19522 24304
rect 19578 24248 19583 24304
rect 15285 24246 19583 24248
rect 15285 24243 15351 24246
rect 19517 24243 19583 24246
rect 20161 24306 20227 24309
rect 21357 24306 21423 24309
rect 20161 24304 21423 24306
rect 20161 24248 20166 24304
rect 20222 24248 21362 24304
rect 21418 24248 21423 24304
rect 20161 24246 21423 24248
rect 20161 24243 20227 24246
rect 21357 24243 21423 24246
rect 2037 24170 2103 24173
rect 9029 24170 9095 24173
rect 2037 24168 9095 24170
rect 2037 24112 2042 24168
rect 2098 24112 9034 24168
rect 9090 24112 9095 24168
rect 2037 24110 9095 24112
rect 2037 24107 2103 24110
rect 9029 24107 9095 24110
rect 10685 24170 10751 24173
rect 11329 24170 11395 24173
rect 15469 24170 15535 24173
rect 10685 24168 15535 24170
rect 10685 24112 10690 24168
rect 10746 24112 11334 24168
rect 11390 24112 15474 24168
rect 15530 24112 15535 24168
rect 10685 24110 15535 24112
rect 10685 24107 10751 24110
rect 11329 24107 11395 24110
rect 15469 24107 15535 24110
rect 18965 24170 19031 24173
rect 22645 24170 22711 24173
rect 18965 24168 22711 24170
rect 18965 24112 18970 24168
rect 19026 24112 22650 24168
rect 22706 24112 22711 24168
rect 18965 24110 22711 24112
rect 18965 24107 19031 24110
rect 22645 24107 22711 24110
rect 0 24034 480 24064
rect 1577 24034 1643 24037
rect 0 24032 1643 24034
rect 0 23976 1582 24032
rect 1638 23976 1643 24032
rect 0 23974 1643 23976
rect 0 23944 480 23974
rect 1577 23971 1643 23974
rect 17493 24034 17559 24037
rect 18321 24034 18387 24037
rect 19517 24034 19583 24037
rect 17493 24032 19583 24034
rect 17493 23976 17498 24032
rect 17554 23976 18326 24032
rect 18382 23976 19522 24032
rect 19578 23976 19583 24032
rect 17493 23974 19583 23976
rect 17493 23971 17559 23974
rect 18321 23971 18387 23974
rect 19517 23971 19583 23974
rect 21817 24034 21883 24037
rect 24117 24034 24183 24037
rect 21817 24032 24183 24034
rect 21817 23976 21822 24032
rect 21878 23976 24122 24032
rect 24178 23976 24183 24032
rect 21817 23974 24183 23976
rect 21817 23971 21883 23974
rect 24117 23971 24183 23974
rect 24669 24034 24735 24037
rect 27520 24034 28000 24064
rect 24669 24032 28000 24034
rect 24669 23976 24674 24032
rect 24730 23976 28000 24032
rect 24669 23974 28000 23976
rect 24669 23971 24735 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 27520 23944 28000 23974
rect 24277 23903 24597 23904
rect 6361 23898 6427 23901
rect 8753 23898 8819 23901
rect 6361 23896 8819 23898
rect 6361 23840 6366 23896
rect 6422 23840 8758 23896
rect 8814 23840 8819 23896
rect 6361 23838 8819 23840
rect 6361 23835 6427 23838
rect 8753 23835 8819 23838
rect 10133 23898 10199 23901
rect 11237 23898 11303 23901
rect 10133 23896 11303 23898
rect 10133 23840 10138 23896
rect 10194 23840 11242 23896
rect 11298 23840 11303 23896
rect 10133 23838 11303 23840
rect 10133 23835 10199 23838
rect 11237 23835 11303 23838
rect 15653 23898 15719 23901
rect 21449 23898 21515 23901
rect 15653 23896 21515 23898
rect 15653 23840 15658 23896
rect 15714 23840 21454 23896
rect 21510 23840 21515 23896
rect 15653 23838 21515 23840
rect 15653 23835 15719 23838
rect 21449 23835 21515 23838
rect 8661 23762 8727 23765
rect 14181 23762 14247 23765
rect 8661 23760 14247 23762
rect 8661 23704 8666 23760
rect 8722 23704 14186 23760
rect 14242 23704 14247 23760
rect 8661 23702 14247 23704
rect 8661 23699 8727 23702
rect 14181 23699 14247 23702
rect 14641 23762 14707 23765
rect 20713 23762 20779 23765
rect 14641 23760 20779 23762
rect 14641 23704 14646 23760
rect 14702 23704 20718 23760
rect 20774 23704 20779 23760
rect 14641 23702 20779 23704
rect 14641 23699 14707 23702
rect 20713 23699 20779 23702
rect 8201 23626 8267 23629
rect 10225 23626 10291 23629
rect 11053 23626 11119 23629
rect 15469 23626 15535 23629
rect 8201 23624 10794 23626
rect 8201 23568 8206 23624
rect 8262 23568 10230 23624
rect 10286 23568 10794 23624
rect 8201 23566 10794 23568
rect 8201 23563 8267 23566
rect 10225 23563 10291 23566
rect 0 23490 480 23520
rect 565 23490 631 23493
rect 0 23488 631 23490
rect 0 23432 570 23488
rect 626 23432 631 23488
rect 0 23430 631 23432
rect 0 23400 480 23430
rect 565 23427 631 23430
rect 3969 23490 4035 23493
rect 9581 23490 9647 23493
rect 3969 23488 9647 23490
rect 3969 23432 3974 23488
rect 4030 23432 9586 23488
rect 9642 23432 9647 23488
rect 3969 23430 9647 23432
rect 3969 23427 4035 23430
rect 9581 23427 9647 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 9857 23354 9923 23357
rect 7054 23352 9923 23354
rect 7054 23296 9862 23352
rect 9918 23296 9923 23352
rect 7054 23294 9923 23296
rect 10734 23354 10794 23566
rect 11053 23624 15535 23626
rect 11053 23568 11058 23624
rect 11114 23568 15474 23624
rect 15530 23568 15535 23624
rect 11053 23566 15535 23568
rect 11053 23563 11119 23566
rect 15469 23563 15535 23566
rect 19241 23626 19307 23629
rect 21357 23626 21423 23629
rect 19241 23624 21423 23626
rect 19241 23568 19246 23624
rect 19302 23568 21362 23624
rect 21418 23568 21423 23624
rect 19241 23566 21423 23568
rect 19241 23563 19307 23566
rect 21357 23563 21423 23566
rect 13261 23490 13327 23493
rect 16297 23490 16363 23493
rect 13261 23488 16363 23490
rect 13261 23432 13266 23488
rect 13322 23432 16302 23488
rect 16358 23432 16363 23488
rect 13261 23430 16363 23432
rect 13261 23427 13327 23430
rect 16297 23427 16363 23430
rect 20069 23490 20135 23493
rect 23657 23490 23723 23493
rect 27520 23490 28000 23520
rect 20069 23488 23723 23490
rect 20069 23432 20074 23488
rect 20130 23432 23662 23488
rect 23718 23432 23723 23488
rect 20069 23430 23723 23432
rect 20069 23427 20135 23430
rect 23657 23427 23723 23430
rect 25592 23430 28000 23490
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 25592 23357 25652 23430
rect 27520 23400 28000 23430
rect 15285 23354 15351 23357
rect 10734 23352 15351 23354
rect 10734 23296 15290 23352
rect 15346 23296 15351 23352
rect 10734 23294 15351 23296
rect 3693 23218 3759 23221
rect 6913 23218 6979 23221
rect 7054 23218 7114 23294
rect 9857 23291 9923 23294
rect 15285 23291 15351 23294
rect 25589 23352 25655 23357
rect 25589 23296 25594 23352
rect 25650 23296 25655 23352
rect 25589 23291 25655 23296
rect 3693 23216 7114 23218
rect 3693 23160 3698 23216
rect 3754 23160 6918 23216
rect 6974 23160 7114 23216
rect 3693 23158 7114 23160
rect 8569 23218 8635 23221
rect 23381 23218 23447 23221
rect 8569 23216 23447 23218
rect 8569 23160 8574 23216
rect 8630 23160 23386 23216
rect 23442 23160 23447 23216
rect 8569 23158 23447 23160
rect 3693 23155 3759 23158
rect 6913 23155 6979 23158
rect 8569 23155 8635 23158
rect 23381 23155 23447 23158
rect 2589 23082 2655 23085
rect 6729 23082 6795 23085
rect 2589 23080 6795 23082
rect 2589 23024 2594 23080
rect 2650 23024 6734 23080
rect 6790 23024 6795 23080
rect 2589 23022 6795 23024
rect 2589 23019 2655 23022
rect 6729 23019 6795 23022
rect 8201 23082 8267 23085
rect 8477 23082 8543 23085
rect 18137 23082 18203 23085
rect 8201 23080 18203 23082
rect 8201 23024 8206 23080
rect 8262 23024 8482 23080
rect 8538 23024 18142 23080
rect 18198 23024 18203 23080
rect 8201 23022 18203 23024
rect 8201 23019 8267 23022
rect 8477 23019 8543 23022
rect 18137 23019 18203 23022
rect 18781 23082 18847 23085
rect 24761 23082 24827 23085
rect 18781 23080 24827 23082
rect 18781 23024 18786 23080
rect 18842 23024 24766 23080
rect 24822 23024 24827 23080
rect 18781 23022 24827 23024
rect 18781 23019 18847 23022
rect 24761 23019 24827 23022
rect 9397 22946 9463 22949
rect 9673 22946 9739 22949
rect 14181 22946 14247 22949
rect 9397 22944 14247 22946
rect 9397 22888 9402 22944
rect 9458 22888 9678 22944
rect 9734 22888 14186 22944
rect 14242 22888 14247 22944
rect 9397 22886 14247 22888
rect 9397 22883 9463 22886
rect 9673 22883 9739 22886
rect 14181 22883 14247 22886
rect 16113 22946 16179 22949
rect 20713 22946 20779 22949
rect 16113 22944 20779 22946
rect 16113 22888 16118 22944
rect 16174 22888 20718 22944
rect 20774 22888 20779 22944
rect 16113 22886 20779 22888
rect 16113 22883 16179 22886
rect 20713 22883 20779 22886
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 2773 22810 2839 22813
rect 0 22808 2839 22810
rect 0 22752 2778 22808
rect 2834 22752 2839 22808
rect 0 22750 2839 22752
rect 0 22720 480 22750
rect 2773 22747 2839 22750
rect 11237 22810 11303 22813
rect 14365 22810 14431 22813
rect 27520 22810 28000 22840
rect 11237 22808 14431 22810
rect 11237 22752 11242 22808
rect 11298 22752 14370 22808
rect 14426 22752 14431 22808
rect 11237 22750 14431 22752
rect 11237 22747 11303 22750
rect 14365 22747 14431 22750
rect 24718 22750 28000 22810
rect 1761 22674 1827 22677
rect 5349 22674 5415 22677
rect 1761 22672 5415 22674
rect 1761 22616 1766 22672
rect 1822 22616 5354 22672
rect 5410 22616 5415 22672
rect 1761 22614 5415 22616
rect 1761 22611 1827 22614
rect 5349 22611 5415 22614
rect 9857 22674 9923 22677
rect 12893 22674 12959 22677
rect 9857 22672 12959 22674
rect 9857 22616 9862 22672
rect 9918 22616 12898 22672
rect 12954 22616 12959 22672
rect 9857 22614 12959 22616
rect 9857 22611 9923 22614
rect 12893 22611 12959 22614
rect 13353 22674 13419 22677
rect 15377 22674 15443 22677
rect 13353 22672 15443 22674
rect 13353 22616 13358 22672
rect 13414 22616 15382 22672
rect 15438 22616 15443 22672
rect 13353 22614 15443 22616
rect 13353 22611 13419 22614
rect 15377 22611 15443 22614
rect 16297 22674 16363 22677
rect 19425 22674 19491 22677
rect 19701 22674 19767 22677
rect 16297 22672 19767 22674
rect 16297 22616 16302 22672
rect 16358 22616 19430 22672
rect 19486 22616 19706 22672
rect 19762 22616 19767 22672
rect 16297 22614 19767 22616
rect 16297 22611 16363 22614
rect 19425 22611 19491 22614
rect 19701 22611 19767 22614
rect 23841 22674 23907 22677
rect 24718 22674 24778 22750
rect 27520 22720 28000 22750
rect 23841 22672 24778 22674
rect 23841 22616 23846 22672
rect 23902 22616 24778 22672
rect 23841 22614 24778 22616
rect 23841 22611 23907 22614
rect 2037 22538 2103 22541
rect 10593 22538 10659 22541
rect 2037 22536 10659 22538
rect 2037 22480 2042 22536
rect 2098 22480 10598 22536
rect 10654 22480 10659 22536
rect 2037 22478 10659 22480
rect 2037 22475 2103 22478
rect 10593 22475 10659 22478
rect 10777 22538 10843 22541
rect 12709 22538 12775 22541
rect 10777 22536 12775 22538
rect 10777 22480 10782 22536
rect 10838 22480 12714 22536
rect 12770 22480 12775 22536
rect 10777 22478 12775 22480
rect 10777 22475 10843 22478
rect 12709 22475 12775 22478
rect 14181 22538 14247 22541
rect 16021 22538 16087 22541
rect 23473 22538 23539 22541
rect 14181 22536 16087 22538
rect 14181 22480 14186 22536
rect 14242 22480 16026 22536
rect 16082 22480 16087 22536
rect 14181 22478 16087 22480
rect 14181 22475 14247 22478
rect 16021 22475 16087 22478
rect 17910 22536 23539 22538
rect 17910 22480 23478 22536
rect 23534 22480 23539 22536
rect 17910 22478 23539 22480
rect 2957 22402 3023 22405
rect 3325 22402 3391 22405
rect 7649 22402 7715 22405
rect 17769 22402 17835 22405
rect 2957 22400 7715 22402
rect 2957 22344 2962 22400
rect 3018 22344 3330 22400
rect 3386 22344 7654 22400
rect 7710 22344 7715 22400
rect 2957 22342 7715 22344
rect 2957 22339 3023 22342
rect 3325 22339 3391 22342
rect 7649 22339 7715 22342
rect 13310 22400 17835 22402
rect 13310 22344 17774 22400
rect 17830 22344 17835 22400
rect 13310 22342 17835 22344
rect 10277 22336 10597 22337
rect 0 22266 480 22296
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 1393 22266 1459 22269
rect 0 22264 1459 22266
rect 0 22208 1398 22264
rect 1454 22208 1459 22264
rect 0 22206 1459 22208
rect 0 22176 480 22206
rect 1393 22203 1459 22206
rect 7833 22266 7899 22269
rect 8109 22266 8175 22269
rect 7833 22264 8175 22266
rect 7833 22208 7838 22264
rect 7894 22208 8114 22264
rect 8170 22208 8175 22264
rect 7833 22206 8175 22208
rect 7833 22203 7899 22206
rect 8109 22203 8175 22206
rect 1393 22130 1459 22133
rect 13310 22130 13370 22342
rect 17769 22339 17835 22342
rect 13445 22266 13511 22269
rect 17910 22266 17970 22478
rect 23473 22475 23539 22478
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 13445 22264 17970 22266
rect 13445 22208 13450 22264
rect 13506 22208 17970 22264
rect 13445 22206 17970 22208
rect 24761 22266 24827 22269
rect 27520 22266 28000 22296
rect 24761 22264 28000 22266
rect 24761 22208 24766 22264
rect 24822 22208 28000 22264
rect 24761 22206 28000 22208
rect 13445 22203 13511 22206
rect 24761 22203 24827 22206
rect 27520 22176 28000 22206
rect 14273 22132 14339 22133
rect 1393 22128 13370 22130
rect 1393 22072 1398 22128
rect 1454 22072 13370 22128
rect 1393 22070 13370 22072
rect 1393 22067 1459 22070
rect 14222 22068 14228 22132
rect 14292 22130 14339 22132
rect 15745 22130 15811 22133
rect 19149 22130 19215 22133
rect 20345 22130 20411 22133
rect 14292 22128 14384 22130
rect 14334 22072 14384 22128
rect 14292 22070 14384 22072
rect 15745 22128 20411 22130
rect 15745 22072 15750 22128
rect 15806 22072 19154 22128
rect 19210 22072 20350 22128
rect 20406 22072 20411 22128
rect 15745 22070 20411 22072
rect 14292 22068 14339 22070
rect 14273 22067 14339 22068
rect 15745 22067 15811 22070
rect 19149 22067 19215 22070
rect 20345 22067 20411 22070
rect 21265 22130 21331 22133
rect 24669 22130 24735 22133
rect 21265 22128 24735 22130
rect 21265 22072 21270 22128
rect 21326 22072 24674 22128
rect 24730 22072 24735 22128
rect 21265 22070 24735 22072
rect 21265 22067 21331 22070
rect 24669 22067 24735 22070
rect 7741 21994 7807 21997
rect 10501 21994 10567 21997
rect 7741 21992 10567 21994
rect 7741 21936 7746 21992
rect 7802 21936 10506 21992
rect 10562 21936 10567 21992
rect 7741 21934 10567 21936
rect 7741 21931 7807 21934
rect 10501 21931 10567 21934
rect 14181 21994 14247 21997
rect 25589 21994 25655 21997
rect 14181 21992 25655 21994
rect 14181 21936 14186 21992
rect 14242 21936 25594 21992
rect 25650 21936 25655 21992
rect 14181 21934 25655 21936
rect 14181 21931 14247 21934
rect 25589 21931 25655 21934
rect 7833 21858 7899 21861
rect 14641 21858 14707 21861
rect 7833 21856 14707 21858
rect 7833 21800 7838 21856
rect 7894 21800 14646 21856
rect 14702 21800 14707 21856
rect 7833 21798 14707 21800
rect 7833 21795 7899 21798
rect 14641 21795 14707 21798
rect 19425 21858 19491 21861
rect 21909 21858 21975 21861
rect 19425 21856 21975 21858
rect 19425 21800 19430 21856
rect 19486 21800 21914 21856
rect 21970 21800 21975 21856
rect 19425 21798 21975 21800
rect 19425 21795 19491 21798
rect 21909 21795 21975 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 1761 21722 1827 21725
rect 5349 21722 5415 21725
rect 1761 21720 5415 21722
rect 1761 21664 1766 21720
rect 1822 21664 5354 21720
rect 5410 21664 5415 21720
rect 1761 21662 5415 21664
rect 1761 21659 1827 21662
rect 5349 21659 5415 21662
rect 0 21586 480 21616
rect 1485 21586 1551 21589
rect 0 21584 1551 21586
rect 0 21528 1490 21584
rect 1546 21528 1551 21584
rect 0 21526 1551 21528
rect 0 21496 480 21526
rect 1485 21523 1551 21526
rect 8109 21586 8175 21589
rect 8753 21586 8819 21589
rect 16113 21586 16179 21589
rect 8109 21584 16179 21586
rect 8109 21528 8114 21584
rect 8170 21528 8758 21584
rect 8814 21528 16118 21584
rect 16174 21528 16179 21584
rect 8109 21526 16179 21528
rect 8109 21523 8175 21526
rect 8753 21523 8819 21526
rect 16113 21523 16179 21526
rect 24669 21586 24735 21589
rect 27520 21586 28000 21616
rect 24669 21584 28000 21586
rect 24669 21528 24674 21584
rect 24730 21528 28000 21584
rect 24669 21526 28000 21528
rect 24669 21523 24735 21526
rect 27520 21496 28000 21526
rect 9857 21450 9923 21453
rect 15929 21450 15995 21453
rect 9857 21448 15995 21450
rect 9857 21392 9862 21448
rect 9918 21392 15934 21448
rect 15990 21392 15995 21448
rect 9857 21390 15995 21392
rect 9857 21387 9923 21390
rect 15929 21387 15995 21390
rect 17902 21388 17908 21452
rect 17972 21450 17978 21452
rect 18413 21450 18479 21453
rect 17972 21448 18479 21450
rect 17972 21392 18418 21448
rect 18474 21392 18479 21448
rect 17972 21390 18479 21392
rect 17972 21388 17978 21390
rect 18413 21387 18479 21390
rect 20529 21450 20595 21453
rect 25037 21450 25103 21453
rect 20529 21448 25103 21450
rect 20529 21392 20534 21448
rect 20590 21392 25042 21448
rect 25098 21392 25103 21448
rect 20529 21390 25103 21392
rect 20529 21387 20595 21390
rect 25037 21387 25103 21390
rect 1393 21314 1459 21317
rect 6085 21314 6151 21317
rect 1393 21312 6151 21314
rect 1393 21256 1398 21312
rect 1454 21256 6090 21312
rect 6146 21256 6151 21312
rect 1393 21254 6151 21256
rect 1393 21251 1459 21254
rect 6085 21251 6151 21254
rect 12382 21252 12388 21316
rect 12452 21314 12458 21316
rect 17401 21314 17467 21317
rect 12452 21312 17467 21314
rect 12452 21256 17406 21312
rect 17462 21256 17467 21312
rect 12452 21254 17467 21256
rect 12452 21252 12458 21254
rect 17401 21251 17467 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 1485 21178 1551 21181
rect 4613 21178 4679 21181
rect 1485 21176 4679 21178
rect 1485 21120 1490 21176
rect 1546 21120 4618 21176
rect 4674 21120 4679 21176
rect 1485 21118 4679 21120
rect 1485 21115 1551 21118
rect 4613 21115 4679 21118
rect 7741 21178 7807 21181
rect 10133 21178 10199 21181
rect 7741 21176 10199 21178
rect 7741 21120 7746 21176
rect 7802 21120 10138 21176
rect 10194 21120 10199 21176
rect 7741 21118 10199 21120
rect 7741 21115 7807 21118
rect 10133 21115 10199 21118
rect 10777 21178 10843 21181
rect 14089 21178 14155 21181
rect 10777 21176 14155 21178
rect 10777 21120 10782 21176
rect 10838 21120 14094 21176
rect 14150 21120 14155 21176
rect 10777 21118 14155 21120
rect 10777 21115 10843 21118
rect 14089 21115 14155 21118
rect 14549 21178 14615 21181
rect 17493 21178 17559 21181
rect 18413 21178 18479 21181
rect 14549 21176 18479 21178
rect 14549 21120 14554 21176
rect 14610 21120 17498 21176
rect 17554 21120 18418 21176
rect 18474 21120 18479 21176
rect 14549 21118 18479 21120
rect 14549 21115 14615 21118
rect 17493 21115 17559 21118
rect 18413 21115 18479 21118
rect 0 21042 480 21072
rect 5717 21042 5783 21045
rect 0 21040 5783 21042
rect 0 20984 5722 21040
rect 5778 20984 5783 21040
rect 0 20982 5783 20984
rect 0 20952 480 20982
rect 5717 20979 5783 20982
rect 8661 21042 8727 21045
rect 14089 21042 14155 21045
rect 8661 21040 14155 21042
rect 8661 20984 8666 21040
rect 8722 20984 14094 21040
rect 14150 20984 14155 21040
rect 8661 20982 14155 20984
rect 8661 20979 8727 20982
rect 14089 20979 14155 20982
rect 14273 21042 14339 21045
rect 17033 21042 17099 21045
rect 14273 21040 17099 21042
rect 14273 20984 14278 21040
rect 14334 20984 17038 21040
rect 17094 20984 17099 21040
rect 14273 20982 17099 20984
rect 14273 20979 14339 20982
rect 17033 20979 17099 20982
rect 23790 20980 23796 21044
rect 23860 21042 23866 21044
rect 27520 21042 28000 21072
rect 23860 20982 28000 21042
rect 23860 20980 23866 20982
rect 27520 20952 28000 20982
rect 6177 20906 6243 20909
rect 10041 20906 10107 20909
rect 15377 20906 15443 20909
rect 6177 20904 15443 20906
rect 6177 20848 6182 20904
rect 6238 20848 10046 20904
rect 10102 20848 15382 20904
rect 15438 20848 15443 20904
rect 6177 20846 15443 20848
rect 6177 20843 6243 20846
rect 10041 20843 10107 20846
rect 15377 20843 15443 20846
rect 2221 20770 2287 20773
rect 2497 20770 2563 20773
rect 2630 20770 2636 20772
rect 2221 20768 2636 20770
rect 2221 20712 2226 20768
rect 2282 20712 2502 20768
rect 2558 20712 2636 20768
rect 2221 20710 2636 20712
rect 2221 20707 2287 20710
rect 2497 20707 2563 20710
rect 2630 20708 2636 20710
rect 2700 20708 2706 20772
rect 6729 20770 6795 20773
rect 9213 20770 9279 20773
rect 6729 20768 9279 20770
rect 6729 20712 6734 20768
rect 6790 20712 9218 20768
rect 9274 20712 9279 20768
rect 6729 20710 9279 20712
rect 6729 20707 6795 20710
rect 9213 20707 9279 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10777 20634 10843 20637
rect 14457 20634 14523 20637
rect 10777 20632 14523 20634
rect 10777 20576 10782 20632
rect 10838 20576 14462 20632
rect 14518 20576 14523 20632
rect 10777 20574 14523 20576
rect 10777 20571 10843 20574
rect 14457 20571 14523 20574
rect 15745 20634 15811 20637
rect 19517 20634 19583 20637
rect 21633 20634 21699 20637
rect 15745 20632 21699 20634
rect 15745 20576 15750 20632
rect 15806 20576 19522 20632
rect 19578 20576 21638 20632
rect 21694 20576 21699 20632
rect 15745 20574 21699 20576
rect 15745 20571 15811 20574
rect 19517 20571 19583 20574
rect 21633 20571 21699 20574
rect 7097 20498 7163 20501
rect 12382 20498 12388 20500
rect 7097 20496 12388 20498
rect 7097 20440 7102 20496
rect 7158 20440 12388 20496
rect 7097 20438 12388 20440
rect 7097 20435 7163 20438
rect 12382 20436 12388 20438
rect 12452 20436 12458 20500
rect 20713 20498 20779 20501
rect 12574 20496 20779 20498
rect 12574 20440 20718 20496
rect 20774 20440 20779 20496
rect 12574 20438 20779 20440
rect 0 20362 480 20392
rect 2865 20362 2931 20365
rect 0 20360 2931 20362
rect 0 20304 2870 20360
rect 2926 20304 2931 20360
rect 0 20302 2931 20304
rect 0 20272 480 20302
rect 2865 20299 2931 20302
rect 7557 20362 7623 20365
rect 9397 20362 9463 20365
rect 7557 20360 9463 20362
rect 7557 20304 7562 20360
rect 7618 20304 9402 20360
rect 9458 20304 9463 20360
rect 7557 20302 9463 20304
rect 7557 20299 7623 20302
rect 9397 20299 9463 20302
rect 11329 20362 11395 20365
rect 12574 20362 12634 20438
rect 20713 20435 20779 20438
rect 11329 20360 12634 20362
rect 11329 20304 11334 20360
rect 11390 20304 12634 20360
rect 11329 20302 12634 20304
rect 12985 20362 13051 20365
rect 19333 20362 19399 20365
rect 12985 20360 19399 20362
rect 12985 20304 12990 20360
rect 13046 20304 19338 20360
rect 19394 20304 19399 20360
rect 12985 20302 19399 20304
rect 11329 20299 11395 20302
rect 12985 20299 13051 20302
rect 19333 20299 19399 20302
rect 23657 20362 23723 20365
rect 27520 20362 28000 20392
rect 23657 20360 28000 20362
rect 23657 20304 23662 20360
rect 23718 20304 28000 20360
rect 23657 20302 28000 20304
rect 23657 20299 23723 20302
rect 27520 20272 28000 20302
rect 2037 20226 2103 20229
rect 4613 20226 4679 20229
rect 2037 20224 4679 20226
rect 2037 20168 2042 20224
rect 2098 20168 4618 20224
rect 4674 20168 4679 20224
rect 2037 20166 4679 20168
rect 2037 20163 2103 20166
rect 4613 20163 4679 20166
rect 6637 20226 6703 20229
rect 9489 20226 9555 20229
rect 6637 20224 9555 20226
rect 6637 20168 6642 20224
rect 6698 20168 9494 20224
rect 9550 20168 9555 20224
rect 6637 20166 9555 20168
rect 6637 20163 6703 20166
rect 9489 20163 9555 20166
rect 11053 20226 11119 20229
rect 11973 20226 12039 20229
rect 13997 20226 14063 20229
rect 14273 20228 14339 20229
rect 14222 20226 14228 20228
rect 11053 20224 14063 20226
rect 11053 20168 11058 20224
rect 11114 20168 11978 20224
rect 12034 20168 14002 20224
rect 14058 20168 14063 20224
rect 11053 20166 14063 20168
rect 14182 20166 14228 20226
rect 14292 20224 14339 20228
rect 14334 20168 14339 20224
rect 11053 20163 11119 20166
rect 11973 20163 12039 20166
rect 13997 20163 14063 20166
rect 14222 20164 14228 20166
rect 14292 20164 14339 20168
rect 14273 20163 14339 20164
rect 15285 20226 15351 20229
rect 18505 20226 18571 20229
rect 15285 20224 18571 20226
rect 15285 20168 15290 20224
rect 15346 20168 18510 20224
rect 18566 20168 18571 20224
rect 15285 20166 18571 20168
rect 15285 20163 15351 20166
rect 18505 20163 18571 20166
rect 23013 20226 23079 20229
rect 24209 20226 24275 20229
rect 23013 20224 24275 20226
rect 23013 20168 23018 20224
rect 23074 20168 24214 20224
rect 24270 20168 24275 20224
rect 23013 20166 24275 20168
rect 23013 20163 23079 20166
rect 24209 20163 24275 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 3693 20090 3759 20093
rect 5073 20090 5139 20093
rect 16481 20090 16547 20093
rect 26049 20090 26115 20093
rect 3693 20088 5139 20090
rect 3693 20032 3698 20088
rect 3754 20032 5078 20088
rect 5134 20032 5139 20088
rect 3693 20030 5139 20032
rect 3693 20027 3759 20030
rect 5073 20027 5139 20030
rect 13080 20088 16547 20090
rect 13080 20032 16486 20088
rect 16542 20032 16547 20088
rect 13080 20030 16547 20032
rect 6361 19954 6427 19957
rect 13080 19954 13140 20030
rect 16481 20027 16547 20030
rect 22694 20088 26115 20090
rect 22694 20032 26054 20088
rect 26110 20032 26115 20088
rect 22694 20030 26115 20032
rect 6361 19952 13140 19954
rect 6361 19896 6366 19952
rect 6422 19896 13140 19952
rect 6361 19894 13140 19896
rect 14641 19954 14707 19957
rect 16849 19954 16915 19957
rect 20897 19954 20963 19957
rect 14641 19952 15578 19954
rect 14641 19896 14646 19952
rect 14702 19896 15578 19952
rect 14641 19894 15578 19896
rect 6361 19891 6427 19894
rect 14641 19891 14707 19894
rect 0 19818 480 19848
rect 1577 19818 1643 19821
rect 0 19816 1643 19818
rect 0 19760 1582 19816
rect 1638 19760 1643 19816
rect 0 19758 1643 19760
rect 0 19728 480 19758
rect 1577 19755 1643 19758
rect 2865 19818 2931 19821
rect 4705 19818 4771 19821
rect 2865 19816 15394 19818
rect 2865 19760 2870 19816
rect 2926 19760 4710 19816
rect 4766 19760 15394 19816
rect 2865 19758 15394 19760
rect 2865 19755 2931 19758
rect 4705 19755 4771 19758
rect 9581 19682 9647 19685
rect 11329 19682 11395 19685
rect 9581 19680 11395 19682
rect 9581 19624 9586 19680
rect 9642 19624 11334 19680
rect 11390 19624 11395 19680
rect 9581 19622 11395 19624
rect 9581 19619 9647 19622
rect 11329 19619 11395 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 6913 19546 6979 19549
rect 9949 19546 10015 19549
rect 6913 19544 10015 19546
rect 6913 19488 6918 19544
rect 6974 19488 9954 19544
rect 10010 19488 10015 19544
rect 6913 19486 10015 19488
rect 15334 19546 15394 19758
rect 15518 19682 15578 19894
rect 16849 19952 20963 19954
rect 16849 19896 16854 19952
rect 16910 19896 20902 19952
rect 20958 19896 20963 19952
rect 16849 19894 20963 19896
rect 16849 19891 16915 19894
rect 20897 19891 20963 19894
rect 19149 19818 19215 19821
rect 22461 19818 22527 19821
rect 19149 19816 22527 19818
rect 19149 19760 19154 19816
rect 19210 19760 22466 19816
rect 22522 19760 22527 19816
rect 19149 19758 22527 19760
rect 19149 19755 19215 19758
rect 22461 19755 22527 19758
rect 20345 19682 20411 19685
rect 15518 19680 20411 19682
rect 15518 19624 20350 19680
rect 20406 19624 20411 19680
rect 15518 19622 20411 19624
rect 20345 19619 20411 19622
rect 22694 19546 22754 20030
rect 26049 20027 26115 20030
rect 23381 19954 23447 19957
rect 23381 19952 25330 19954
rect 23381 19896 23386 19952
rect 23442 19896 25330 19952
rect 23381 19894 25330 19896
rect 23381 19891 23447 19894
rect 22829 19818 22895 19821
rect 25129 19818 25195 19821
rect 22829 19816 25195 19818
rect 22829 19760 22834 19816
rect 22890 19760 25134 19816
rect 25190 19760 25195 19816
rect 22829 19758 25195 19760
rect 25270 19818 25330 19894
rect 27520 19818 28000 19848
rect 25270 19758 28000 19818
rect 22829 19755 22895 19758
rect 25129 19755 25195 19758
rect 27520 19728 28000 19758
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 15334 19486 22754 19546
rect 6913 19483 6979 19486
rect 9949 19483 10015 19486
rect 4889 19410 4955 19413
rect 12617 19410 12683 19413
rect 4889 19408 12683 19410
rect 4889 19352 4894 19408
rect 4950 19352 12622 19408
rect 12678 19352 12683 19408
rect 4889 19350 12683 19352
rect 4889 19347 4955 19350
rect 12617 19347 12683 19350
rect 13077 19410 13143 19413
rect 15653 19410 15719 19413
rect 13077 19408 15719 19410
rect 13077 19352 13082 19408
rect 13138 19352 15658 19408
rect 15714 19352 15719 19408
rect 13077 19350 15719 19352
rect 13077 19347 13143 19350
rect 15653 19347 15719 19350
rect 18229 19410 18295 19413
rect 19701 19410 19767 19413
rect 18229 19408 19767 19410
rect 18229 19352 18234 19408
rect 18290 19352 19706 19408
rect 19762 19352 19767 19408
rect 18229 19350 19767 19352
rect 18229 19347 18295 19350
rect 19701 19347 19767 19350
rect 24025 19410 24091 19413
rect 25405 19410 25471 19413
rect 24025 19408 25471 19410
rect 24025 19352 24030 19408
rect 24086 19352 25410 19408
rect 25466 19352 25471 19408
rect 24025 19350 25471 19352
rect 24025 19347 24091 19350
rect 25405 19347 25471 19350
rect 8661 19274 8727 19277
rect 14365 19274 14431 19277
rect 8661 19272 14431 19274
rect 8661 19216 8666 19272
rect 8722 19216 14370 19272
rect 14426 19216 14431 19272
rect 8661 19214 14431 19216
rect 8661 19211 8727 19214
rect 14365 19211 14431 19214
rect 18505 19274 18571 19277
rect 22277 19274 22343 19277
rect 18505 19272 22343 19274
rect 18505 19216 18510 19272
rect 18566 19216 22282 19272
rect 22338 19216 22343 19272
rect 18505 19214 22343 19216
rect 18505 19211 18571 19214
rect 22277 19211 22343 19214
rect 0 19138 480 19168
rect 3969 19138 4035 19141
rect 0 19136 4035 19138
rect 0 19080 3974 19136
rect 4030 19080 4035 19136
rect 0 19078 4035 19080
rect 0 19048 480 19078
rect 3969 19075 4035 19078
rect 10685 19138 10751 19141
rect 15469 19138 15535 19141
rect 10685 19136 15535 19138
rect 10685 19080 10690 19136
rect 10746 19080 15474 19136
rect 15530 19080 15535 19136
rect 10685 19078 15535 19080
rect 10685 19075 10751 19078
rect 15469 19075 15535 19078
rect 21725 19138 21791 19141
rect 27520 19138 28000 19168
rect 21725 19136 28000 19138
rect 21725 19080 21730 19136
rect 21786 19080 28000 19136
rect 21725 19078 28000 19080
rect 21725 19075 21791 19078
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 27520 19048 28000 19078
rect 19610 19007 19930 19008
rect 2497 19002 2563 19005
rect 6361 19002 6427 19005
rect 6913 19002 6979 19005
rect 2497 19000 6979 19002
rect 2497 18944 2502 19000
rect 2558 18944 6366 19000
rect 6422 18944 6918 19000
rect 6974 18944 6979 19000
rect 2497 18942 6979 18944
rect 2497 18939 2563 18942
rect 6361 18939 6427 18942
rect 6913 18939 6979 18942
rect 10777 19002 10843 19005
rect 15009 19002 15075 19005
rect 17769 19002 17835 19005
rect 10777 19000 15075 19002
rect 10777 18944 10782 19000
rect 10838 18944 15014 19000
rect 15070 18944 15075 19000
rect 10777 18942 15075 18944
rect 10777 18939 10843 18942
rect 15009 18939 15075 18942
rect 16254 19000 17835 19002
rect 16254 18944 17774 19000
rect 17830 18944 17835 19000
rect 16254 18942 17835 18944
rect 1853 18866 1919 18869
rect 16254 18866 16314 18942
rect 17769 18939 17835 18942
rect 21541 19002 21607 19005
rect 21909 19002 21975 19005
rect 25037 19002 25103 19005
rect 21541 19000 25103 19002
rect 21541 18944 21546 19000
rect 21602 18944 21914 19000
rect 21970 18944 25042 19000
rect 25098 18944 25103 19000
rect 21541 18942 25103 18944
rect 21541 18939 21607 18942
rect 21909 18939 21975 18942
rect 25037 18939 25103 18942
rect 1853 18864 16314 18866
rect 1853 18808 1858 18864
rect 1914 18808 16314 18864
rect 1853 18806 16314 18808
rect 16481 18866 16547 18869
rect 24117 18866 24183 18869
rect 16481 18864 24183 18866
rect 16481 18808 16486 18864
rect 16542 18808 24122 18864
rect 24178 18808 24183 18864
rect 16481 18806 24183 18808
rect 1853 18803 1919 18806
rect 12344 18772 12450 18806
rect 16481 18803 16547 18806
rect 24117 18803 24183 18806
rect 2405 18730 2471 18733
rect 7741 18730 7807 18733
rect 11973 18730 12039 18733
rect 2405 18728 7666 18730
rect 2405 18672 2410 18728
rect 2466 18672 7666 18728
rect 2405 18670 7666 18672
rect 2405 18667 2471 18670
rect 0 18594 480 18624
rect 5441 18594 5507 18597
rect 0 18592 5507 18594
rect 0 18536 5446 18592
rect 5502 18536 5507 18592
rect 0 18534 5507 18536
rect 7606 18594 7666 18670
rect 7741 18728 12039 18730
rect 7741 18672 7746 18728
rect 7802 18672 11978 18728
rect 12034 18672 12039 18728
rect 7741 18670 12039 18672
rect 7741 18667 7807 18670
rect 11973 18667 12039 18670
rect 18413 18730 18479 18733
rect 20989 18730 21055 18733
rect 23473 18730 23539 18733
rect 18413 18728 23539 18730
rect 18413 18672 18418 18728
rect 18474 18672 20994 18728
rect 21050 18672 23478 18728
rect 23534 18672 23539 18728
rect 18413 18670 23539 18672
rect 18413 18667 18479 18670
rect 20989 18667 21055 18670
rect 23473 18667 23539 18670
rect 24894 18668 24900 18732
rect 24964 18730 24970 18732
rect 25589 18730 25655 18733
rect 24964 18728 25655 18730
rect 24964 18672 25594 18728
rect 25650 18672 25655 18728
rect 24964 18670 25655 18672
rect 24964 18668 24970 18670
rect 25589 18667 25655 18670
rect 22093 18594 22159 18597
rect 23381 18594 23447 18597
rect 27520 18594 28000 18624
rect 7606 18534 10794 18594
rect 0 18504 480 18534
rect 5441 18531 5507 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 6821 18458 6887 18461
rect 10593 18458 10659 18461
rect 6821 18456 10659 18458
rect 6821 18400 6826 18456
rect 6882 18400 10598 18456
rect 10654 18400 10659 18456
rect 6821 18398 10659 18400
rect 6821 18395 6887 18398
rect 10593 18395 10659 18398
rect 5717 18186 5783 18189
rect 8477 18186 8543 18189
rect 5717 18184 8543 18186
rect 5717 18128 5722 18184
rect 5778 18128 8482 18184
rect 8538 18128 8543 18184
rect 5717 18126 8543 18128
rect 5717 18123 5783 18126
rect 8477 18123 8543 18126
rect 3233 18050 3299 18053
rect 6821 18050 6887 18053
rect 3233 18048 6887 18050
rect 3233 17992 3238 18048
rect 3294 17992 6826 18048
rect 6882 17992 6887 18048
rect 3233 17990 6887 17992
rect 10734 18050 10794 18534
rect 22093 18592 23447 18594
rect 22093 18536 22098 18592
rect 22154 18536 23386 18592
rect 23442 18536 23447 18592
rect 22093 18534 23447 18536
rect 22093 18531 22159 18534
rect 23381 18531 23447 18534
rect 24902 18534 28000 18594
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 13486 18396 13492 18460
rect 13556 18458 13562 18460
rect 14089 18458 14155 18461
rect 13556 18456 14155 18458
rect 13556 18400 14094 18456
rect 14150 18400 14155 18456
rect 13556 18398 14155 18400
rect 13556 18396 13562 18398
rect 14089 18395 14155 18398
rect 18781 18458 18847 18461
rect 22645 18458 22711 18461
rect 18781 18456 22711 18458
rect 18781 18400 18786 18456
rect 18842 18400 22650 18456
rect 22706 18400 22711 18456
rect 18781 18398 22711 18400
rect 18781 18395 18847 18398
rect 22645 18395 22711 18398
rect 11881 18322 11947 18325
rect 19425 18322 19491 18325
rect 11881 18320 19491 18322
rect 11881 18264 11886 18320
rect 11942 18264 19430 18320
rect 19486 18264 19491 18320
rect 11881 18262 19491 18264
rect 11881 18259 11947 18262
rect 19425 18259 19491 18262
rect 11421 18186 11487 18189
rect 24902 18186 24962 18534
rect 27520 18504 28000 18534
rect 11421 18184 24962 18186
rect 11421 18128 11426 18184
rect 11482 18128 24962 18184
rect 11421 18126 24962 18128
rect 11421 18123 11487 18126
rect 17125 18050 17191 18053
rect 10734 18048 17191 18050
rect 10734 17992 17130 18048
rect 17186 17992 17191 18048
rect 10734 17990 17191 17992
rect 3233 17987 3299 17990
rect 6821 17987 6887 17990
rect 17125 17987 17191 17990
rect 17309 18050 17375 18053
rect 19333 18050 19399 18053
rect 17309 18048 19399 18050
rect 17309 17992 17314 18048
rect 17370 17992 19338 18048
rect 19394 17992 19399 18048
rect 17309 17990 19399 17992
rect 17309 17987 17375 17990
rect 19333 17987 19399 17990
rect 22277 18050 22343 18053
rect 25681 18050 25747 18053
rect 22277 18048 25747 18050
rect 22277 17992 22282 18048
rect 22338 17992 25686 18048
rect 25742 17992 25747 18048
rect 22277 17990 25747 17992
rect 22277 17987 22343 17990
rect 25681 17987 25747 17990
rect 10277 17984 10597 17985
rect 0 17914 480 17944
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3785 17914 3851 17917
rect 0 17912 3851 17914
rect 0 17856 3790 17912
rect 3846 17856 3851 17912
rect 0 17854 3851 17856
rect 0 17824 480 17854
rect 3785 17851 3851 17854
rect 11789 17914 11855 17917
rect 14641 17914 14707 17917
rect 11789 17912 14707 17914
rect 11789 17856 11794 17912
rect 11850 17856 14646 17912
rect 14702 17856 14707 17912
rect 11789 17854 14707 17856
rect 11789 17851 11855 17854
rect 14641 17851 14707 17854
rect 25773 17914 25839 17917
rect 27520 17914 28000 17944
rect 25773 17912 28000 17914
rect 25773 17856 25778 17912
rect 25834 17856 28000 17912
rect 25773 17854 28000 17856
rect 25773 17851 25839 17854
rect 27520 17824 28000 17854
rect 1669 17778 1735 17781
rect 6177 17778 6243 17781
rect 1669 17776 6243 17778
rect 1669 17720 1674 17776
rect 1730 17720 6182 17776
rect 6238 17720 6243 17776
rect 1669 17718 6243 17720
rect 1669 17715 1735 17718
rect 6177 17715 6243 17718
rect 8017 17778 8083 17781
rect 14457 17778 14523 17781
rect 8017 17776 14523 17778
rect 8017 17720 8022 17776
rect 8078 17720 14462 17776
rect 14518 17720 14523 17776
rect 8017 17718 14523 17720
rect 8017 17715 8083 17718
rect 14457 17715 14523 17718
rect 17033 17778 17099 17781
rect 19241 17778 19307 17781
rect 22277 17778 22343 17781
rect 17033 17776 22343 17778
rect 17033 17720 17038 17776
rect 17094 17720 19246 17776
rect 19302 17720 22282 17776
rect 22338 17720 22343 17776
rect 17033 17718 22343 17720
rect 17033 17715 17099 17718
rect 19241 17715 19307 17718
rect 22277 17715 22343 17718
rect 2221 17642 2287 17645
rect 6085 17642 6151 17645
rect 2221 17640 6151 17642
rect 2221 17584 2226 17640
rect 2282 17584 6090 17640
rect 6146 17584 6151 17640
rect 2221 17582 6151 17584
rect 2221 17579 2287 17582
rect 6085 17579 6151 17582
rect 6269 17642 6335 17645
rect 14917 17642 14983 17645
rect 6269 17640 14983 17642
rect 6269 17584 6274 17640
rect 6330 17584 14922 17640
rect 14978 17584 14983 17640
rect 6269 17582 14983 17584
rect 6269 17579 6335 17582
rect 14917 17579 14983 17582
rect 15101 17642 15167 17645
rect 17769 17642 17835 17645
rect 15101 17640 17835 17642
rect 15101 17584 15106 17640
rect 15162 17584 17774 17640
rect 17830 17584 17835 17640
rect 15101 17582 17835 17584
rect 15101 17579 15167 17582
rect 17769 17579 17835 17582
rect 21633 17642 21699 17645
rect 24710 17642 24716 17644
rect 21633 17640 24716 17642
rect 21633 17584 21638 17640
rect 21694 17584 24716 17640
rect 21633 17582 24716 17584
rect 21633 17579 21699 17582
rect 24710 17580 24716 17582
rect 24780 17580 24786 17644
rect 9673 17506 9739 17509
rect 13997 17506 14063 17509
rect 9673 17504 14063 17506
rect 9673 17448 9678 17504
rect 9734 17448 14002 17504
rect 14058 17448 14063 17504
rect 9673 17446 14063 17448
rect 9673 17443 9739 17446
rect 13997 17443 14063 17446
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 7557 17370 7623 17373
rect 13813 17370 13879 17373
rect 0 17310 5136 17370
rect 0 17280 480 17310
rect 5076 17234 5136 17310
rect 7557 17368 13879 17370
rect 7557 17312 7562 17368
rect 7618 17312 13818 17368
rect 13874 17312 13879 17368
rect 7557 17310 13879 17312
rect 7557 17307 7623 17310
rect 13813 17307 13879 17310
rect 26141 17370 26207 17373
rect 27520 17370 28000 17400
rect 26141 17368 28000 17370
rect 26141 17312 26146 17368
rect 26202 17312 28000 17368
rect 26141 17310 28000 17312
rect 26141 17307 26207 17310
rect 27520 17280 28000 17310
rect 7005 17234 7071 17237
rect 5076 17232 7071 17234
rect 5076 17176 7010 17232
rect 7066 17176 7071 17232
rect 5076 17174 7071 17176
rect 7005 17171 7071 17174
rect 7925 17234 7991 17237
rect 8753 17234 8819 17237
rect 14917 17234 14983 17237
rect 7925 17232 14983 17234
rect 7925 17176 7930 17232
rect 7986 17176 8758 17232
rect 8814 17176 14922 17232
rect 14978 17176 14983 17232
rect 7925 17174 14983 17176
rect 7925 17171 7991 17174
rect 8753 17171 8819 17174
rect 14917 17171 14983 17174
rect 3509 17098 3575 17101
rect 6729 17098 6795 17101
rect 11145 17098 11211 17101
rect 3509 17096 6795 17098
rect 3509 17040 3514 17096
rect 3570 17040 6734 17096
rect 6790 17040 6795 17096
rect 3509 17038 6795 17040
rect 3509 17035 3575 17038
rect 6729 17035 6795 17038
rect 10136 17096 11211 17098
rect 10136 17040 11150 17096
rect 11206 17040 11211 17096
rect 10136 17038 11211 17040
rect 10136 16965 10196 17038
rect 11145 17035 11211 17038
rect 5533 16962 5599 16965
rect 10133 16962 10199 16965
rect 5533 16960 10199 16962
rect 5533 16904 5538 16960
rect 5594 16904 10138 16960
rect 10194 16904 10199 16960
rect 5533 16902 10199 16904
rect 5533 16899 5599 16902
rect 10133 16899 10199 16902
rect 23013 16962 23079 16965
rect 23013 16960 25514 16962
rect 23013 16904 23018 16960
rect 23074 16904 25514 16960
rect 23013 16902 25514 16904
rect 23013 16899 23079 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 5349 16826 5415 16829
rect 8017 16826 8083 16829
rect 8569 16826 8635 16829
rect 10133 16826 10199 16829
rect 5349 16824 10199 16826
rect 5349 16768 5354 16824
rect 5410 16768 8022 16824
rect 8078 16768 8574 16824
rect 8630 16768 10138 16824
rect 10194 16768 10199 16824
rect 5349 16766 10199 16768
rect 5349 16763 5415 16766
rect 8017 16763 8083 16766
rect 8569 16763 8635 16766
rect 10133 16763 10199 16766
rect 22921 16826 22987 16829
rect 25129 16826 25195 16829
rect 22921 16824 25195 16826
rect 22921 16768 22926 16824
rect 22982 16768 25134 16824
rect 25190 16768 25195 16824
rect 22921 16766 25195 16768
rect 22921 16763 22987 16766
rect 25129 16763 25195 16766
rect 0 16690 480 16720
rect 3141 16690 3207 16693
rect 9581 16690 9647 16693
rect 0 16630 1410 16690
rect 0 16600 480 16630
rect 1350 16554 1410 16630
rect 3141 16688 9647 16690
rect 3141 16632 3146 16688
rect 3202 16632 9586 16688
rect 9642 16632 9647 16688
rect 3141 16630 9647 16632
rect 3141 16627 3207 16630
rect 9581 16627 9647 16630
rect 13261 16690 13327 16693
rect 15469 16690 15535 16693
rect 13261 16688 15535 16690
rect 13261 16632 13266 16688
rect 13322 16632 15474 16688
rect 15530 16632 15535 16688
rect 13261 16630 15535 16632
rect 13261 16627 13327 16630
rect 15469 16627 15535 16630
rect 20805 16690 20871 16693
rect 22461 16690 22527 16693
rect 25221 16690 25287 16693
rect 20805 16688 20914 16690
rect 20805 16632 20810 16688
rect 20866 16632 20914 16688
rect 20805 16627 20914 16632
rect 22461 16688 25287 16690
rect 22461 16632 22466 16688
rect 22522 16632 25226 16688
rect 25282 16632 25287 16688
rect 22461 16630 25287 16632
rect 25454 16690 25514 16902
rect 27520 16690 28000 16720
rect 25454 16630 28000 16690
rect 22461 16627 22527 16630
rect 25221 16627 25287 16630
rect 1485 16554 1551 16557
rect 1350 16552 1551 16554
rect 1350 16496 1490 16552
rect 1546 16496 1551 16552
rect 1350 16494 1551 16496
rect 1485 16491 1551 16494
rect 7833 16554 7899 16557
rect 14457 16554 14523 16557
rect 15377 16554 15443 16557
rect 7833 16552 14336 16554
rect 7833 16496 7838 16552
rect 7894 16496 14336 16552
rect 7833 16494 14336 16496
rect 7833 16491 7899 16494
rect 8937 16418 9003 16421
rect 13905 16418 13971 16421
rect 8937 16416 13971 16418
rect 8937 16360 8942 16416
rect 8998 16360 13910 16416
rect 13966 16360 13971 16416
rect 8937 16358 13971 16360
rect 8937 16355 9003 16358
rect 13905 16355 13971 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 6637 16282 6703 16285
rect 9213 16282 9279 16285
rect 6637 16280 9279 16282
rect 6637 16224 6642 16280
rect 6698 16224 9218 16280
rect 9274 16224 9279 16280
rect 6637 16222 9279 16224
rect 6637 16219 6703 16222
rect 9213 16219 9279 16222
rect 10777 16282 10843 16285
rect 13997 16282 14063 16285
rect 10777 16280 14063 16282
rect 10777 16224 10782 16280
rect 10838 16224 14002 16280
rect 14058 16224 14063 16280
rect 10777 16222 14063 16224
rect 10777 16219 10843 16222
rect 13997 16219 14063 16222
rect 0 16146 480 16176
rect 4061 16146 4127 16149
rect 0 16144 4127 16146
rect 0 16088 4066 16144
rect 4122 16088 4127 16144
rect 0 16086 4127 16088
rect 0 16056 480 16086
rect 4061 16083 4127 16086
rect 10961 16146 11027 16149
rect 12801 16146 12867 16149
rect 10961 16144 12867 16146
rect 10961 16088 10966 16144
rect 11022 16088 12806 16144
rect 12862 16088 12867 16144
rect 10961 16086 12867 16088
rect 14276 16146 14336 16494
rect 14457 16552 15443 16554
rect 14457 16496 14462 16552
rect 14518 16496 15382 16552
rect 15438 16496 15443 16552
rect 14457 16494 15443 16496
rect 14457 16491 14523 16494
rect 15377 16491 15443 16494
rect 16481 16554 16547 16557
rect 18505 16554 18571 16557
rect 16481 16552 18571 16554
rect 16481 16496 16486 16552
rect 16542 16496 18510 16552
rect 18566 16496 18571 16552
rect 16481 16494 18571 16496
rect 16481 16491 16547 16494
rect 18505 16491 18571 16494
rect 16665 16418 16731 16421
rect 20854 16418 20914 16627
rect 27520 16600 28000 16630
rect 24669 16554 24735 16557
rect 25129 16554 25195 16557
rect 24669 16552 25195 16554
rect 24669 16496 24674 16552
rect 24730 16496 25134 16552
rect 25190 16496 25195 16552
rect 24669 16494 25195 16496
rect 24669 16491 24735 16494
rect 25129 16491 25195 16494
rect 23606 16418 23612 16420
rect 16665 16416 23612 16418
rect 16665 16360 16670 16416
rect 16726 16360 23612 16416
rect 16665 16358 23612 16360
rect 16665 16355 16731 16358
rect 23606 16356 23612 16358
rect 23676 16356 23682 16420
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 20897 16146 20963 16149
rect 14276 16144 20963 16146
rect 14276 16088 20902 16144
rect 20958 16088 20963 16144
rect 14276 16086 20963 16088
rect 10961 16083 11027 16086
rect 12801 16083 12867 16086
rect 20897 16083 20963 16086
rect 23749 16146 23815 16149
rect 27520 16146 28000 16176
rect 23749 16144 28000 16146
rect 23749 16088 23754 16144
rect 23810 16088 28000 16144
rect 23749 16086 28000 16088
rect 23749 16083 23815 16086
rect 27520 16056 28000 16086
rect 9857 16010 9923 16013
rect 12433 16010 12499 16013
rect 9857 16008 12499 16010
rect 9857 15952 9862 16008
rect 9918 15952 12438 16008
rect 12494 15952 12499 16008
rect 9857 15950 12499 15952
rect 9857 15947 9923 15950
rect 12433 15947 12499 15950
rect 13905 16010 13971 16013
rect 16665 16010 16731 16013
rect 13905 16008 16731 16010
rect 13905 15952 13910 16008
rect 13966 15952 16670 16008
rect 16726 15952 16731 16008
rect 13905 15950 16731 15952
rect 13905 15947 13971 15950
rect 16665 15947 16731 15950
rect 16849 16010 16915 16013
rect 19977 16010 20043 16013
rect 16849 16008 20043 16010
rect 16849 15952 16854 16008
rect 16910 15952 19982 16008
rect 20038 15952 20043 16008
rect 16849 15950 20043 15952
rect 16849 15947 16915 15950
rect 19977 15947 20043 15950
rect 20253 16010 20319 16013
rect 23473 16010 23539 16013
rect 20253 16008 23539 16010
rect 20253 15952 20258 16008
rect 20314 15952 23478 16008
rect 23534 15952 23539 16008
rect 20253 15950 23539 15952
rect 20253 15947 20319 15950
rect 23473 15947 23539 15950
rect 3509 15874 3575 15877
rect 4981 15874 5047 15877
rect 3509 15872 5047 15874
rect 3509 15816 3514 15872
rect 3570 15816 4986 15872
rect 5042 15816 5047 15872
rect 3509 15814 5047 15816
rect 3509 15811 3575 15814
rect 4981 15811 5047 15814
rect 14457 15874 14523 15877
rect 16849 15874 16915 15877
rect 14457 15872 16915 15874
rect 14457 15816 14462 15872
rect 14518 15816 16854 15872
rect 16910 15816 16915 15872
rect 14457 15814 16915 15816
rect 14457 15811 14523 15814
rect 16849 15811 16915 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 13169 15738 13235 15741
rect 13302 15738 13308 15740
rect 13169 15736 13308 15738
rect 13169 15680 13174 15736
rect 13230 15680 13308 15736
rect 13169 15678 13308 15680
rect 13169 15675 13235 15678
rect 13302 15676 13308 15678
rect 13372 15738 13378 15740
rect 13372 15678 19442 15738
rect 13372 15676 13378 15678
rect 1577 15602 1643 15605
rect 6637 15602 6703 15605
rect 1577 15600 6703 15602
rect 1577 15544 1582 15600
rect 1638 15544 6642 15600
rect 6698 15544 6703 15600
rect 1577 15542 6703 15544
rect 1577 15539 1643 15542
rect 6637 15539 6703 15542
rect 9489 15602 9555 15605
rect 11145 15602 11211 15605
rect 9489 15600 11211 15602
rect 9489 15544 9494 15600
rect 9550 15544 11150 15600
rect 11206 15544 11211 15600
rect 9489 15542 11211 15544
rect 9489 15539 9555 15542
rect 11145 15539 11211 15542
rect 12985 15602 13051 15605
rect 19382 15602 19442 15678
rect 20253 15602 20319 15605
rect 12985 15600 16866 15602
rect 12985 15544 12990 15600
rect 13046 15544 16866 15600
rect 12985 15542 16866 15544
rect 19382 15600 20319 15602
rect 19382 15544 20258 15600
rect 20314 15544 20319 15600
rect 19382 15542 20319 15544
rect 12985 15539 13051 15542
rect 0 15466 480 15496
rect 3693 15466 3759 15469
rect 0 15464 3759 15466
rect 0 15408 3698 15464
rect 3754 15408 3759 15464
rect 0 15406 3759 15408
rect 0 15376 480 15406
rect 3693 15403 3759 15406
rect 3969 15466 4035 15469
rect 4613 15466 4679 15469
rect 5257 15466 5323 15469
rect 16573 15466 16639 15469
rect 3969 15464 16639 15466
rect 3969 15408 3974 15464
rect 4030 15408 4618 15464
rect 4674 15408 5262 15464
rect 5318 15408 16578 15464
rect 16634 15408 16639 15464
rect 3969 15406 16639 15408
rect 3969 15403 4035 15406
rect 4613 15403 4679 15406
rect 5257 15403 5323 15406
rect 16573 15403 16639 15406
rect 8569 15330 8635 15333
rect 10041 15330 10107 15333
rect 8569 15328 10107 15330
rect 8569 15272 8574 15328
rect 8630 15272 10046 15328
rect 10102 15272 10107 15328
rect 8569 15270 10107 15272
rect 16806 15330 16866 15542
rect 20253 15539 20319 15542
rect 17769 15466 17835 15469
rect 22645 15466 22711 15469
rect 17769 15464 22711 15466
rect 17769 15408 17774 15464
rect 17830 15408 22650 15464
rect 22706 15408 22711 15464
rect 17769 15406 22711 15408
rect 17769 15403 17835 15406
rect 22645 15403 22711 15406
rect 23841 15466 23907 15469
rect 24669 15466 24735 15469
rect 27520 15466 28000 15496
rect 23841 15464 24042 15466
rect 23841 15408 23846 15464
rect 23902 15408 24042 15464
rect 23841 15406 24042 15408
rect 23841 15403 23907 15406
rect 20621 15330 20687 15333
rect 16806 15328 20687 15330
rect 16806 15272 20626 15328
rect 20682 15272 20687 15328
rect 16806 15270 20687 15272
rect 8569 15267 8635 15270
rect 10041 15267 10107 15270
rect 20621 15267 20687 15270
rect 22001 15330 22067 15333
rect 23841 15330 23907 15333
rect 22001 15328 23907 15330
rect 22001 15272 22006 15328
rect 22062 15272 23846 15328
rect 23902 15272 23907 15328
rect 22001 15270 23907 15272
rect 22001 15267 22067 15270
rect 23841 15267 23907 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 14641 15194 14707 15197
rect 17861 15194 17927 15197
rect 18689 15194 18755 15197
rect 21449 15194 21515 15197
rect 12390 15192 14707 15194
rect 12390 15160 14646 15192
rect 12344 15136 14646 15160
rect 14702 15136 14707 15192
rect 12344 15134 14707 15136
rect 12344 15100 12450 15134
rect 14641 15131 14707 15134
rect 15334 15192 21515 15194
rect 15334 15136 17866 15192
rect 17922 15136 18694 15192
rect 18750 15136 21454 15192
rect 21510 15136 21515 15192
rect 15334 15134 21515 15136
rect 749 15058 815 15061
rect 12344 15058 12404 15100
rect 749 15056 12404 15058
rect 749 15000 754 15056
rect 810 15000 12404 15056
rect 749 14998 12404 15000
rect 13721 15058 13787 15061
rect 15334 15058 15394 15134
rect 17861 15131 17927 15134
rect 18689 15131 18755 15134
rect 21449 15131 21515 15134
rect 22553 15058 22619 15061
rect 13721 15056 15394 15058
rect 13721 15000 13726 15056
rect 13782 15000 15394 15056
rect 13721 14998 15394 15000
rect 17174 15056 22619 15058
rect 17174 15000 22558 15056
rect 22614 15000 22619 15056
rect 17174 14998 22619 15000
rect 749 14995 815 14998
rect 13721 14995 13787 14998
rect 0 14922 480 14952
rect 3141 14922 3207 14925
rect 0 14920 3207 14922
rect 0 14864 3146 14920
rect 3202 14864 3207 14920
rect 0 14862 3207 14864
rect 0 14832 480 14862
rect 3141 14859 3207 14862
rect 3785 14922 3851 14925
rect 5809 14922 5875 14925
rect 3785 14920 5875 14922
rect 3785 14864 3790 14920
rect 3846 14864 5814 14920
rect 5870 14864 5875 14920
rect 3785 14862 5875 14864
rect 3785 14859 3851 14862
rect 5809 14859 5875 14862
rect 7189 14922 7255 14925
rect 17174 14922 17234 14998
rect 22553 14995 22619 14998
rect 7189 14920 17234 14922
rect 7189 14864 7194 14920
rect 7250 14864 17234 14920
rect 7189 14862 17234 14864
rect 17309 14922 17375 14925
rect 23381 14922 23447 14925
rect 17309 14920 23447 14922
rect 17309 14864 17314 14920
rect 17370 14864 23386 14920
rect 23442 14864 23447 14920
rect 17309 14862 23447 14864
rect 23982 14922 24042 15406
rect 24669 15464 28000 15466
rect 24669 15408 24674 15464
rect 24730 15408 28000 15464
rect 24669 15406 28000 15408
rect 24669 15403 24735 15406
rect 27520 15376 28000 15406
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 24853 15194 24919 15197
rect 25957 15194 26023 15197
rect 24853 15192 26023 15194
rect 24853 15136 24858 15192
rect 24914 15136 25962 15192
rect 26018 15136 26023 15192
rect 24853 15134 26023 15136
rect 24853 15131 24919 15134
rect 25957 15131 26023 15134
rect 27520 14922 28000 14952
rect 23982 14862 28000 14922
rect 7189 14859 7255 14862
rect 17309 14859 17375 14862
rect 23381 14859 23447 14862
rect 27520 14832 28000 14862
rect 10685 14786 10751 14789
rect 12801 14786 12867 14789
rect 10685 14784 12867 14786
rect 10685 14728 10690 14784
rect 10746 14728 12806 14784
rect 12862 14728 12867 14784
rect 10685 14726 12867 14728
rect 10685 14723 10751 14726
rect 12801 14723 12867 14726
rect 23422 14724 23428 14788
rect 23492 14786 23498 14788
rect 25037 14786 25103 14789
rect 23492 14784 25103 14786
rect 23492 14728 25042 14784
rect 25098 14728 25103 14784
rect 23492 14726 25103 14728
rect 23492 14724 23498 14726
rect 25037 14723 25103 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1577 14650 1643 14653
rect 4613 14650 4679 14653
rect 1577 14648 4679 14650
rect 1577 14592 1582 14648
rect 1638 14592 4618 14648
rect 4674 14592 4679 14648
rect 1577 14590 4679 14592
rect 1577 14587 1643 14590
rect 4613 14587 4679 14590
rect 12934 14588 12940 14652
rect 13004 14650 13010 14652
rect 13445 14650 13511 14653
rect 13004 14648 13511 14650
rect 13004 14592 13450 14648
rect 13506 14592 13511 14648
rect 13004 14590 13511 14592
rect 13004 14588 13010 14590
rect 13445 14587 13511 14590
rect 2589 14514 2655 14517
rect 10133 14514 10199 14517
rect 14089 14514 14155 14517
rect 2589 14512 4124 14514
rect 2589 14456 2594 14512
rect 2650 14456 4124 14512
rect 2589 14454 4124 14456
rect 2589 14451 2655 14454
rect 0 14378 480 14408
rect 3918 14378 3924 14380
rect 0 14318 3924 14378
rect 0 14288 480 14318
rect 3918 14316 3924 14318
rect 3988 14316 3994 14380
rect 4064 14378 4124 14454
rect 10133 14512 14155 14514
rect 10133 14456 10138 14512
rect 10194 14456 14094 14512
rect 14150 14456 14155 14512
rect 10133 14454 14155 14456
rect 10133 14451 10199 14454
rect 14089 14451 14155 14454
rect 21541 14514 21607 14517
rect 23749 14514 23815 14517
rect 21541 14512 23815 14514
rect 21541 14456 21546 14512
rect 21602 14456 23754 14512
rect 23810 14456 23815 14512
rect 21541 14454 23815 14456
rect 21541 14451 21607 14454
rect 23749 14451 23815 14454
rect 23565 14378 23631 14381
rect 4064 14376 23631 14378
rect 4064 14320 23570 14376
rect 23626 14320 23631 14376
rect 4064 14318 23631 14320
rect 23565 14315 23631 14318
rect 26049 14378 26115 14381
rect 27520 14378 28000 14408
rect 26049 14376 28000 14378
rect 26049 14320 26054 14376
rect 26110 14320 28000 14376
rect 26049 14318 28000 14320
rect 26049 14315 26115 14318
rect 27520 14288 28000 14318
rect 2037 14242 2103 14245
rect 4429 14242 4495 14245
rect 2037 14240 4495 14242
rect 2037 14184 2042 14240
rect 2098 14184 4434 14240
rect 4490 14184 4495 14240
rect 2037 14182 4495 14184
rect 2037 14179 2103 14182
rect 4429 14179 4495 14182
rect 7281 14242 7347 14245
rect 11237 14242 11303 14245
rect 7281 14240 11303 14242
rect 7281 14184 7286 14240
rect 7342 14184 11242 14240
rect 11298 14184 11303 14240
rect 7281 14182 11303 14184
rect 7281 14179 7347 14182
rect 11237 14179 11303 14182
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 2405 14106 2471 14109
rect 2773 14106 2839 14109
rect 2405 14104 2839 14106
rect 2405 14048 2410 14104
rect 2466 14048 2778 14104
rect 2834 14048 2839 14104
rect 2405 14046 2839 14048
rect 2405 14043 2471 14046
rect 2773 14043 2839 14046
rect 2589 13970 2655 13973
rect 2957 13970 3023 13973
rect 3141 13970 3207 13973
rect 2589 13968 3207 13970
rect 2589 13912 2594 13968
rect 2650 13912 2962 13968
rect 3018 13912 3146 13968
rect 3202 13912 3207 13968
rect 2589 13910 3207 13912
rect 2589 13907 2655 13910
rect 2957 13907 3023 13910
rect 3141 13907 3207 13910
rect 12893 13834 12959 13837
rect 14457 13834 14523 13837
rect 12893 13832 14523 13834
rect 12893 13776 12898 13832
rect 12954 13776 14462 13832
rect 14518 13776 14523 13832
rect 12893 13774 14523 13776
rect 12893 13771 12959 13774
rect 14457 13771 14523 13774
rect 24894 13772 24900 13836
rect 24964 13834 24970 13836
rect 25037 13834 25103 13837
rect 24964 13832 25103 13834
rect 24964 13776 25042 13832
rect 25098 13776 25103 13832
rect 24964 13774 25103 13776
rect 24964 13772 24970 13774
rect 25037 13771 25103 13774
rect 0 13698 480 13728
rect 4797 13698 4863 13701
rect 8385 13698 8451 13701
rect 0 13638 4538 13698
rect 0 13608 480 13638
rect 4478 13426 4538 13638
rect 4797 13696 8451 13698
rect 4797 13640 4802 13696
rect 4858 13640 8390 13696
rect 8446 13640 8451 13696
rect 4797 13638 8451 13640
rect 4797 13635 4863 13638
rect 8385 13635 8451 13638
rect 14089 13698 14155 13701
rect 17677 13698 17743 13701
rect 14089 13696 17743 13698
rect 14089 13640 14094 13696
rect 14150 13640 17682 13696
rect 17738 13640 17743 13696
rect 14089 13638 17743 13640
rect 14089 13635 14155 13638
rect 17677 13635 17743 13638
rect 22001 13698 22067 13701
rect 23381 13698 23447 13701
rect 22001 13696 23447 13698
rect 22001 13640 22006 13696
rect 22062 13640 23386 13696
rect 23442 13640 23447 13696
rect 22001 13638 23447 13640
rect 22001 13635 22067 13638
rect 23381 13635 23447 13638
rect 24710 13636 24716 13700
rect 24780 13698 24786 13700
rect 27520 13698 28000 13728
rect 24780 13638 28000 13698
rect 24780 13636 24786 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 27520 13608 28000 13638
rect 19610 13567 19930 13568
rect 6269 13562 6335 13565
rect 8477 13562 8543 13565
rect 6269 13560 8543 13562
rect 6269 13504 6274 13560
rect 6330 13504 8482 13560
rect 8538 13504 8543 13560
rect 6269 13502 8543 13504
rect 6269 13499 6335 13502
rect 8477 13499 8543 13502
rect 11605 13426 11671 13429
rect 4478 13424 11671 13426
rect 4478 13368 11610 13424
rect 11666 13368 11671 13424
rect 4478 13366 11671 13368
rect 11605 13363 11671 13366
rect 14825 13426 14891 13429
rect 21909 13426 21975 13429
rect 14825 13424 21975 13426
rect 14825 13368 14830 13424
rect 14886 13368 21914 13424
rect 21970 13368 21975 13424
rect 14825 13366 21975 13368
rect 14825 13363 14891 13366
rect 21909 13363 21975 13366
rect 10777 13290 10843 13293
rect 10910 13290 10916 13292
rect 10777 13288 10916 13290
rect 10777 13232 10782 13288
rect 10838 13232 10916 13288
rect 10777 13230 10916 13232
rect 10777 13227 10843 13230
rect 10910 13228 10916 13230
rect 10980 13228 10986 13292
rect 0 13154 480 13184
rect 9581 13154 9647 13157
rect 10685 13154 10751 13157
rect 11605 13154 11671 13157
rect 0 13094 2698 13154
rect 0 13064 480 13094
rect 2638 13018 2698 13094
rect 9581 13152 11671 13154
rect 9581 13096 9586 13152
rect 9642 13096 10690 13152
rect 10746 13096 11610 13152
rect 11666 13096 11671 13152
rect 9581 13094 11671 13096
rect 9581 13091 9647 13094
rect 10685 13091 10751 13094
rect 11605 13091 11671 13094
rect 23657 13154 23723 13157
rect 23790 13154 23796 13156
rect 23657 13152 23796 13154
rect 23657 13096 23662 13152
rect 23718 13096 23796 13152
rect 23657 13094 23796 13096
rect 23657 13091 23723 13094
rect 23790 13092 23796 13094
rect 23860 13092 23866 13156
rect 24761 13154 24827 13157
rect 27520 13154 28000 13184
rect 24761 13152 28000 13154
rect 24761 13096 24766 13152
rect 24822 13096 28000 13152
rect 24761 13094 28000 13096
rect 24761 13091 24827 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 7557 13018 7623 13021
rect 14089 13018 14155 13021
rect 2638 12958 3986 13018
rect 3926 12746 3986 12958
rect 7557 13016 14155 13018
rect 7557 12960 7562 13016
rect 7618 12960 14094 13016
rect 14150 12960 14155 13016
rect 7557 12958 14155 12960
rect 7557 12955 7623 12958
rect 14089 12955 14155 12958
rect 8661 12882 8727 12885
rect 11145 12882 11211 12885
rect 8661 12880 11211 12882
rect 8661 12824 8666 12880
rect 8722 12824 11150 12880
rect 11206 12824 11211 12880
rect 8661 12822 11211 12824
rect 8661 12819 8727 12822
rect 11145 12819 11211 12822
rect 11789 12882 11855 12885
rect 12985 12882 13051 12885
rect 11789 12880 13051 12882
rect 11789 12824 11794 12880
rect 11850 12824 12990 12880
rect 13046 12824 13051 12880
rect 11789 12822 13051 12824
rect 11789 12819 11855 12822
rect 12985 12819 13051 12822
rect 19149 12746 19215 12749
rect 3926 12686 17786 12746
rect 8385 12610 8451 12613
rect 8518 12610 8524 12612
rect 8385 12608 8524 12610
rect 8385 12552 8390 12608
rect 8446 12552 8524 12608
rect 8385 12550 8524 12552
rect 8385 12547 8451 12550
rect 8518 12548 8524 12550
rect 8588 12548 8594 12612
rect 10277 12544 10597 12545
rect 0 12474 480 12504
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 7557 12474 7623 12477
rect 0 12472 7623 12474
rect 0 12416 7562 12472
rect 7618 12416 7623 12472
rect 0 12414 7623 12416
rect 0 12384 480 12414
rect 7557 12411 7623 12414
rect 11237 12474 11303 12477
rect 17309 12474 17375 12477
rect 11237 12472 17375 12474
rect 11237 12416 11242 12472
rect 11298 12416 17314 12472
rect 17370 12416 17375 12472
rect 11237 12414 17375 12416
rect 11237 12411 11303 12414
rect 17309 12411 17375 12414
rect 3049 12338 3115 12341
rect 7373 12338 7439 12341
rect 3049 12336 7439 12338
rect 3049 12280 3054 12336
rect 3110 12280 7378 12336
rect 7434 12280 7439 12336
rect 3049 12278 7439 12280
rect 3049 12275 3115 12278
rect 7373 12275 7439 12278
rect 8845 12338 8911 12341
rect 12985 12338 13051 12341
rect 8845 12336 13051 12338
rect 8845 12280 8850 12336
rect 8906 12280 12990 12336
rect 13046 12280 13051 12336
rect 8845 12278 13051 12280
rect 8845 12275 8911 12278
rect 12985 12275 13051 12278
rect 13302 12276 13308 12340
rect 13372 12338 13378 12340
rect 13445 12338 13511 12341
rect 13372 12336 13511 12338
rect 13372 12280 13450 12336
rect 13506 12280 13511 12336
rect 13372 12278 13511 12280
rect 17726 12338 17786 12686
rect 19149 12744 22018 12746
rect 19149 12688 19154 12744
rect 19210 12688 22018 12744
rect 19149 12686 22018 12688
rect 19149 12683 19215 12686
rect 19425 12612 19491 12613
rect 19374 12548 19380 12612
rect 19444 12610 19491 12612
rect 21958 12610 22018 12686
rect 19444 12608 19536 12610
rect 19486 12552 19536 12608
rect 19444 12550 19536 12552
rect 21958 12550 22202 12610
rect 19444 12548 19491 12550
rect 19425 12547 19491 12548
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 22142 12474 22202 12550
rect 23790 12548 23796 12612
rect 23860 12610 23866 12612
rect 23933 12610 23999 12613
rect 23860 12608 23999 12610
rect 23860 12552 23938 12608
rect 23994 12552 23999 12608
rect 23860 12550 23999 12552
rect 23860 12548 23866 12550
rect 23933 12547 23999 12550
rect 27520 12474 28000 12504
rect 22142 12414 28000 12474
rect 27520 12384 28000 12414
rect 22553 12338 22619 12341
rect 17726 12336 22619 12338
rect 17726 12280 22558 12336
rect 22614 12280 22619 12336
rect 17726 12278 22619 12280
rect 13372 12276 13378 12278
rect 13445 12275 13511 12278
rect 22553 12275 22619 12278
rect 22737 12338 22803 12341
rect 23422 12338 23428 12340
rect 22737 12336 23428 12338
rect 22737 12280 22742 12336
rect 22798 12280 23428 12336
rect 22737 12278 23428 12280
rect 22737 12275 22803 12278
rect 23422 12276 23428 12278
rect 23492 12276 23498 12340
rect 7741 12202 7807 12205
rect 13353 12202 13419 12205
rect 7741 12200 13419 12202
rect 7741 12144 7746 12200
rect 7802 12144 13358 12200
rect 13414 12144 13419 12200
rect 7741 12142 13419 12144
rect 7741 12139 7807 12142
rect 13353 12139 13419 12142
rect 21265 12202 21331 12205
rect 25221 12202 25287 12205
rect 21265 12200 25287 12202
rect 21265 12144 21270 12200
rect 21326 12144 25226 12200
rect 25282 12144 25287 12200
rect 21265 12142 25287 12144
rect 21265 12139 21331 12142
rect 25221 12139 25287 12142
rect 15561 12066 15627 12069
rect 22737 12066 22803 12069
rect 15561 12064 22803 12066
rect 15561 12008 15566 12064
rect 15622 12008 22742 12064
rect 22798 12008 22803 12064
rect 15561 12006 22803 12008
rect 15561 12003 15627 12006
rect 22737 12003 22803 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 4981 11932 5047 11933
rect 4981 11930 5028 11932
rect 0 11870 4860 11930
rect 4936 11928 5028 11930
rect 4936 11872 4986 11928
rect 4936 11870 5028 11872
rect 0 11840 480 11870
rect 4800 11794 4860 11870
rect 4981 11868 5028 11870
rect 5092 11868 5098 11932
rect 18781 11930 18847 11933
rect 22277 11930 22343 11933
rect 27520 11930 28000 11960
rect 18781 11928 22343 11930
rect 18781 11872 18786 11928
rect 18842 11872 22282 11928
rect 22338 11872 22343 11928
rect 18781 11870 22343 11872
rect 4981 11867 5047 11868
rect 18781 11867 18847 11870
rect 22277 11867 22343 11870
rect 25270 11870 28000 11930
rect 11973 11794 12039 11797
rect 4800 11792 12039 11794
rect 4800 11736 11978 11792
rect 12034 11736 12039 11792
rect 4800 11734 12039 11736
rect 11973 11731 12039 11734
rect 14549 11794 14615 11797
rect 25037 11794 25103 11797
rect 14549 11792 25103 11794
rect 14549 11736 14554 11792
rect 14610 11736 25042 11792
rect 25098 11736 25103 11792
rect 14549 11734 25103 11736
rect 14549 11731 14615 11734
rect 25037 11731 25103 11734
rect 3693 11658 3759 11661
rect 13721 11658 13787 11661
rect 3693 11656 13787 11658
rect 3693 11600 3698 11656
rect 3754 11600 13726 11656
rect 13782 11600 13787 11656
rect 3693 11598 13787 11600
rect 3693 11595 3759 11598
rect 13721 11595 13787 11598
rect 16481 11658 16547 11661
rect 23473 11658 23539 11661
rect 16481 11656 23539 11658
rect 16481 11600 16486 11656
rect 16542 11600 23478 11656
rect 23534 11600 23539 11656
rect 16481 11598 23539 11600
rect 16481 11595 16547 11598
rect 23473 11595 23539 11598
rect 24485 11658 24551 11661
rect 25270 11658 25330 11870
rect 27520 11840 28000 11870
rect 24485 11656 25330 11658
rect 24485 11600 24490 11656
rect 24546 11600 25330 11656
rect 24485 11598 25330 11600
rect 24485 11595 24551 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 22645 11386 22711 11389
rect 22645 11384 25146 11386
rect 22645 11328 22650 11384
rect 22706 11328 25146 11384
rect 22645 11326 25146 11328
rect 22645 11323 22711 11326
rect 0 11250 480 11280
rect 4061 11250 4127 11253
rect 0 11248 4127 11250
rect 0 11192 4066 11248
rect 4122 11192 4127 11248
rect 0 11190 4127 11192
rect 0 11160 480 11190
rect 4061 11187 4127 11190
rect 13905 11250 13971 11253
rect 17309 11250 17375 11253
rect 13905 11248 17375 11250
rect 13905 11192 13910 11248
rect 13966 11192 17314 11248
rect 17370 11192 17375 11248
rect 13905 11190 17375 11192
rect 13905 11187 13971 11190
rect 17309 11187 17375 11190
rect 23606 11188 23612 11252
rect 23676 11250 23682 11252
rect 24577 11250 24643 11253
rect 23676 11248 24643 11250
rect 23676 11192 24582 11248
rect 24638 11192 24643 11248
rect 23676 11190 24643 11192
rect 25086 11250 25146 11326
rect 27520 11250 28000 11280
rect 25086 11190 28000 11250
rect 23676 11188 23682 11190
rect 24577 11187 24643 11190
rect 27520 11160 28000 11190
rect 3417 11114 3483 11117
rect 4429 11114 4495 11117
rect 3417 11112 4495 11114
rect 3417 11056 3422 11112
rect 3478 11056 4434 11112
rect 4490 11056 4495 11112
rect 3417 11054 4495 11056
rect 3417 11051 3483 11054
rect 4429 11051 4495 11054
rect 17585 11114 17651 11117
rect 23197 11114 23263 11117
rect 17585 11112 23263 11114
rect 17585 11056 17590 11112
rect 17646 11056 23202 11112
rect 23258 11056 23263 11112
rect 17585 11054 23263 11056
rect 17585 11051 17651 11054
rect 23197 11051 23263 11054
rect 23013 10978 23079 10981
rect 15334 10976 23079 10978
rect 15334 10920 23018 10976
rect 23074 10920 23079 10976
rect 15334 10918 23079 10920
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 5993 10842 6059 10845
rect 5993 10840 14520 10842
rect 5993 10784 5998 10840
rect 6054 10784 14520 10840
rect 5993 10782 14520 10784
rect 5993 10779 6059 10782
rect 0 10706 480 10736
rect 565 10706 631 10709
rect 0 10704 631 10706
rect 0 10648 570 10704
rect 626 10648 631 10704
rect 0 10646 631 10648
rect 14460 10706 14520 10782
rect 15334 10706 15394 10918
rect 23013 10915 23079 10918
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 16389 10842 16455 10845
rect 20989 10842 21055 10845
rect 23749 10842 23815 10845
rect 16389 10840 23815 10842
rect 16389 10784 16394 10840
rect 16450 10784 20994 10840
rect 21050 10784 23754 10840
rect 23810 10784 23815 10840
rect 16389 10782 23815 10784
rect 16389 10779 16455 10782
rect 20989 10779 21055 10782
rect 23749 10779 23815 10782
rect 14460 10646 15394 10706
rect 21633 10706 21699 10709
rect 27520 10706 28000 10736
rect 21633 10704 28000 10706
rect 21633 10648 21638 10704
rect 21694 10648 28000 10704
rect 21633 10646 28000 10648
rect 0 10616 480 10646
rect 565 10643 631 10646
rect 21633 10643 21699 10646
rect 27520 10616 28000 10646
rect 4061 10570 4127 10573
rect 12341 10570 12407 10573
rect 21173 10570 21239 10573
rect 4061 10568 21239 10570
rect 4061 10512 4066 10568
rect 4122 10512 12346 10568
rect 12402 10512 21178 10568
rect 21234 10512 21239 10568
rect 4061 10510 21239 10512
rect 4061 10507 4127 10510
rect 12341 10507 12407 10510
rect 21173 10507 21239 10510
rect 13169 10434 13235 10437
rect 13486 10434 13492 10436
rect 13169 10432 13492 10434
rect 13169 10376 13174 10432
rect 13230 10376 13492 10432
rect 13169 10374 13492 10376
rect 13169 10371 13235 10374
rect 13486 10372 13492 10374
rect 13556 10372 13562 10436
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 10777 10298 10843 10301
rect 13077 10298 13143 10301
rect 10777 10296 13143 10298
rect 10777 10240 10782 10296
rect 10838 10240 13082 10296
rect 13138 10240 13143 10296
rect 10777 10238 13143 10240
rect 10777 10235 10843 10238
rect 13077 10235 13143 10238
rect 23790 10236 23796 10300
rect 23860 10298 23866 10300
rect 23860 10238 24778 10298
rect 23860 10236 23866 10238
rect 8937 10162 9003 10165
rect 614 10160 9003 10162
rect 614 10104 8942 10160
rect 8998 10104 9003 10160
rect 614 10102 9003 10104
rect 0 10026 480 10056
rect 614 10026 674 10102
rect 8937 10099 9003 10102
rect 11513 10162 11579 10165
rect 24393 10162 24459 10165
rect 11513 10160 24459 10162
rect 11513 10104 11518 10160
rect 11574 10104 24398 10160
rect 24454 10104 24459 10160
rect 11513 10102 24459 10104
rect 11513 10099 11579 10102
rect 24393 10099 24459 10102
rect 0 9966 674 10026
rect 3877 10026 3943 10029
rect 12341 10026 12407 10029
rect 24718 10026 24778 10238
rect 27520 10026 28000 10056
rect 3877 10024 6194 10026
rect 3877 9968 3882 10024
rect 3938 9968 6194 10024
rect 3877 9966 6194 9968
rect 0 9936 480 9966
rect 3877 9963 3943 9966
rect 6134 9890 6194 9966
rect 12341 10024 17234 10026
rect 12341 9968 12346 10024
rect 12402 9968 17234 10024
rect 12341 9966 17234 9968
rect 24718 9966 28000 10026
rect 12341 9963 12407 9966
rect 13261 9890 13327 9893
rect 6134 9888 13327 9890
rect 6134 9832 13266 9888
rect 13322 9832 13327 9888
rect 6134 9830 13327 9832
rect 17174 9890 17234 9966
rect 27520 9936 28000 9966
rect 23841 9890 23907 9893
rect 17174 9888 23907 9890
rect 17174 9832 23846 9888
rect 23902 9832 23907 9888
rect 17174 9830 23907 9832
rect 13261 9827 13327 9830
rect 23841 9827 23907 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 13854 9692 13860 9756
rect 13924 9754 13930 9756
rect 24117 9754 24183 9757
rect 13924 9694 14842 9754
rect 13924 9692 13930 9694
rect 13537 9618 13603 9621
rect 614 9616 13603 9618
rect 614 9560 13542 9616
rect 13598 9560 13603 9616
rect 614 9558 13603 9560
rect 14782 9618 14842 9694
rect 15334 9752 24183 9754
rect 15334 9696 24122 9752
rect 24178 9696 24183 9752
rect 15334 9694 24183 9696
rect 15334 9618 15394 9694
rect 24117 9691 24183 9694
rect 14782 9558 15394 9618
rect 17125 9618 17191 9621
rect 24393 9618 24459 9621
rect 17125 9616 24459 9618
rect 17125 9560 17130 9616
rect 17186 9560 24398 9616
rect 24454 9560 24459 9616
rect 17125 9558 24459 9560
rect 0 9482 480 9512
rect 614 9482 674 9558
rect 13537 9555 13603 9558
rect 17125 9555 17191 9558
rect 24393 9555 24459 9558
rect 0 9422 674 9482
rect 4061 9482 4127 9485
rect 13445 9482 13511 9485
rect 4061 9480 13511 9482
rect 4061 9424 4066 9480
rect 4122 9424 13450 9480
rect 13506 9424 13511 9480
rect 4061 9422 13511 9424
rect 0 9392 480 9422
rect 4061 9419 4127 9422
rect 13445 9419 13511 9422
rect 22369 9482 22435 9485
rect 27520 9482 28000 9512
rect 22369 9480 28000 9482
rect 22369 9424 22374 9480
rect 22430 9424 28000 9480
rect 22369 9422 28000 9424
rect 22369 9419 22435 9422
rect 27520 9392 28000 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 24761 9210 24827 9213
rect 26325 9210 26391 9213
rect 24761 9208 26391 9210
rect 24761 9152 24766 9208
rect 24822 9152 26330 9208
rect 26386 9152 26391 9208
rect 24761 9150 26391 9152
rect 24761 9147 24827 9150
rect 26325 9147 26391 9150
rect 24117 9074 24183 9077
rect 25865 9074 25931 9077
rect 24117 9072 25931 9074
rect 24117 9016 24122 9072
rect 24178 9016 25870 9072
rect 25926 9016 25931 9072
rect 24117 9014 25931 9016
rect 24117 9011 24183 9014
rect 25865 9011 25931 9014
rect 15745 8938 15811 8941
rect 24761 8938 24827 8941
rect 15745 8936 24827 8938
rect 15745 8880 15750 8936
rect 15806 8880 24766 8936
rect 24822 8880 24827 8936
rect 15745 8878 24827 8880
rect 15745 8875 15811 8878
rect 24761 8875 24827 8878
rect 0 8802 480 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 480 8742
rect 4061 8739 4127 8742
rect 24669 8802 24735 8805
rect 27520 8802 28000 8832
rect 24669 8800 28000 8802
rect 24669 8744 24674 8800
rect 24730 8744 28000 8800
rect 24669 8742 28000 8744
rect 24669 8739 24735 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 27520 8712 28000 8742
rect 24277 8671 24597 8672
rect 12525 8394 12591 8397
rect 20437 8394 20503 8397
rect 12525 8392 20503 8394
rect 12525 8336 12530 8392
rect 12586 8336 20442 8392
rect 20498 8336 20503 8392
rect 12525 8334 20503 8336
rect 12525 8331 12591 8334
rect 20437 8331 20503 8334
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 20069 8258 20135 8261
rect 27520 8258 28000 8288
rect 20069 8256 28000 8258
rect 20069 8200 20074 8256
rect 20130 8200 28000 8256
rect 20069 8198 28000 8200
rect 20069 8195 20135 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 27520 8168 28000 8198
rect 19610 8127 19930 8128
rect 16389 7986 16455 7989
rect 2776 7984 16455 7986
rect 2776 7928 16394 7984
rect 16450 7928 16455 7984
rect 2776 7926 16455 7928
rect 2776 7714 2836 7926
rect 16389 7923 16455 7926
rect 4061 7850 4127 7853
rect 23933 7850 23999 7853
rect 4061 7848 23999 7850
rect 4061 7792 4066 7848
rect 4122 7792 23938 7848
rect 23994 7792 23999 7848
rect 4061 7790 23999 7792
rect 4061 7787 4127 7790
rect 23933 7787 23999 7790
rect 2638 7654 2836 7714
rect 0 7578 480 7608
rect 2638 7578 2698 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 27520 7578 28000 7608
rect 0 7518 2698 7578
rect 24902 7518 28000 7578
rect 0 7488 480 7518
rect 16849 7442 16915 7445
rect 3006 7440 16915 7442
rect 3006 7384 16854 7440
rect 16910 7384 16915 7440
rect 3006 7382 16915 7384
rect 565 7306 631 7309
rect 3006 7306 3066 7382
rect 16849 7379 16915 7382
rect 22001 7442 22067 7445
rect 24902 7442 24962 7518
rect 27520 7488 28000 7518
rect 22001 7440 24962 7442
rect 22001 7384 22006 7440
rect 22062 7384 24962 7440
rect 22001 7382 24962 7384
rect 22001 7379 22067 7382
rect 565 7304 3066 7306
rect 565 7248 570 7304
rect 626 7248 3066 7304
rect 565 7246 3066 7248
rect 565 7243 631 7246
rect 10277 7104 10597 7105
rect 0 7034 480 7064
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 565 7034 631 7037
rect 0 7032 631 7034
rect 0 6976 570 7032
rect 626 6976 631 7032
rect 0 6974 631 6976
rect 0 6944 480 6974
rect 565 6971 631 6974
rect 20161 7034 20227 7037
rect 27520 7034 28000 7064
rect 20161 7032 28000 7034
rect 20161 6976 20166 7032
rect 20222 6976 28000 7032
rect 20161 6974 28000 6976
rect 20161 6971 20227 6974
rect 27520 6944 28000 6974
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 3877 6354 3943 6357
rect 0 6352 3943 6354
rect 0 6296 3882 6352
rect 3938 6296 3943 6352
rect 0 6294 3943 6296
rect 0 6264 480 6294
rect 3877 6291 3943 6294
rect 17493 6354 17559 6357
rect 27520 6354 28000 6384
rect 17493 6352 28000 6354
rect 17493 6296 17498 6352
rect 17554 6296 28000 6352
rect 17493 6294 28000 6296
rect 17493 6291 17559 6294
rect 27520 6264 28000 6294
rect 24669 6082 24735 6085
rect 24669 6080 26618 6082
rect 24669 6024 24674 6080
rect 24730 6024 26618 6080
rect 24669 6022 26618 6024
rect 24669 6019 24735 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 24669 5946 24735 5949
rect 26417 5946 26483 5949
rect 24669 5944 26483 5946
rect 24669 5888 24674 5944
rect 24730 5888 26422 5944
rect 26478 5888 26483 5944
rect 24669 5886 26483 5888
rect 24669 5883 24735 5886
rect 26417 5883 26483 5886
rect 0 5810 480 5840
rect 24485 5810 24551 5813
rect 0 5808 24551 5810
rect 0 5752 24490 5808
rect 24546 5752 24551 5808
rect 0 5750 24551 5752
rect 26558 5810 26618 6022
rect 27520 5810 28000 5840
rect 26558 5750 28000 5810
rect 0 5720 480 5750
rect 24485 5747 24551 5750
rect 27520 5720 28000 5750
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 0 5130 480 5160
rect 3693 5130 3759 5133
rect 0 5128 3759 5130
rect 0 5072 3698 5128
rect 3754 5072 3759 5128
rect 0 5070 3759 5072
rect 0 5040 480 5070
rect 3693 5067 3759 5070
rect 23473 5130 23539 5133
rect 27520 5130 28000 5160
rect 23473 5128 28000 5130
rect 23473 5072 23478 5128
rect 23534 5072 28000 5128
rect 23473 5070 28000 5072
rect 23473 5067 23539 5070
rect 27520 5040 28000 5070
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 24117 4722 24183 4725
rect 24485 4722 24551 4725
rect 2776 4720 24551 4722
rect 2776 4664 24122 4720
rect 24178 4664 24490 4720
rect 24546 4664 24551 4720
rect 2776 4662 24551 4664
rect 0 4586 480 4616
rect 0 4526 2698 4586
rect 0 4496 480 4526
rect 2638 4450 2698 4526
rect 2776 4450 2836 4662
rect 24117 4659 24183 4662
rect 24485 4659 24551 4662
rect 24761 4586 24827 4589
rect 27520 4586 28000 4616
rect 24761 4584 28000 4586
rect 24761 4528 24766 4584
rect 24822 4528 28000 4584
rect 24761 4526 28000 4528
rect 24761 4523 24827 4526
rect 27520 4496 28000 4526
rect 2638 4390 2836 4450
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 17033 4042 17099 4045
rect 4846 4040 17099 4042
rect 4846 3984 17038 4040
rect 17094 3984 17099 4040
rect 4846 3982 17099 3984
rect 0 3906 480 3936
rect 4846 3906 4906 3982
rect 17033 3979 17099 3982
rect 0 3846 4906 3906
rect 24577 3906 24643 3909
rect 27520 3906 28000 3936
rect 24577 3904 28000 3906
rect 24577 3848 24582 3904
rect 24638 3848 28000 3904
rect 24577 3846 28000 3848
rect 0 3816 480 3846
rect 24577 3843 24643 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 27520 3816 28000 3846
rect 19610 3775 19930 3776
rect 9489 3634 9555 3637
rect 13905 3634 13971 3637
rect 9489 3632 13971 3634
rect 9489 3576 9494 3632
rect 9550 3576 13910 3632
rect 13966 3576 13971 3632
rect 9489 3574 13971 3576
rect 9489 3571 9555 3574
rect 13905 3571 13971 3574
rect 17309 3634 17375 3637
rect 17309 3632 24962 3634
rect 17309 3576 17314 3632
rect 17370 3576 24962 3632
rect 17309 3574 24962 3576
rect 17309 3571 17375 3574
rect 2773 3498 2839 3501
rect 12157 3498 12223 3501
rect 2773 3496 12223 3498
rect 2773 3440 2778 3496
rect 2834 3440 12162 3496
rect 12218 3440 12223 3496
rect 2773 3438 12223 3440
rect 2773 3435 2839 3438
rect 12157 3435 12223 3438
rect 12893 3498 12959 3501
rect 23473 3498 23539 3501
rect 12893 3496 23539 3498
rect 12893 3440 12898 3496
rect 12954 3440 23478 3496
rect 23534 3440 23539 3496
rect 12893 3438 23539 3440
rect 12893 3435 12959 3438
rect 23473 3435 23539 3438
rect 0 3362 480 3392
rect 2957 3362 3023 3365
rect 0 3360 3023 3362
rect 0 3304 2962 3360
rect 3018 3304 3023 3360
rect 0 3302 3023 3304
rect 24902 3362 24962 3574
rect 27520 3362 28000 3392
rect 24902 3302 28000 3362
rect 0 3272 480 3302
rect 2957 3299 3023 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 27520 3272 28000 3302
rect 24277 3231 24597 3232
rect 8293 2954 8359 2957
rect 12433 2954 12499 2957
rect 8293 2952 12499 2954
rect 8293 2896 8298 2952
rect 8354 2896 12438 2952
rect 12494 2896 12499 2952
rect 8293 2894 12499 2896
rect 8293 2891 8359 2894
rect 12433 2891 12499 2894
rect 10277 2752 10597 2753
rect 0 2682 480 2712
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 3509 2682 3575 2685
rect 0 2680 3575 2682
rect 0 2624 3514 2680
rect 3570 2624 3575 2680
rect 0 2622 3575 2624
rect 0 2592 480 2622
rect 3509 2619 3575 2622
rect 23749 2682 23815 2685
rect 27520 2682 28000 2712
rect 23749 2680 28000 2682
rect 23749 2624 23754 2680
rect 23810 2624 28000 2680
rect 23749 2622 28000 2624
rect 23749 2619 23815 2622
rect 27520 2592 28000 2622
rect 1301 2410 1367 2413
rect 18505 2410 18571 2413
rect 1301 2408 18571 2410
rect 1301 2352 1306 2408
rect 1362 2352 18510 2408
rect 18566 2352 18571 2408
rect 1301 2350 18571 2352
rect 1301 2347 1367 2350
rect 18505 2347 18571 2350
rect 23841 2410 23907 2413
rect 23841 2408 25514 2410
rect 23841 2352 23846 2408
rect 23902 2352 25514 2408
rect 23841 2350 25514 2352
rect 23841 2347 23907 2350
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 5165 2138 5231 2141
rect 0 2136 5231 2138
rect 0 2080 5170 2136
rect 5226 2080 5231 2136
rect 0 2078 5231 2080
rect 25454 2138 25514 2350
rect 27520 2138 28000 2168
rect 25454 2078 28000 2138
rect 0 2048 480 2078
rect 5165 2075 5231 2078
rect 27520 2048 28000 2078
rect 0 1458 480 1488
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1368 480 1398
rect 2865 1395 2931 1398
rect 20437 1458 20503 1461
rect 27520 1458 28000 1488
rect 20437 1456 28000 1458
rect 20437 1400 20442 1456
rect 20498 1400 28000 1456
rect 20437 1398 28000 1400
rect 20437 1395 20503 1398
rect 27520 1368 28000 1398
rect 0 914 480 944
rect 4061 914 4127 917
rect 0 912 4127 914
rect 0 856 4066 912
rect 4122 856 4127 912
rect 0 854 4127 856
rect 0 824 480 854
rect 4061 851 4127 854
rect 23473 914 23539 917
rect 27520 914 28000 944
rect 23473 912 28000 914
rect 23473 856 23478 912
rect 23534 856 28000 912
rect 23473 854 28000 856
rect 23473 851 23539 854
rect 27520 824 28000 854
rect 0 370 480 400
rect 3417 370 3483 373
rect 27520 370 28000 400
rect 0 368 3483 370
rect 0 312 3422 368
rect 3478 312 3483 368
rect 0 310 3483 312
rect 0 280 480 310
rect 3417 307 3483 310
rect 27478 280 28000 370
rect 14457 98 14523 101
rect 27478 98 27538 280
rect 14457 96 27538 98
rect 14457 40 14462 96
rect 14518 40 27538 96
rect 14457 38 27538 40
rect 14457 35 14523 38
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 11284 24516 11348 24580
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 13860 24380 13924 24444
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 14228 22128 14292 22132
rect 14228 22072 14278 22128
rect 14278 22072 14292 22128
rect 14228 22068 14292 22072
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 17908 21388 17972 21452
rect 12388 21252 12452 21316
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 23796 20980 23860 21044
rect 2636 20708 2700 20772
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 12388 20436 12452 20500
rect 14228 20224 14292 20228
rect 14228 20168 14278 20224
rect 14278 20168 14292 20224
rect 14228 20164 14292 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 24900 18668 24964 18732
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 13492 18396 13556 18460
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 24716 17580 24780 17644
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 23612 16356 23676 16420
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 13308 15676 13372 15740
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 23428 14724 23492 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 12940 14588 13004 14652
rect 3924 14316 3988 14380
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 24900 13772 24964 13836
rect 24716 13636 24780 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 10916 13228 10980 13292
rect 23796 13092 23860 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 8524 12548 8588 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 13308 12276 13372 12340
rect 19380 12608 19444 12612
rect 19380 12552 19430 12608
rect 19430 12552 19444 12608
rect 19380 12548 19444 12552
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 23796 12548 23860 12612
rect 23428 12276 23492 12340
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 5028 11928 5092 11932
rect 5028 11872 5042 11928
rect 5042 11872 5092 11928
rect 5028 11868 5092 11872
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 23612 11188 23676 11252
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 13492 10372 13556 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 23796 10236 23860 10300
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 13860 9692 13924 9756
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 2638 20773 2698 21302
rect 2635 20772 2701 20773
rect 2635 20708 2636 20772
rect 2700 20708 2701 20772
rect 2635 20707 2701 20708
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 3923 14380 3989 14381
rect 3923 14316 3924 14380
rect 3988 14316 3989 14380
rect 3923 14315 3989 14316
rect 3926 14058 3986 14315
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 11283 24580 11349 24581
rect 11283 24516 11284 24580
rect 11348 24516 11349 24580
rect 11283 24515 11349 24516
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 11286 18818 11346 24515
rect 13859 24444 13925 24445
rect 13859 24380 13860 24444
rect 13924 24380 13925 24444
rect 13859 24379 13925 24380
rect 12387 21316 12453 21317
rect 12387 21252 12388 21316
rect 12452 21252 12453 21316
rect 12387 21251 12453 21252
rect 12390 20501 12450 21251
rect 12387 20500 12453 20501
rect 12387 20436 12388 20500
rect 12452 20436 12453 20500
rect 12387 20435 12453 20436
rect 13491 18460 13557 18461
rect 13491 18396 13492 18460
rect 13556 18396 13557 18460
rect 13491 18395 13557 18396
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 13307 15740 13373 15741
rect 13307 15676 13308 15740
rect 13372 15676 13373 15740
rect 13307 15675 13373 15676
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 12939 14652 13005 14653
rect 12939 14588 12940 14652
rect 13004 14588 13005 14652
rect 12939 14587 13005 14588
rect 12942 14058 13002 14587
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 11456 10597 12480
rect 13310 12341 13370 15675
rect 13307 12340 13373 12341
rect 13307 12276 13308 12340
rect 13372 12276 13373 12340
rect 13307 12275 13373 12276
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 13494 10437 13554 18395
rect 13862 12018 13922 24379
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14227 22132 14293 22133
rect 14227 22068 14228 22132
rect 14292 22068 14293 22132
rect 14227 22067 14293 22068
rect 14230 20229 14290 22067
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14227 20228 14293 20229
rect 14227 20164 14228 20228
rect 14292 20164 14293 20228
rect 14227 20163 14293 20164
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 23795 21044 23861 21045
rect 23795 20980 23796 21044
rect 23860 20980 23861 21044
rect 23795 20979 23861 20980
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 23611 16420 23677 16421
rect 23611 16356 23612 16420
rect 23676 16356 23677 16420
rect 23611 16355 23677 16356
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 23427 14788 23493 14789
rect 23427 14724 23428 14788
rect 23492 14724 23493 14788
rect 23427 14723 23493 14724
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 13491 10436 13557 10437
rect 13491 10372 13492 10436
rect 13556 10372 13557 10436
rect 13491 10371 13557 10372
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 13862 9757 13922 11782
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 13859 9756 13925 9757
rect 13859 9692 13860 9756
rect 13924 9692 13925 9756
rect 13859 9691 13925 9692
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 11456 19930 12480
rect 23430 12341 23490 14723
rect 23427 12340 23493 12341
rect 23427 12276 23428 12340
rect 23492 12276 23493 12340
rect 23427 12275 23493 12276
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 23614 11253 23674 16355
rect 23798 13157 23858 20979
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24715 17644 24781 17645
rect 24715 17580 24716 17644
rect 24780 17580 24781 17644
rect 24715 17579 24781 17580
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 23795 13156 23861 13157
rect 23795 13092 23796 13156
rect 23860 13092 23861 13156
rect 23795 13091 23861 13092
rect 24277 13088 24597 14112
rect 24718 13701 24778 17579
rect 24899 13836 24965 13837
rect 24899 13772 24900 13836
rect 24964 13772 24965 13836
rect 24899 13771 24965 13772
rect 24715 13700 24781 13701
rect 24715 13636 24716 13700
rect 24780 13636 24781 13700
rect 24715 13635 24781 13636
rect 24902 13378 24962 13771
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23795 12612 23861 12613
rect 23795 12548 23796 12612
rect 23860 12548 23861 12612
rect 23795 12547 23861 12548
rect 23611 11252 23677 11253
rect 23611 11188 23612 11252
rect 23676 11188 23677 11252
rect 23611 11187 23677 11188
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 23798 10301 23858 12547
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 23795 10300 23861 10301
rect 23795 10236 23796 10300
rect 23860 10236 23861 10300
rect 23795 10235 23861 10236
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 2550 21302 2786 21538
rect 3838 13822 4074 14058
rect 4942 11932 5178 12018
rect 4942 11868 5028 11932
rect 5028 11868 5092 11932
rect 5092 11868 5178 11932
rect 4942 11782 5178 11868
rect 11198 18582 11434 18818
rect 12854 13822 13090 14058
rect 8438 12612 8674 12698
rect 8438 12548 8524 12612
rect 8524 12548 8588 12612
rect 8588 12548 8674 12612
rect 8438 12462 8674 12548
rect 10830 13292 11066 13378
rect 10830 13228 10916 13292
rect 10916 13228 10980 13292
rect 10980 13228 11066 13292
rect 10830 13142 11066 13228
rect 17822 21452 18058 21538
rect 17822 21388 17908 21452
rect 17908 21388 17972 21452
rect 17972 21388 18058 21452
rect 17822 21302 18058 21388
rect 13774 11782 14010 12018
rect 19294 12612 19530 12698
rect 19294 12548 19380 12612
rect 19380 12548 19444 12612
rect 19444 12548 19530 12612
rect 19294 12462 19530 12548
rect 24814 18732 25050 18818
rect 24814 18668 24900 18732
rect 24900 18668 24964 18732
rect 24964 18668 25050 18732
rect 24814 18582 25050 18668
rect 24814 13142 25050 13378
<< metal5 >>
rect 2508 21538 18100 21580
rect 2508 21302 2550 21538
rect 2786 21302 17822 21538
rect 18058 21302 18100 21538
rect 2508 21260 18100 21302
rect 11156 18818 25092 18860
rect 11156 18582 11198 18818
rect 11434 18582 24814 18818
rect 25050 18582 25092 18818
rect 11156 18540 25092 18582
rect 3796 14058 13132 14100
rect 3796 13822 3838 14058
rect 4074 13822 12854 14058
rect 13090 13822 13132 14058
rect 3796 13780 13132 13822
rect 10788 13378 25092 13420
rect 10788 13142 10830 13378
rect 11066 13142 24814 13378
rect 25050 13142 25092 13378
rect 10788 13100 25092 13142
rect 8396 12698 19572 12740
rect 8396 12462 8438 12698
rect 8674 12462 19294 12698
rect 19530 12462 19572 12698
rect 8396 12420 19572 12462
rect 4900 12018 14052 12060
rect 4900 11782 4942 12018
rect 5178 11782 13774 12018
rect 14010 11782 14052 12018
rect 4900 11740 14052 11782
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1604681595
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _056_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604681595
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 1604681595
transform 1 0 18676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_195
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_207
timestamp 1604681595
transform 1 0 20148 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604681595
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604681595
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604681595
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1604681595
transform 1 0 24380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1604681595
transform 1 0 25484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_269
timestamp 1604681595
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604681595
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604681595
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604681595
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604681595
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604681595
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_252
timestamp 1604681595
transform 1 0 24288 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_256
timestamp 1604681595
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_260
timestamp 1604681595
transform 1 0 25024 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_272
timestamp 1604681595
transform 1 0 26128 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_276
timestamp 1604681595
transform 1 0 26496 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 24104 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_239
timestamp 1604681595
transform 1 0 23092 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_247
timestamp 1604681595
transform 1 0 23828 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_259
timestamp 1604681595
transform 1 0 24932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_271
timestamp 1604681595
transform 1 0 26036 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604681595
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_253
timestamp 1604681595
transform 1 0 24380 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_256
timestamp 1604681595
transform 1 0 24656 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_268
timestamp 1604681595
transform 1 0 25760 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_276
timestamp 1604681595
transform 1 0 26496 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1604681595
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604681595
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604681595
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604681595
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604681595
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604681595
transform 1 0 24472 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1604681595
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1604681595
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_269
timestamp 1604681595
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604681595
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1604681595
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604681595
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604681595
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1604681595
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1604681595
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1604681595
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1604681595
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1604681595
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1604681595
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1604681595
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_269
timestamp 1604681595
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1604681595
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1604681595
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1604681595
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1604681595
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1604681595
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1604681595
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1604681595
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604681595
transform 1 0 23920 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604681595
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1604681595
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_256
timestamp 1604681595
transform 1 0 24656 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_260
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_272
timestamp 1604681595
transform 1 0 26128 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_276
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1604681595
transform 1 0 14076 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_144
timestamp 1604681595
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1604681595
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1604681595
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604681595
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604681595
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_251
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_259
timestamp 1604681595
transform 1 0 24932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1604681595
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_125
timestamp 1604681595
transform 1 0 12604 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp 1604681595
transform 1 0 12880 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12696 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12696 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1604681595
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1604681595
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_136
timestamp 1604681595
transform 1 0 13616 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1604681595
transform 1 0 14720 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _029_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1604681595
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1604681595
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1604681595
transform 1 0 16284 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_172
timestamp 1604681595
transform 1 0 16928 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1604681595
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1604681595
transform 1 0 17388 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1604681595
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_189
timestamp 1604681595
transform 1 0 18492 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1604681595
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1604681595
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_235
timestamp 1604681595
transform 1 0 22724 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_231
timestamp 1604681595
transform 1 0 22356 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604681595
transform 1 0 22448 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_247
timestamp 1604681595
transform 1 0 23828 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1604681595
transform 1 0 24012 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604681595
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604681595
transform 1 0 23460 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604681595
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604681595
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604681595
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604681595
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_263
timestamp 1604681595
transform 1 0 25300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1604681595
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_20
timestamp 1604681595
transform 1 0 2944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_24
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_36
timestamp 1604681595
transform 1 0 4416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_48
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1604681595
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1604681595
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1604681595
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_147
timestamp 1604681595
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1604681595
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_164
timestamp 1604681595
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16836 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_168
timestamp 1604681595
transform 1 0 16560 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_173
timestamp 1604681595
transform 1 0 17020 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1604681595
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604681595
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_220
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604681595
transform 1 0 22540 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1604681595
transform 1 0 22816 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604681595
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604681595
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604681595
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_263
timestamp 1604681595
transform 1 0 25300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_275
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604681595
transform 1 0 1564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 1604681595
transform 1 0 2760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1604681595
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1604681595
transform 1 0 3496 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1604681595
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1604681595
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_40
timestamp 1604681595
transform 1 0 4784 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_52
timestamp 1604681595
transform 1 0 5888 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_76
timestamp 1604681595
transform 1 0 8096 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1604681595
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604681595
transform 1 0 11040 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12052 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_107
timestamp 1604681595
transform 1 0 10948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1604681595
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1604681595
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1604681595
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 16284 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604681595
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16652 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1604681595
transform 1 0 16468 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_180
timestamp 1604681595
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1604681595
transform 1 0 18032 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1604681595
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1604681595
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_218
timestamp 1604681595
transform 1 0 21160 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604681595
transform 1 0 23000 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23920 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_230
timestamp 1604681595
transform 1 0 22264 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_242
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1604681595
transform 1 0 24104 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604681595
transform 1 0 24564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24288 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_254
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_259
timestamp 1604681595
transform 1 0 24932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_271
timestamp 1604681595
transform 1 0 26036 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3864 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 3496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_24
timestamp 1604681595
transform 1 0 3312 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_28
timestamp 1604681595
transform 1 0 3680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1604681595
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_45
timestamp 1604681595
transform 1 0 5244 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1604681595
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_78
timestamp 1604681595
transform 1 0 8280 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10580 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1604681595
transform 1 0 9384 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_94
timestamp 1604681595
transform 1 0 9752 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_97
timestamp 1604681595
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_101
timestamp 1604681595
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1604681595
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_140
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_144
timestamp 1604681595
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16100 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14536 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15916 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1604681595
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_159
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1604681595
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_192
timestamp 1604681595
transform 1 0 18768 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_203
timestamp 1604681595
transform 1 0 19780 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604681595
transform 1 0 21896 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604681595
transform 1 0 21160 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_215
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_224
timestamp 1604681595
transform 1 0 21712 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_228
timestamp 1604681595
transform 1 0 22080 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604681595
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604681595
transform 1 0 25484 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_257
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_261
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_269
timestamp 1604681595
transform 1 0 25852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604681595
transform 1 0 26036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_273
timestamp 1604681595
transform 1 0 26220 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1604681595
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5520 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_50
timestamp 1604681595
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1604681595
transform 1 0 6072 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_64
timestamp 1604681595
transform 1 0 6992 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_81
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1604681595
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_99
timestamp 1604681595
transform 1 0 10212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1604681595
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10948 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13432 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1604681595
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1604681595
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1604681595
transform 1 0 17664 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_187
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18400 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1604681595
transform 1 0 19228 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1604681595
transform 1 0 19596 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1604681595
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_225
timestamp 1604681595
transform 1 0 21804 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604681595
transform 1 0 22540 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23092 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_237
timestamp 1604681595
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_241
timestamp 1604681595
transform 1 0 23276 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_264
timestamp 1604681595
transform 1 0 25392 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_272
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_7
timestamp 1604681595
transform 1 0 1748 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2024 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604681595
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_36
timestamp 1604681595
transform 1 0 4416 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604681595
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604681595
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1604681595
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9108 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_85
timestamp 1604681595
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604681595
transform 1 0 9292 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_103
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604681595
transform 1 0 9752 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10212 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_122
timestamp 1604681595
transform 1 0 12328 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1604681595
transform 1 0 11960 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_19_141
timestamp 1604681595
transform 1 0 14076 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14812 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_146
timestamp 1604681595
transform 1 0 14536 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_177
timestamp 1604681595
transform 1 0 17388 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_173
timestamp 1604681595
transform 1 0 17020 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604681595
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18124 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17940 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 19688 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 1604681595
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_202
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_206
timestamp 1604681595
transform 1 0 20056 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_215
timestamp 1604681595
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1604681595
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21068 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1604681595
transform 1 0 22080 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_228
timestamp 1604681595
transform 1 0 22080 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 21896 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21252 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_236
timestamp 1604681595
transform 1 0 22816 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_236
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_232
timestamp 1604681595
transform 1 0 22448 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604681595
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22632 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 22264 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604681595
transform 1 0 22448 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_244
timestamp 1604681595
transform 1 0 23552 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_240
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_240
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23828 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_38.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_19_266
timestamp 1604681595
transform 1 0 25576 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1604681595
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2668 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_13
timestamp 1604681595
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_36
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_79
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8832 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_107
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11132 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604681595
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_140
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_144
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1604681595
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1604681595
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_179
timestamp 1604681595
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1604681595
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1604681595
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_228
timestamp 1604681595
transform 1 0 22080 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604681595
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_254
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604681595
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_268
timestamp 1604681595
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_272
timestamp 1604681595
transform 1 0 26128 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_276
timestamp 1604681595
transform 1 0 26496 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1472 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4140 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 5704 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 8648 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1604681595
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604681595
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_101
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11132 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_108
timestamp 1604681595
transform 1 0 11040 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1604681595
transform 1 0 11960 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1604681595
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_125
timestamp 1604681595
transform 1 0 12604 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_135
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1604681595
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1604681595
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17572 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_173
timestamp 1604681595
transform 1 0 17020 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_177
timestamp 1604681595
transform 1 0 17388 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1604681595
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_204
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_208
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 22816 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_234
timestamp 1604681595
transform 1 0 22632 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 1604681595
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_251
timestamp 1604681595
transform 1 0 24196 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_255
timestamp 1604681595
transform 1 0 24564 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_265
timestamp 1604681595
transform 1 0 25484 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_273
timestamp 1604681595
transform 1 0 26220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1604681595
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1604681595
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1604681595
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_45
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604681595
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1604681595
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_82
timestamp 1604681595
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 9568 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_86
timestamp 1604681595
transform 1 0 9016 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_111
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_115
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604681595
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13984 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_136
timestamp 1604681595
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1604681595
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1604681595
transform 1 0 15180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604681595
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 19964 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1604681595
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_207
timestamp 1604681595
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1604681595
transform 1 0 20884 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1604681595
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_224
timestamp 1604681595
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_228
timestamp 1604681595
transform 1 0 22080 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604681595
transform 1 0 22448 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23736 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604681595
transform 1 0 22264 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604681595
transform 1 0 25300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_255
timestamp 1604681595
transform 1 0 24564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_259
timestamp 1604681595
transform 1 0 24932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_267
timestamp 1604681595
transform 1 0 25668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_271
timestamp 1604681595
transform 1 0 26036 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_18
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3496 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_24
timestamp 1604681595
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1604681595
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_40
timestamp 1604681595
transform 1 0 4784 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5520 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 4968 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_47
timestamp 1604681595
transform 1 0 5428 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1604681595
transform 1 0 6348 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_61
timestamp 1604681595
transform 1 0 6716 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604681595
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604681595
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1604681595
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604681595
transform 1 0 9844 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10856 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604681595
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15732 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15548 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1604681595
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604681595
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604681595
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604681595
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_195
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1604681595
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604681595
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_224
timestamp 1604681595
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 1604681595
transform 1 0 22080 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23368 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 22448 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1604681595
transform 1 0 22724 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_239
timestamp 1604681595
transform 1 0 23092 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_261
timestamp 1604681595
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_273
timestamp 1604681595
transform 1 0 26220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_9
timestamp 1604681595
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1604681595
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_31
timestamp 1604681595
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 8188 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1604681595
transform 1 0 7452 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1604681595
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_96
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 13984 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1604681595
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1604681595
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604681595
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_149
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_156
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1604681595
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604681595
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604681595
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1604681595
transform 1 0 20148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1604681595
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23736 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1604681595
transform 1 0 22816 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 24748 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_255
timestamp 1604681595
transform 1 0 24564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_259
timestamp 1604681595
transform 1 0 24932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_267
timestamp 1604681595
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_271
timestamp 1604681595
transform 1 0 26036 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_10
timestamp 1604681595
transform 1 0 2024 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 1840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_34
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_30
timestamp 1604681595
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_38
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4876 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1604681595
transform 1 0 5244 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_42
timestamp 1604681595
transform 1 0 4968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5060 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5336 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1604681595
transform 1 0 7452 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_65
timestamp 1604681595
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604681595
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_77
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8280 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1604681595
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_97
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604681595
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13340 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_135
timestamp 1604681595
transform 1 0 13524 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604681595
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_163
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_159
timestamp 1604681595
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_172
timestamp 1604681595
transform 1 0 16928 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1604681595
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604681595
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 17020 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_192
timestamp 1604681595
transform 1 0 18768 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1604681595
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_201
timestamp 1604681595
transform 1 0 19596 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604681595
transform 1 0 19504 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_206
timestamp 1604681595
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_204
timestamp 1604681595
transform 1 0 19872 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19872 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_208
timestamp 1604681595
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_229
timestamp 1604681595
transform 1 0 22172 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_237
timestamp 1604681595
transform 1 0 22908 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_233
timestamp 1604681595
transform 1 0 22540 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_238
timestamp 1604681595
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604681595
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_242
timestamp 1604681595
transform 1 0 23368 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23552 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23736 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_265
timestamp 1604681595
transform 1 0 25484 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_268
timestamp 1604681595
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 1604681595
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_272
timestamp 1604681595
transform 1 0 26128 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1604681595
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_25
timestamp 1604681595
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604681595
transform 1 0 6532 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1604681595
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1604681595
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1604681595
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1604681595
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1604681595
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_107
timestamp 1604681595
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 13524 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1604681595
transform 1 0 13340 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_137
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604681595
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 17756 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17572 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1604681595
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1604681595
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1604681595
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_204
timestamp 1604681595
transform 1 0 19872 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1604681595
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1604681595
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604681595
transform 1 0 22448 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23644 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23460 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_236
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_242
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_264
timestamp 1604681595
transform 1 0 25392 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_272
timestamp 1604681595
transform 1 0 26128 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2300 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1604681595
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_12
timestamp 1604681595
transform 1 0 2208 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_32
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604681595
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1604681595
transform 1 0 4784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_53
timestamp 1604681595
transform 1 0 5980 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_77
timestamp 1604681595
transform 1 0 8188 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1604681595
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_103
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604681595
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_107
timestamp 1604681595
transform 1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12972 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_152
timestamp 1604681595
transform 1 0 15088 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604681595
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 19964 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19780 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21528 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_214
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1604681595
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1604681595
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1604681595
transform 1 0 22724 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604681595
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1604681595
transform 1 0 25392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_268
timestamp 1604681595
transform 1 0 25760 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604681595
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 2024 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_19
timestamp 1604681595
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 3036 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604681595
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4784 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6440 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_49
timestamp 1604681595
transform 1 0 5612 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1604681595
transform 1 0 6072 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1604681595
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_120
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_125
timestamp 1604681595
transform 1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12880 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13984 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1604681595
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16284 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1604681595
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_150
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1604681595
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17572 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_167
timestamp 1604681595
transform 1 0 16468 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_175
timestamp 1604681595
transform 1 0 17204 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19320 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19136 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1604681595
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_204
timestamp 1604681595
transform 1 0 19872 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_208
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_228
timestamp 1604681595
transform 1 0 22080 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604681595
transform 1 0 22448 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23460 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22264 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604681595
transform 1 0 25024 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 24472 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_252
timestamp 1604681595
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_256
timestamp 1604681595
transform 1 0 24656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_264
timestamp 1604681595
transform 1 0 25392 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604681595
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 2392 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1604681595
transform 1 0 1932 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_13
timestamp 1604681595
transform 1 0 2300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_16
timestamp 1604681595
transform 1 0 2576 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 4232 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1604681595
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1604681595
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1604681595
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_75
timestamp 1604681595
transform 1 0 8004 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_79
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1604681595
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_95
timestamp 1604681595
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_108
timestamp 1604681595
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_112
timestamp 1604681595
transform 1 0 11408 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1604681595
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1604681595
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604681595
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_193
timestamp 1604681595
transform 1 0 18860 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1604681595
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_205
timestamp 1604681595
transform 1 0 19964 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 20792 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1604681595
transform 1 0 20424 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23736 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1604681595
transform 1 0 22540 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_255
timestamp 1604681595
transform 1 0 24564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_259
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_269
timestamp 1604681595
transform 1 0 25852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 26036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_273
timestamp 1604681595
transform 1 0 26220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604681595
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_6
timestamp 1604681595
transform 1 0 1656 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_10
timestamp 1604681595
transform 1 0 2024 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604681595
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4232 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4784 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1604681595
transform 1 0 6532 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7268 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8648 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1604681595
transform 1 0 8096 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_88
timestamp 1604681595
transform 1 0 9200 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_99
timestamp 1604681595
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604681595
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18216 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17756 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 17572 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_173
timestamp 1604681595
transform 1 0 17020 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1604681595
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604681595
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_205
timestamp 1604681595
transform 1 0 19964 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 20976 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_209
timestamp 1604681595
transform 1 0 20332 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23736 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23092 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_235
timestamp 1604681595
transform 1 0 22724 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_241
timestamp 1604681595
transform 1 0 23276 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_245
timestamp 1604681595
transform 1 0 23644 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1604681595
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604681595
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_6
timestamp 1604681595
transform 1 0 1656 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1604681595
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604681595
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_10
timestamp 1604681595
transform 1 0 2024 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_11
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1604681595
transform 1 0 2576 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_23
timestamp 1604681595
transform 1 0 3220 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_25
timestamp 1604681595
transform 1 0 3404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3404 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 1604681595
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_36
timestamp 1604681595
transform 1 0 4416 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1604681595
transform 1 0 4140 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4600 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4232 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4876 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_45
timestamp 1604681595
transform 1 0 5244 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1604681595
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604681595
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_60
timestamp 1604681595
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_64
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1604681595
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_68
timestamp 1604681595
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604681595
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_81
timestamp 1604681595
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_77
timestamp 1604681595
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8096 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_89
timestamp 1604681595
transform 1 0 9292 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1604681595
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1604681595
transform 1 0 10028 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_95
timestamp 1604681595
transform 1 0 9844 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 10396 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10580 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604681595
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_122
timestamp 1604681595
transform 1 0 12328 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604681595
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13064 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_143
timestamp 1604681595
transform 1 0 14260 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_139
timestamp 1604681595
transform 1 0 13892 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_144
timestamp 1604681595
transform 1 0 14352 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_140
timestamp 1604681595
transform 1 0 13984 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604681595
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14168 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15640 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 14628 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_147
timestamp 1604681595
transform 1 0 14628 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_176
timestamp 1604681595
transform 1 0 17296 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_170
timestamp 1604681595
transform 1 0 16744 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 17112 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 17664 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 17480 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17572 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_177
timestamp 1604681595
transform 1 0 17388 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_181
timestamp 1604681595
transform 1 0 17756 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 17940 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18124 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18676 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19136 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_188
timestamp 1604681595
transform 1 0 18400 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1604681595
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_198
timestamp 1604681595
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1604681595
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1604681595
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_217
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_214
timestamp 1604681595
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_210
timestamp 1604681595
transform 1 0 20424 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_224
timestamp 1604681595
transform 1 0 21712 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_223
timestamp 1604681595
transform 1 0 21620 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 21804 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_229
timestamp 1604681595
transform 1 0 22172 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_239
timestamp 1604681595
transform 1 0 23092 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_235
timestamp 1604681595
transform 1 0 22724 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22908 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604681595
transform 1 0 22448 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604681595
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23276 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 23460 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604681595
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604681595
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1604681595
transform 1 0 25576 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_262
timestamp 1604681595
transform 1 0 25208 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25392 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 25208 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_268
timestamp 1604681595
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_276
timestamp 1604681595
transform 1 0 26496 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1472 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2852 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_13
timestamp 1604681595
transform 1 0 2300 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_17
timestamp 1604681595
transform 1 0 2668 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 3036 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_35_40
timestamp 1604681595
transform 1 0 4784 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604681595
transform 1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604681595
transform 1 0 5520 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1604681595
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1604681595
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7728 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 7544 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_68
timestamp 1604681595
transform 1 0 7360 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10028 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_91
timestamp 1604681595
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604681595
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1604681595
transform 1 0 10212 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_103
timestamp 1604681595
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1604681595
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13432 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_132
timestamp 1604681595
transform 1 0 13248 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1604681595
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1604681595
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1604681595
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_170
timestamp 1604681595
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_174
timestamp 1604681595
transform 1 0 17112 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604681595
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1604681595
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18768 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_35_189
timestamp 1604681595
transform 1 0 18492 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604681595
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21804 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1604681595
transform 1 0 20884 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_223
timestamp 1604681595
transform 1 0 21620 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 23644 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1604681595
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_240
timestamp 1604681595
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_264
timestamp 1604681595
transform 1 0 25392 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_268
timestamp 1604681595
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_272
timestamp 1604681595
transform 1 0 26128 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_276
timestamp 1604681595
transform 1 0 26496 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 1840 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_6
timestamp 1604681595
transform 1 0 1656 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_10
timestamp 1604681595
transform 1 0 2024 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 3772 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_23
timestamp 1604681595
transform 1 0 3220 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_41
timestamp 1604681595
transform 1 0 4876 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5980 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_45
timestamp 1604681595
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_49
timestamp 1604681595
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_62
timestamp 1604681595
transform 1 0 6808 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8556 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_66
timestamp 1604681595
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_79
timestamp 1604681595
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_83
timestamp 1604681595
transform 1 0 8740 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8924 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_87
timestamp 1604681595
transform 1 0 9108 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604681595
transform 1 0 12328 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 12144 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11408 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1604681595
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1604681595
transform 1 0 11224 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_114
timestamp 1604681595
transform 1 0 11592 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_118
timestamp 1604681595
transform 1 0 11960 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_131
timestamp 1604681595
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_135
timestamp 1604681595
transform 1 0 13524 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1604681595
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_163
timestamp 1604681595
transform 1 0 16100 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17020 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18308 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17940 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_167
timestamp 1604681595
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_171
timestamp 1604681595
transform 1 0 16836 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_179
timestamp 1604681595
transform 1 0 17572 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_185
timestamp 1604681595
transform 1 0 18124 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19320 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20148 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_196
timestamp 1604681595
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_200
timestamp 1604681595
transform 1 0 19504 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_205
timestamp 1604681595
transform 1 0 19964 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_215
timestamp 1604681595
transform 1 0 20884 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1604681595
transform 1 0 20700 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_209
timestamp 1604681595
transform 1 0 20332 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 20516 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604681595
transform 1 0 20976 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_224
timestamp 1604681595
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_220
timestamp 1604681595
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 21528 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_22.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 22080 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24012 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_247
timestamp 1604681595
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24564 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604681595
transform 1 0 25576 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_251
timestamp 1604681595
transform 1 0 24196 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1604681595
transform 1 0 25392 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_268
timestamp 1604681595
transform 1 0 25760 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1604681595
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604681595
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 2944 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604681595
transform 1 0 2760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2392 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_10
timestamp 1604681595
transform 1 0 2024 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_16
timestamp 1604681595
transform 1 0 2576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 4876 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604681595
transform 1 0 5428 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604681595
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5244 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_43
timestamp 1604681595
transform 1 0 5060 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_55
timestamp 1604681595
transform 1 0 6164 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 7360 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6992 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_66
timestamp 1604681595
transform 1 0 7176 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9476 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_87
timestamp 1604681595
transform 1 0 9108 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_93
timestamp 1604681595
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_97
timestamp 1604681595
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_101
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604681595
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604681595
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14352 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1604681595
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15456 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15272 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 14904 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_146
timestamp 1604681595
transform 1 0 14536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_152
timestamp 1604681595
transform 1 0 15088 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18216 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604681595
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604681595
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_184
timestamp 1604681595
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19780 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19228 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_195
timestamp 1604681595
transform 1 0 19044 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_199
timestamp 1604681595
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21712 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22080 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1604681595
transform 1 0 21528 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_226
timestamp 1604681595
transform 1 0 21896 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23644 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 22264 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1604681595
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_240
timestamp 1604681595
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604681595
transform 1 0 25208 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604681595
transform 1 0 25760 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24656 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_254
timestamp 1604681595
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_258
timestamp 1604681595
transform 1 0 24840 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_266
timestamp 1604681595
transform 1 0 25576 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_270
timestamp 1604681595
transform 1 0 25944 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604681595
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604681595
transform 1 0 2760 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1472 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_10
timestamp 1604681595
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_14
timestamp 1604681595
transform 1 0 2392 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4232 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_22
timestamp 1604681595
transform 1 0 3128 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_26
timestamp 1604681595
transform 1 0 3496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1604681595
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6716 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6532 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6164 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_53
timestamp 1604681595
transform 1 0 5980 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_57
timestamp 1604681595
transform 1 0 6348 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604681595
transform 1 0 8096 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7728 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_70
timestamp 1604681595
transform 1 0 7544 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_74
timestamp 1604681595
transform 1 0 7912 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9844 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9292 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_84
timestamp 1604681595
transform 1 0 8832 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1604681595
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_104
timestamp 1604681595
transform 1 0 10672 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11408 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10856 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11224 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1604681595
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13892 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13340 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_131
timestamp 1604681595
transform 1 0 13156 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_135
timestamp 1604681595
transform 1 0 13524 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1604681595
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 15364 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1604681595
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 1604681595
transform 1 0 15272 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17940 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17296 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 17756 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_174
timestamp 1604681595
transform 1 0 17112 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_178
timestamp 1604681595
transform 1 0 17480 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18676 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_189
timestamp 1604681595
transform 1 0 18492 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_193
timestamp 1604681595
transform 1 0 18860 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_206
timestamp 1604681595
transform 1 0 20056 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21160 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20608 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_210
timestamp 1604681595
transform 1 0 20424 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_215
timestamp 1604681595
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_20.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 23460 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_237
timestamp 1604681595
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_241
timestamp 1604681595
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604681595
transform 1 0 25208 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_254
timestamp 1604681595
transform 1 0 24472 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_266
timestamp 1604681595
transform 1 0 25576 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604681595
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1604681595
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604681595
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604681595
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1604681595
transform 1 0 2116 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_17
timestamp 1604681595
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_13
timestamp 1604681595
transform 1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_9
timestamp 1604681595
transform 1 0 1932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604681595
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604681595
transform 1 0 2116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1604681595
transform 1 0 2852 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1604681595
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_21
timestamp 1604681595
transform 1 0 3036 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_40
timestamp 1604681595
transform 1 0 4784 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_36
timestamp 1604681595
transform 1 0 4416 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_40
timestamp 1604681595
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_36
timestamp 1604681595
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604681595
transform 1 0 4600 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_46
timestamp 1604681595
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604681595
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604681595
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5704 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604681595
transform 1 0 8464 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8740 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1604681595
transform 1 0 8556 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_69
timestamp 1604681595
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_73
timestamp 1604681595
transform 1 0 7820 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_77
timestamp 1604681595
transform 1 0 8188 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_90
timestamp 1604681595
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_84
timestamp 1604681595
transform 1 0 8832 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_85
timestamp 1604681595
transform 1 0 8924 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9200 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9108 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9292 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_102
timestamp 1604681595
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_102
timestamp 1604681595
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_110
timestamp 1604681595
transform 1 0 11224 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_106
timestamp 1604681595
transform 1 0 10856 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604681595
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_106
timestamp 1604681595
transform 1 0 10856 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11040 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11316 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1604681595
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_117
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604681595
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12420 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604681595
transform 1 0 12604 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604681595
transform 1 0 14168 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 13800 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_142
timestamp 1604681595
transform 1 0 14168 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_134
timestamp 1604681595
transform 1 0 13432 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_140
timestamp 1604681595
transform 1 0 13984 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_148
timestamp 1604681595
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1604681595
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604681595
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_152
timestamp 1604681595
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_164
timestamp 1604681595
transform 1 0 16192 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_160
timestamp 1604681595
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1604681595
transform 1 0 16284 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 16008 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15456 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_174
timestamp 1604681595
transform 1 0 17112 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_170
timestamp 1604681595
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 16560 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_187
timestamp 1604681595
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_184
timestamp 1604681595
transform 1 0 18032 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604681595
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604681595
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 18124 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_18.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 16560 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19044 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 18860 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1604681595
transform 1 0 19872 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_208
timestamp 1604681595
transform 1 0 20240 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_191
timestamp 1604681595
transform 1 0 18676 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_204
timestamp 1604681595
transform 1 0 19872 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_208
timestamp 1604681595
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_215
timestamp 1604681595
transform 1 0 20884 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_212
timestamp 1604681595
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_211
timestamp 1604681595
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604681595
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604681595
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20884 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21068 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_226
timestamp 1604681595
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_228
timestamp 1604681595
transform 1 0 22080 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604681595
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22080 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_230
timestamp 1604681595
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_236
timestamp 1604681595
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22448 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22264 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604681595
transform 1 0 23000 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604681595
transform 1 0 22448 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_247
timestamp 1604681595
transform 1 0 23828 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_243
timestamp 1604681595
transform 1 0 23460 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_240
timestamp 1604681595
transform 1 0 23184 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 23644 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604681595
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 23644 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604681595
transform 1 0 24932 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604681595
transform 1 0 24564 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604681595
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604681595
transform 1 0 25484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1604681595
transform 1 0 24196 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_257
timestamp 1604681595
transform 1 0 24748 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_263
timestamp 1604681595
transform 1 0 25300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_267
timestamp 1604681595
transform 1 0 25668 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_259
timestamp 1604681595
transform 1 0 24932 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604681595
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604681595
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_271
timestamp 1604681595
transform 1 0 26036 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604681595
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604681595
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604681595
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604681595
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604681595
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1604681595
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604681595
transform 1 0 4692 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604681595
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604681595
transform 1 0 4140 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604681595
transform 1 0 4508 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604681595
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604681595
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1604681595
transform 1 0 4324 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604681595
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_43
timestamp 1604681595
transform 1 0 5060 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1604681595
transform 1 0 5428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1604681595
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7176 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8648 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_68
timestamp 1604681595
transform 1 0 7360 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_80
timestamp 1604681595
transform 1 0 8464 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9200 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604681595
transform 1 0 10672 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604681595
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_84
timestamp 1604681595
transform 1 0 8832 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_97
timestamp 1604681595
transform 1 0 10028 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_102
timestamp 1604681595
transform 1 0 10488 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604681595
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604681595
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_106
timestamp 1604681595
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604681595
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604681595
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1604681595
transform 1 0 13064 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 12880 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14076 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_127
timestamp 1604681595
transform 1 0 12788 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_139
timestamp 1604681595
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_3_
timestamp 1604681595
transform 1 0 16192 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__A1
timestamp 1604681595
transform 1 0 16008 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15640 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_156
timestamp 1604681595
transform 1 0 15456 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_160
timestamp 1604681595
transform 1 0 15824 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604681595
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_3__S
timestamp 1604681595
transform 1 0 17204 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_173
timestamp 1604681595
transform 1 0 17020 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1604681595
transform 1 0 17388 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19596 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1604681595
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_197
timestamp 1604681595
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21160 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20976 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22172 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_210
timestamp 1604681595
transform 1 0 20424 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_214
timestamp 1604681595
transform 1 0 20792 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_227
timestamp 1604681595
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604681595
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 22540 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 22908 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_231
timestamp 1604681595
transform 1 0 22356 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_235
timestamp 1604681595
transform 1 0 22724 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1604681595
transform 1 0 23092 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1604681595
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1604681595
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604681595
transform 1 0 24564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604681595
transform 1 0 25116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604681595
transform 1 0 24380 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_259
timestamp 1604681595
transform 1 0 24932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_263
timestamp 1604681595
transform 1 0 25300 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_275
timestamp 1604681595
transform 1 0 26404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_7
timestamp 1604681595
transform 1 0 1748 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_19
timestamp 1604681595
transform 1 0 2852 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604681595
transform 1 0 5152 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604681595
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7176 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_42_63
timestamp 1604681595
transform 1 0 6900 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_75
timestamp 1604681595
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604681595
transform 1 0 10304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_87
timestamp 1604681595
transform 1 0 9108 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_90
timestamp 1604681595
transform 1 0 9384 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_94
timestamp 1604681595
transform 1 0 9752 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1604681595
transform 1 0 10672 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604681595
transform 1 0 11408 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604681595
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_116
timestamp 1604681595
transform 1 0 11776 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_125
timestamp 1604681595
transform 1 0 12604 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604681595
transform 1 0 12696 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13800 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A0
timestamp 1604681595
transform 1 0 13248 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_130
timestamp 1604681595
transform 1 0 13064 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_134
timestamp 1604681595
transform 1 0 13432 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15732 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604681595
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604681595
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1604681595
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1604681595
transform 1 0 15456 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18308 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604681595
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_168
timestamp 1604681595
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1604681595
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604681595
transform 1 0 19872 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19596 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_196
timestamp 1604681595
transform 1 0 19136 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_200
timestamp 1604681595
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_203
timestamp 1604681595
transform 1 0 19780 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_208
timestamp 1604681595
transform 1 0 20240 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 21160 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604681595
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_214
timestamp 1604681595
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_227
timestamp 1604681595
transform 1 0 21988 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604681595
transform 1 0 22816 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604681595
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_235
timestamp 1604681595
transform 1 0 22724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_240
timestamp 1604681595
transform 1 0 23184 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_249
timestamp 1604681595
transform 1 0 24012 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604681595
transform 1 0 24564 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_259
timestamp 1604681595
transform 1 0 24932 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_271
timestamp 1604681595
transform 1 0 26036 0 -1 25568
box -38 -48 590 592
<< labels >>
rlabel metal2 s 19522 0 19578 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 294 27520 350 28000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 25134 0 25190 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 8298 0 8354 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 13910 0 13966 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 12384 480 12504 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 14288 480 14408 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 14832 480 14952 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 15376 480 15496 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 4496 480 4616 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 6944 480 7064 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 22720 480 22840 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 23400 480 23520 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 23944 480 24064 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 24624 480 24744 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 25168 480 25288 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 25848 480 25968 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 26392 480 26512 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 27072 480 27192 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 27616 480 27736 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 20272 480 20392 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 20952 480 21072 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 27520 3816 28000 3936 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 27520 9936 28000 10056 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 27520 10616 28000 10736 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 27520 11160 28000 11280 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 27520 12384 28000 12504 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 27520 4496 28000 4616 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 27520 5040 28000 5160 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 27520 5720 28000 5840 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 27520 6264 28000 6384 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 27520 7488 28000 7608 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 27520 8168 28000 8288 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 27520 8712 28000 8832 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 27520 9392 28000 9512 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 27520 16056 28000 16176 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 27520 22176 28000 22296 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 27520 22720 28000 22840 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 27520 23400 28000 23520 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 27520 23944 28000 24064 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 27520 24624 28000 24744 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 27520 25168 28000 25288 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 27520 25848 28000 25968 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 27520 26392 28000 26512 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 27520 27072 28000 27192 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 27520 27616 28000 27736 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 27520 17280 28000 17400 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 27520 17824 28000 17944 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 27520 18504 28000 18624 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 27520 19048 28000 19168 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 27520 19728 28000 19848 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 27520 20272 28000 20392 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 27520 20952 28000 21072 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 27520 21496 28000 21616 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 5262 27520 5318 28000 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 10874 27520 10930 28000 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 11426 27520 11482 28000 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 11978 27520 12034 28000 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 5814 27520 5870 28000 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 6366 27520 6422 28000 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 6918 27520 6974 28000 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 7562 27520 7618 28000 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 8114 27520 8170 28000 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 8666 27520 8722 28000 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 9218 27520 9274 28000 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 10322 27520 10378 28000 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 16486 27520 16542 28000 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 22098 27520 22154 28000 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 22650 27520 22706 28000 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 23202 27520 23258 28000 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 23754 27520 23810 28000 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 24306 27520 24362 28000 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 24858 27520 24914 28000 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 25410 27520 25466 28000 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 25962 27520 26018 28000 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 17590 27520 17646 28000 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 18142 27520 18198 28000 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 18694 27520 18750 28000 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 19246 27520 19302 28000 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 19798 27520 19854 28000 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 20350 27520 20406 28000 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 20902 27520 20958 28000 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 21546 27520 21602 28000 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 left_bottom_grid_pin_11_
port 126 nsew default input
rlabel metal3 s 0 280 480 400 6 left_bottom_grid_pin_1_
port 127 nsew default input
rlabel metal3 s 0 824 480 944 6 left_bottom_grid_pin_3_
port 128 nsew default input
rlabel metal3 s 0 1368 480 1488 6 left_bottom_grid_pin_5_
port 129 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_7_
port 130 nsew default input
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_9_
port 131 nsew default input
rlabel metal2 s 2778 0 2834 480 6 prog_clk
port 132 nsew default input
rlabel metal3 s 27520 3272 28000 3392 6 right_bottom_grid_pin_11_
port 133 nsew default input
rlabel metal3 s 27520 280 28000 400 6 right_bottom_grid_pin_1_
port 134 nsew default input
rlabel metal3 s 27520 824 28000 944 6 right_bottom_grid_pin_3_
port 135 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 right_bottom_grid_pin_5_
port 136 nsew default input
rlabel metal3 s 27520 2048 28000 2168 6 right_bottom_grid_pin_7_
port 137 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 right_bottom_grid_pin_9_
port 138 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_42_
port 139 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_43_
port 140 nsew default input
rlabel metal2 s 1950 27520 2006 28000 6 top_left_grid_pin_44_
port 141 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 top_left_grid_pin_45_
port 142 nsew default input
rlabel metal2 s 3054 27520 3110 28000 6 top_left_grid_pin_46_
port 143 nsew default input
rlabel metal2 s 3606 27520 3662 28000 6 top_left_grid_pin_47_
port 144 nsew default input
rlabel metal2 s 4158 27520 4214 28000 6 top_left_grid_pin_48_
port 145 nsew default input
rlabel metal2 s 4710 27520 4766 28000 6 top_left_grid_pin_49_
port 146 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 147 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 148 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
